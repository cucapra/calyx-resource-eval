
module std_fp_mult_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    input  logic             go,
    input  logic             clk,
    output logic [WIDTH-1:0] out,
    output logic             done
);
  logic [WIDTH-1:0]          rtmp;
  logic [WIDTH-1:0]          ltmp;
  logic [(WIDTH << 1) - 1:0] out_tmp;
  reg done_buf[1:0];
  always_ff @(posedge clk) begin
    if (go) begin
      rtmp <= right;
      ltmp <= left;
      out_tmp <= ltmp * rtmp;
      out <= out_tmp[(WIDTH << 1) - INT_WIDTH - 1 : WIDTH - INT_WIDTH];

      done <= done_buf[1];
      done_buf[0] <= 1'b1;
      done_buf[1] <= done_buf[0];
    end else begin
      rtmp <= 0;
      ltmp <= 0;
      out_tmp <= 0;
      out <= 0;

      done <= 0;
      done_buf[0] <= 0;
      done_buf[1] <= 0;
    end
  end
endmodule

module std_fp_add #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  assign out = left + right;
endmodule

module std_fp_sub #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module std_fp_gt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic             out
);
  assign out = left > right;
endmodule

module std_fp_add_dwidth #(
    parameter WIDTH1 = 32,
    parameter WIDTH2 = 32,
    parameter INT_WIDTH1 = 8,
    parameter FRACT_WIDTH1 = 24,
    parameter INT_WIDTH2 = 4,
    parameter FRACT_WIDTH2 = 28,
    parameter OUT_WIDTH = 36
) (
    input  logic [   WIDTH1-1:0] left,
    input  logic [   WIDTH2-1:0] right,
    output logic [OUT_WIDTH-1:0] out
);

  localparam BIG_INT = (INT_WIDTH1 >= INT_WIDTH2) ? INT_WIDTH1 : INT_WIDTH2;
  localparam BIG_FRACT = (FRACT_WIDTH1 >= FRACT_WIDTH2) ? FRACT_WIDTH1 : FRACT_WIDTH2;

  if (BIG_INT + BIG_FRACT != OUT_WIDTH)
    $error("std_fp_add_dwidth: Given output width not equal to computed output width");

  logic [INT_WIDTH1-1:0] left_int;
  logic [INT_WIDTH2-1:0] right_int;
  logic [FRACT_WIDTH1-1:0] left_fract;
  logic [FRACT_WIDTH2-1:0] right_fract;

  logic [BIG_INT-1:0] mod_right_int;
  logic [BIG_FRACT-1:0] mod_left_fract;

  logic [BIG_INT-1:0] whole_int;
  logic [BIG_FRACT-1:0] whole_fract;

  assign {left_int, left_fract} = left;
  assign {right_int, right_fract} = right;

  assign mod_left_fract = left_fract * (2 ** (FRACT_WIDTH2 - FRACT_WIDTH1));

  always_comb begin
    if ((mod_left_fract + right_fract) >= 2 ** FRACT_WIDTH2) begin
      whole_int = left_int + right_int + 1;
      whole_fract = mod_left_fract + right_fract - 2 ** FRACT_WIDTH2;
    end else begin
      whole_int = left_int + right_int;
      whole_fract = mod_left_fract + right_fract;
    end
  end

  assign out = {whole_int, whole_fract};
endmodule

/// ========================= Unsynthesizable primitives =====================

module std_fp_mult #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  logic [2*WIDTH-2:0] result;

  assign result = left * right;
  assign out = result[WIDTH+FRACT_WIDTH-1:FRACT_WIDTH];
endmodule

module std_fp_div #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  logic [2*WIDTH-2:0] result;

  assign result = left / right;
  assign out = result[WIDTH+FRACT_WIDTH-1:FRACT_WIDTH];
endmodule
module std_fp_smult_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  signed       [WIDTH-1:0] left,
    input  signed       [WIDTH-1:0] right,
    input  logic                    go,
    input  logic                    clk,
    output logic signed [WIDTH-1:0] out,
    output logic                    done
);
  logic signed [WIDTH-1:0] rtmp;
  logic signed [WIDTH-1:0] ltmp;
  logic signed [(WIDTH << 1) - 1:0] out_tmp;
  reg done_buf[1:0];
  always_ff @(posedge clk) begin
    if (go) begin
      ltmp <= left;
      rtmp <= right;
      // Sign extend by the first bit for the operands.
      out_tmp <= $signed(
                   { {WIDTH{ltmp[WIDTH-1]}}, ltmp} *
                   { {WIDTH{rtmp[WIDTH-1]}}, rtmp}
                 );
      out <= out_tmp[(WIDTH << 1) - INT_WIDTH - 1: WIDTH - INT_WIDTH];

      done <= done_buf[1];
      done_buf[0] <= 1'b1;
      done_buf[1] <= done_buf[0];
    end else begin
      rtmp <= 0;
      ltmp <= 0;
      out_tmp <= 0;
      out <= 0;

      done <= 0;
      done_buf[0] <= 0;
      done_buf[1] <= 0;
    end
  end
endmodule

module std_fp_sadd #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left + right);
endmodule

module std_fp_ssub #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);

  assign out = $signed(left - right);
endmodule

module std_fp_sadd_dwidth #(
    parameter WIDTH1 = 32,
    parameter WIDTH2 = 32,
    parameter INT_WIDTH1 = 8,
    parameter FRACT_WIDTH1 = 24,
    parameter INT_WIDTH2 = 4,
    parameter FRACT_WIDTH2 = 28,
    parameter OUT_WIDTH = 36
) (
    input  logic [   WIDTH1-1:0] left,
    input  logic [   WIDTH2-1:0] right,
    output logic [OUT_WIDTH-1:0] out
);

  logic signed [INT_WIDTH1-1:0] left_int;
  logic signed [INT_WIDTH2-1:0] right_int;
  logic [FRACT_WIDTH1-1:0] left_fract;
  logic [FRACT_WIDTH2-1:0] right_fract;

  localparam BIG_INT = (INT_WIDTH1 >= INT_WIDTH2) ? INT_WIDTH1 : INT_WIDTH2;
  localparam BIG_FRACT = (FRACT_WIDTH1 >= FRACT_WIDTH2) ? FRACT_WIDTH1 : FRACT_WIDTH2;

  logic [BIG_INT-1:0] mod_right_int;
  logic [BIG_FRACT-1:0] mod_left_fract;

  logic [BIG_INT-1:0] whole_int;
  logic [BIG_FRACT-1:0] whole_fract;

  assign {left_int, left_fract} = left;
  assign {right_int, right_fract} = right;

  assign mod_left_fract = left_fract * (2 ** (FRACT_WIDTH2 - FRACT_WIDTH1));

  always_comb begin
    if ((mod_left_fract + right_fract) >= 2 ** FRACT_WIDTH2) begin
      whole_int = $signed(left_int + right_int + 1);
      whole_fract = mod_left_fract + right_fract - 2 ** FRACT_WIDTH2;
    end else begin
      whole_int = $signed(left_int + right_int);
      whole_fract = mod_left_fract + right_fract;
    end
  end

  assign out = {whole_int, whole_fract};
endmodule

module std_fp_sgt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  logic signed [WIDTH-1:0] left,
    input  logic signed [WIDTH-1:0] right,
    output logic signed             out
);
  assign out = $signed(left > right);
endmodule

module std_fp_smult #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);

  logic [2*WIDTH-2:0] result;

  assign result = $signed(left * right);
  assign out = result[WIDTH+FRACT_WIDTH-1:FRACT_WIDTH];
endmodule

module std_fp_sdiv #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);

  logic [2*WIDTH-2:0] result;

  assign result = $signed(left / right);
  assign out = result[WIDTH+FRACT_WIDTH-1:FRACT_WIDTH];
endmodule

/* verilator lint_off WIDTH */
module std_div_pipe #(
    parameter width = 32
) (
    input                    clk,
    input                    go,
    input        [width-1:0] left,
    input        [width-1:0] right,
    output logic [width-1:0] out_remainder,
    output logic [width-1:0] out_quotient,
    output logic             done
);

  logic [width-1:0] dividend;
  logic [(width-1)*2:0] divisor;
  logic [width-1:0] quotient;
  logic [width-1:0] quotient_msk;
  logic start, running, finished;

  assign start = go && !running;
  assign finished = !quotient_msk && running;

  always @(posedge clk) begin
    if (!go) begin
      running <= 0;
      done <= 0;
      out_remainder <= 0;
      out_quotient <= 0;
    end else if (start && left == 0) begin
      out_remainder <= 0;
      out_quotient <= 0;
      done <= 1;
    end

    if (start) begin
      running <= 1;
      dividend <= left;
      divisor <= right << width - 1;
      quotient <= 0;
      quotient_msk <= 1 << width - 1;
    end else if (finished) begin
      running <= 0;
      done <= 1;
      out_remainder <= dividend;
      out_quotient <= quotient;
    end else begin
      if (divisor <= dividend) begin
        dividend <= dividend - divisor;
        quotient <= quotient | quotient_msk;
      end
      divisor <= divisor >> 1;
      quotient_msk <= quotient_msk >> 1;
    end
  end

  `ifdef VERILATOR
    // Simulation self test against unsynthesizable implementation.
    always @(posedge clk) begin
      if (finished && dividend != $unsigned(left % right))
        $error(
          "\nstd_div_pipe (Remainder): Computed and golden outputs do not match!\n",
          "left: %0d", $unsigned(left),
          "  right: %0d\n", $unsigned(right),
          "expected: %0d", $unsigned(left % right),
          "  computed: %0d", $unsigned(dividend)
        );
      if (finished && quotient != $unsigned(left / right))
        $error(
          "\nstd_div_pipe (Quotient): Computed and golden outputs do not match!\n",
          "left: %0d", $unsigned(left),
          "  right: %0d\n", $unsigned(right),
          "expected: %0d", $unsigned(left / right),
          "  computed: %0d", $unsigned(quotient)
        );
    end
  `endif
endmodule

module std_mult_pipe #(
    parameter width = 32
) (
    input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    input  logic             go,
    input  logic             clk,
    output logic [width-1:0] out,
    output logic             done
);
  logic [width-1:0] rtmp;
  logic [width-1:0] ltmp;
  logic [width-1:0] out_tmp;
  reg done_buf[1:0];
  always_ff @(posedge clk) begin
    if (go) begin
      rtmp <= right;
      ltmp <= left;
      out_tmp <= rtmp * ltmp;
      out <= out_tmp;

      done <= done_buf[1];
      done_buf[0] <= 1'b1;
      done_buf[1] <= done_buf[0];
    end else begin
      rtmp <= 0;
      ltmp <= 0;
      out_tmp <= 0;
      out <= 0;

      done <= 0;
      done_buf[0] <= 0;
      done_buf[1] <= 0;
    end
  end
endmodule

// ===============Signed operations that wrap unsigned ones ===============

/* verilator lint_off WIDTH */
module std_sdiv_pipe #(
    parameter width = 32
) (
    input                     clk,
    input                     go,
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output logic  [width-1:0] out_quotient,
    output logic  [width-1:0] out_remainder,
    output logic              done
);

  logic signed [width-1:0] left_abs;
  logic signed [width-1:0] right_abs;
  logic signed [width-1:0] comp_out_q;
  logic signed [width-1:0] comp_out_r;

  assign right_abs = right[width-1] == 1 ? -right : right;
  assign left_abs = left[width-1] == 1 ? -left : left;
  assign out_quotient =
    (left[width-1] == 1) ^ (right[width-1] == 1) ? -comp_out_q : comp_out_q;
  assign out_remainder = left[width-1] == 1 ? $signed(right - comp_out_r) : comp_out_r;

  std_div_pipe #(
    .width(width)
  ) comp (
    .clk(clk),
    .done(done),
    .go(go),
    .left(left_abs),
    .right(right_abs),
    .out_quotient(comp_out_q),
    .out_remainder(comp_out_r)
  );

  `ifdef VERILATOR
    // Simulation self test against unsynthesizable implementation.
    always @(posedge clk) begin
      if (done && out_quotient != $signed(left / right))
        $error(
          "\nstd_sdiv_pipe (Quotient): Computed and golden outputs do not match!\n",
          "left: %0d", left,
          "  right: %0d\n", right,
          "expected: %0d", $signed(left / right),
          "  computed: %0d", $signed(out_quotient)
        );
      if (done && out_remainder != $signed(((left % right) + right) % right))
        $error(
          "\nstd_sdiv_pipe (Remainder): Computed and golden outputs do not match!\n",
          "left: %0d", left,
          "  right: %0d\n", right,
          "expected: %0d", $signed(((left % right) + right) % right),
          "  computed: %0d", $signed(out_remainder)
        );
    end
  `endif
endmodule


//==================== Unsynthesizable primitives =========================
module std_mult #(
    parameter width = 32
) (
    input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    output logic [width-1:0] out
);
  assign out = left * right;
endmodule

module std_div #(
    parameter width = 32
) (
    input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    output logic [width-1:0] out
);
  assign out = left / right;
endmodule

module std_mod #(
    parameter width = 32
) (
    input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    output logic [width-1:0] out
);
  assign out = left % right;
endmodule
/**
* Signed arthimetic primitives for FuTIL.
*/

module std_slsh #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed [width-1:0] out
);
  assign out = left <<< right;
endmodule

module std_srsh #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed [width-1:0] out
);
  assign out = left >>> right;
endmodule

module std_sadd #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed [width-1:0] out
);
  assign out = $signed(left + right);
endmodule

module std_ssub #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed [width-1:0] out
);
  assign out = $signed(left - right);
endmodule

module std_smult_pipe #(
    parameter width = 32
) (
    input  logic                    go,
    input  logic                    clk,
    input  signed       [width-1:0] left,
    input  signed       [width-1:0] right,
    output logic signed [width-1:0] out,
    output logic                    done
);
  logic signed [width-1:0] rtmp;
  logic signed [width-1:0] ltmp;
  logic signed [width-1:0] out_tmp;
  logic done_buf[1:0];

  always_ff @(posedge clk) begin
    if (go) begin
      rtmp <= right;
      ltmp <= left;
      out_tmp <= $signed(rtmp * ltmp);
      out <= out_tmp;

      done <= done_buf[1];
      done_buf[0] <= 1'b1;
      done_buf[1] <= done_buf[0];
    end else begin
      rtmp <= 0;
      ltmp <= 0;
      out_tmp <= 0;
      out <= 0;

      done <= 0;
      done_buf[0] <= 0;
      done_buf[1] <= 0;
    end
  end
endmodule

module std_sgt #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed             out
);
  assign out = $signed(left > right);
endmodule

module std_slt #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed             out
);
  assign out = $signed(left < right);
endmodule

module std_seq #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed             out
);
  assign out = $signed(left == right);
endmodule

module std_sneq #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed             out
);
  assign out = $signed(left != right);
endmodule

module std_sge #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed             out
);
  assign out = $signed(left >= right);
endmodule

module std_sle #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed             out
);
  assign out = $signed(left <= right);
endmodule

module std_sdiv #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed [width-1:0] out
);
  assign out = $signed(left / right);
endmodule

module std_smod #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed [width-1:0] out
);
  assign out = $signed(left % right);
endmodule


module std_smult #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed [width-1:0] out
);
  assign out = $signed(left * right);
endmodule

/**
 * Core primitives for FuTIL.
 * Implements core primitives used by the compiler.
 *
 * Conventions:
 * - All parameter names must be SNAKE_CASE and all caps.
 * - Port names must be snake_case, no caps.
 */
`default_nettype none

module std_mem_d1 #(
    parameter width = 32,
    parameter size = 16,
    parameter idx_size = 4
) (
   input wire                logic [idx_size-1:0] addr0,
   input wire                logic [ width-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   output logic [ width-1:0] read_data,
   output logic              done
);

  logic [width-1:0] mem[size-1:0];

  /* verilator lint_off WIDTH */
  assign read_data = mem[addr0];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0] <= write_data;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module std_mem_d2 #(
    parameter width = 32,
    parameter d0_size = 16,
    parameter d1_size = 16,
    parameter d0_idx_size = 4,
    parameter d1_idx_size = 4
) (
   input wire                logic [d0_idx_size-1:0] addr0,
   input wire                logic [d1_idx_size-1:0] addr1,
   input wire                logic [ width-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   output logic [ width-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [width-1:0] mem[d0_size-1:0][d1_size-1:0];

  assign read_data = mem[addr0][addr1];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0][addr1] <= write_data;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module std_mem_d3 #(
    parameter width = 32,
    parameter d0_size = 16,
    parameter d1_size = 16,
    parameter d2_size = 16,
    parameter d0_idx_size = 4,
    parameter d1_idx_size = 4,
    parameter d2_idx_size = 4
) (
   input wire                logic [d0_idx_size-1:0] addr0,
   input wire                logic [d1_idx_size-1:0] addr1,
   input wire                logic [d2_idx_size-1:0] addr2,
   input wire                logic [ width-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   output logic [ width-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [width-1:0] mem[d0_size-1:0][d1_size-1:0][d2_size-1:0];

  assign read_data = mem[addr0][addr1][addr2];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0][addr1][addr2] <= write_data;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module std_mem_d4 #(
    parameter width = 32,
    parameter d0_size = 16,
    parameter d1_size = 16,
    parameter d2_size = 16,
    parameter d3_size = 16,
    parameter d0_idx_size = 4,
    parameter d1_idx_size = 4,
    parameter d2_idx_size = 4,
    parameter d3_idx_size = 4
) (
   input wire                logic [d0_idx_size-1:0] addr0,
   input wire                logic [d1_idx_size-1:0] addr1,
   input wire                logic [d2_idx_size-1:0] addr2,
   input wire                logic [d3_idx_size-1:0] addr3,
   input wire                logic [ width-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   output logic [ width-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [width-1:0] mem[d0_size-1:0][d1_size-1:0][d2_size-1:0][d3_size-1:0];

  assign read_data = mem[addr0][addr1][addr2][addr3];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0][addr1][addr2][addr3] <= write_data;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module std_reg #(
    parameter width = 32
) (
   input wire [ width-1:0]    in,
   input wire                 write_en,
   input wire                 clk,
    // output
   output logic [width - 1:0] out,
   output logic               done
);

  always_ff @(posedge clk) begin
    if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module std_const #(
    parameter width = 32,
    parameter value = 0
) (
   output logic [width - 1:0] out
);
  assign out = value;
endmodule

module std_slice #(
    parameter in_width  = 32,
    parameter out_width = 32
) (
   input wire                   logic [ in_width-1:0] in,
   output logic [out_width-1:0] out
);
  assign out = in[out_width-1:0];

  `ifdef VERILATOR
    always_comb begin
      if (in_width < out_width)
        $error(
          "std_slice: Input width less than output width\n",
          "in_width: %0d", in_width,
          "out_width: %0d", out_width
        );
    end
  `endif
endmodule

module std_pad #(
    parameter in_width  = 32,
    parameter out_width = 32
) (
   input wire                   logic [ in_width-1:0] in,
   output logic [out_width-1:0] out
);
  localparam EXTEND = out_width - in_width;
  assign out = { {EXTEND {1'b0}}, in};

  `ifdef VERILATOR
    always_comb begin
      if (in_width > out_width)
        $error(
          "std_pad: Output width less than input width\n",
          "in_width: %0d", in_width,
          "out_width: %0d", out_width
        );
    end
  `endif
endmodule

module std_lsh #(
    parameter width = 32
) (
   input wire               logic [width-1:0] left,
   input wire               logic [width-1:0] right,
   output logic [width-1:0] out
);
  assign out = left << right;
endmodule

module std_rsh #(
    parameter width = 32
) (
   input wire               logic [width-1:0] left,
   input wire               logic [width-1:0] right,
   output logic [width-1:0] out
);
  assign out = left >> right;
endmodule

module std_add #(
    parameter width = 32
) (
   input wire               logic [width-1:0] left,
   input wire               logic [width-1:0] right,
   output logic [width-1:0] out
);
  assign out = left + right;
endmodule

module std_sub #(
    parameter width = 32
) (
   input wire               logic [width-1:0] left,
   input wire               logic [width-1:0] right,
   output logic [width-1:0] out
);
  assign out = left - right;
endmodule

module std_not #(
    parameter width = 32
) (
   input wire               logic [width-1:0] in,
   output logic [width-1:0] out
);
  assign out = ~in;
endmodule

module std_and #(
    parameter width = 32
) (
   input wire               logic [width-1:0] left,
   input wire               logic [width-1:0] right,
   output logic [width-1:0] out
);
  assign out = left & right;
endmodule

module std_or #(
    parameter width = 32
) (
   input wire               logic [width-1:0] left,
   input wire               logic [width-1:0] right,
   output logic [width-1:0] out
);
  assign out = left | right;
endmodule

module std_xor #(
    parameter width = 32
) (
   input wire               logic [width-1:0] left,
   input wire               logic [width-1:0] right,
   output logic [width-1:0] out
);
  assign out = left ^ right;
endmodule

module std_gt #(
    parameter width = 32
) (
   input wire   logic [width-1:0] left,
   input wire   logic [width-1:0] right,
   output logic out
);
  assign out = left > right;
endmodule

module std_lt #(
    parameter width = 32
) (
   input wire   logic [width-1:0] left,
   input wire   logic [width-1:0] right,
   output logic out
);
  assign out = left < right;
endmodule

module std_eq #(
    parameter width = 32
) (
   input wire   logic [width-1:0] left,
   input wire   logic [width-1:0] right,
   output logic out
);
  assign out = left == right;
endmodule

module std_neq #(
    parameter width = 32
) (
   input wire   logic [width-1:0] left,
   input wire   logic [width-1:0] right,
   output logic out
);
  assign out = left != right;
endmodule

module std_ge #(
    parameter width = 32
) (
    input wire   logic [width-1:0] left,
    input wire   logic [width-1:0] right,
    output logic out
);
  assign out = left >= right;
endmodule

module std_le #(
    parameter width = 32
) (
   input wire   logic [width-1:0] left,
   input wire   logic [width-1:0] right,
   output logic out
);
  assign out = left <= right;
endmodule

`default_nettype wire
module main (
    input logic go,
    input logic clk,
    output logic done,
    output logic [3:0] t0_addr0,
    output logic [31:0] t0_write_data,
    output logic t0_write_en,
    output logic t0_clk,
    input logic [31:0] t0_read_data,
    input logic t0_done,
    output logic [3:0] t1_addr0,
    output logic [31:0] t1_write_data,
    output logic t1_write_en,
    output logic t1_clk,
    input logic [31:0] t1_read_data,
    input logic t1_done,
    output logic [3:0] t2_addr0,
    output logic [31:0] t2_write_data,
    output logic t2_write_en,
    output logic t2_clk,
    input logic [31:0] t2_read_data,
    input logic t2_done,
    output logic [3:0] t3_addr0,
    output logic [31:0] t3_write_data,
    output logic t3_write_en,
    output logic t3_clk,
    input logic [31:0] t3_read_data,
    input logic t3_done,
    output logic [3:0] t4_addr0,
    output logic [31:0] t4_write_data,
    output logic t4_write_en,
    output logic t4_clk,
    input logic [31:0] t4_read_data,
    input logic t4_done,
    output logic [3:0] t5_addr0,
    output logic [31:0] t5_write_data,
    output logic t5_write_en,
    output logic t5_clk,
    input logic [31:0] t5_read_data,
    input logic t5_done,
    output logic [3:0] t6_addr0,
    output logic [31:0] t6_write_data,
    output logic t6_write_en,
    output logic t6_clk,
    input logic [31:0] t6_read_data,
    input logic t6_done,
    output logic [3:0] t7_addr0,
    output logic [31:0] t7_write_data,
    output logic t7_write_en,
    output logic t7_clk,
    input logic [31:0] t7_read_data,
    input logic t7_done,
    output logic [3:0] l0_addr0,
    output logic [31:0] l0_write_data,
    output logic l0_write_en,
    output logic l0_clk,
    input logic [31:0] l0_read_data,
    input logic l0_done,
    output logic [3:0] l1_addr0,
    output logic [31:0] l1_write_data,
    output logic l1_write_en,
    output logic l1_clk,
    input logic [31:0] l1_read_data,
    input logic l1_done,
    output logic [3:0] l2_addr0,
    output logic [31:0] l2_write_data,
    output logic l2_write_en,
    output logic l2_clk,
    input logic [31:0] l2_read_data,
    input logic l2_done,
    output logic [3:0] l3_addr0,
    output logic [31:0] l3_write_data,
    output logic l3_write_en,
    output logic l3_clk,
    input logic [31:0] l3_read_data,
    input logic l3_done,
    output logic [3:0] l4_addr0,
    output logic [31:0] l4_write_data,
    output logic l4_write_en,
    output logic l4_clk,
    input logic [31:0] l4_read_data,
    input logic l4_done,
    output logic [3:0] l5_addr0,
    output logic [31:0] l5_write_data,
    output logic l5_write_en,
    output logic l5_clk,
    input logic [31:0] l5_read_data,
    input logic l5_done,
    output logic [3:0] l6_addr0,
    output logic [31:0] l6_write_data,
    output logic l6_write_en,
    output logic l6_clk,
    input logic [31:0] l6_read_data,
    input logic l6_done,
    output logic [3:0] l7_addr0,
    output logic [31:0] l7_write_data,
    output logic l7_write_en,
    output logic l7_clk,
    input logic [31:0] l7_read_data,
    input logic l7_done
);
    logic [3:0] t0_idx_in;
    logic t0_idx_write_en;
    logic t0_idx_clk;
    logic [3:0] t0_idx_out;
    logic t0_idx_done;
    logic [3:0] t0_add_left;
    logic [3:0] t0_add_right;
    logic [3:0] t0_add_out;
    logic [3:0] t1_idx_in;
    logic t1_idx_write_en;
    logic t1_idx_clk;
    logic [3:0] t1_idx_out;
    logic t1_idx_done;
    logic [3:0] t1_add_left;
    logic [3:0] t1_add_right;
    logic [3:0] t1_add_out;
    logic [3:0] t2_idx_in;
    logic t2_idx_write_en;
    logic t2_idx_clk;
    logic [3:0] t2_idx_out;
    logic t2_idx_done;
    logic [3:0] t2_add_left;
    logic [3:0] t2_add_right;
    logic [3:0] t2_add_out;
    logic [3:0] t3_idx_in;
    logic t3_idx_write_en;
    logic t3_idx_clk;
    logic [3:0] t3_idx_out;
    logic t3_idx_done;
    logic [3:0] t3_add_left;
    logic [3:0] t3_add_right;
    logic [3:0] t3_add_out;
    logic [3:0] t4_idx_in;
    logic t4_idx_write_en;
    logic t4_idx_clk;
    logic [3:0] t4_idx_out;
    logic t4_idx_done;
    logic [3:0] t4_add_left;
    logic [3:0] t4_add_right;
    logic [3:0] t4_add_out;
    logic [3:0] t5_idx_in;
    logic t5_idx_write_en;
    logic t5_idx_clk;
    logic [3:0] t5_idx_out;
    logic t5_idx_done;
    logic [3:0] t5_add_left;
    logic [3:0] t5_add_right;
    logic [3:0] t5_add_out;
    logic [3:0] t6_idx_in;
    logic t6_idx_write_en;
    logic t6_idx_clk;
    logic [3:0] t6_idx_out;
    logic t6_idx_done;
    logic [3:0] t6_add_left;
    logic [3:0] t6_add_right;
    logic [3:0] t6_add_out;
    logic [3:0] t7_idx_in;
    logic t7_idx_write_en;
    logic t7_idx_clk;
    logic [3:0] t7_idx_out;
    logic t7_idx_done;
    logic [3:0] t7_add_left;
    logic [3:0] t7_add_right;
    logic [3:0] t7_add_out;
    logic [3:0] l0_idx_in;
    logic l0_idx_write_en;
    logic l0_idx_clk;
    logic [3:0] l0_idx_out;
    logic l0_idx_done;
    logic [3:0] l0_add_left;
    logic [3:0] l0_add_right;
    logic [3:0] l0_add_out;
    logic [3:0] l1_idx_in;
    logic l1_idx_write_en;
    logic l1_idx_clk;
    logic [3:0] l1_idx_out;
    logic l1_idx_done;
    logic [3:0] l1_add_left;
    logic [3:0] l1_add_right;
    logic [3:0] l1_add_out;
    logic [3:0] l2_idx_in;
    logic l2_idx_write_en;
    logic l2_idx_clk;
    logic [3:0] l2_idx_out;
    logic l2_idx_done;
    logic [3:0] l2_add_left;
    logic [3:0] l2_add_right;
    logic [3:0] l2_add_out;
    logic [3:0] l3_idx_in;
    logic l3_idx_write_en;
    logic l3_idx_clk;
    logic [3:0] l3_idx_out;
    logic l3_idx_done;
    logic [3:0] l3_add_left;
    logic [3:0] l3_add_right;
    logic [3:0] l3_add_out;
    logic [3:0] l4_idx_in;
    logic l4_idx_write_en;
    logic l4_idx_clk;
    logic [3:0] l4_idx_out;
    logic l4_idx_done;
    logic [3:0] l4_add_left;
    logic [3:0] l4_add_right;
    logic [3:0] l4_add_out;
    logic [3:0] l5_idx_in;
    logic l5_idx_write_en;
    logic l5_idx_clk;
    logic [3:0] l5_idx_out;
    logic l5_idx_done;
    logic [3:0] l5_add_left;
    logic [3:0] l5_add_right;
    logic [3:0] l5_add_out;
    logic [3:0] l6_idx_in;
    logic l6_idx_write_en;
    logic l6_idx_clk;
    logic [3:0] l6_idx_out;
    logic l6_idx_done;
    logic [3:0] l6_add_left;
    logic [3:0] l6_add_right;
    logic [3:0] l6_add_out;
    logic [3:0] l7_idx_in;
    logic l7_idx_write_en;
    logic l7_idx_clk;
    logic [3:0] l7_idx_out;
    logic l7_idx_done;
    logic [3:0] l7_add_left;
    logic [3:0] l7_add_right;
    logic [3:0] l7_add_out;
    logic [31:0] pe_0_0_top;
    logic [31:0] pe_0_0_left;
    logic [31:0] pe_0_0_out;
    logic pe_0_0_go;
    logic pe_0_0_clk;
    logic pe_0_0_done;
    logic [31:0] top_0_0_in;
    logic top_0_0_write_en;
    logic top_0_0_clk;
    logic [31:0] top_0_0_out;
    logic top_0_0_done;
    logic [31:0] left_0_0_in;
    logic left_0_0_write_en;
    logic left_0_0_clk;
    logic [31:0] left_0_0_out;
    logic left_0_0_done;
    logic [31:0] pe_0_1_top;
    logic [31:0] pe_0_1_left;
    logic [31:0] pe_0_1_out;
    logic pe_0_1_go;
    logic pe_0_1_clk;
    logic pe_0_1_done;
    logic [31:0] top_0_1_in;
    logic top_0_1_write_en;
    logic top_0_1_clk;
    logic [31:0] top_0_1_out;
    logic top_0_1_done;
    logic [31:0] left_0_1_in;
    logic left_0_1_write_en;
    logic left_0_1_clk;
    logic [31:0] left_0_1_out;
    logic left_0_1_done;
    logic [31:0] pe_0_2_top;
    logic [31:0] pe_0_2_left;
    logic [31:0] pe_0_2_out;
    logic pe_0_2_go;
    logic pe_0_2_clk;
    logic pe_0_2_done;
    logic [31:0] top_0_2_in;
    logic top_0_2_write_en;
    logic top_0_2_clk;
    logic [31:0] top_0_2_out;
    logic top_0_2_done;
    logic [31:0] left_0_2_in;
    logic left_0_2_write_en;
    logic left_0_2_clk;
    logic [31:0] left_0_2_out;
    logic left_0_2_done;
    logic [31:0] pe_0_3_top;
    logic [31:0] pe_0_3_left;
    logic [31:0] pe_0_3_out;
    logic pe_0_3_go;
    logic pe_0_3_clk;
    logic pe_0_3_done;
    logic [31:0] top_0_3_in;
    logic top_0_3_write_en;
    logic top_0_3_clk;
    logic [31:0] top_0_3_out;
    logic top_0_3_done;
    logic [31:0] left_0_3_in;
    logic left_0_3_write_en;
    logic left_0_3_clk;
    logic [31:0] left_0_3_out;
    logic left_0_3_done;
    logic [31:0] pe_0_4_top;
    logic [31:0] pe_0_4_left;
    logic [31:0] pe_0_4_out;
    logic pe_0_4_go;
    logic pe_0_4_clk;
    logic pe_0_4_done;
    logic [31:0] top_0_4_in;
    logic top_0_4_write_en;
    logic top_0_4_clk;
    logic [31:0] top_0_4_out;
    logic top_0_4_done;
    logic [31:0] left_0_4_in;
    logic left_0_4_write_en;
    logic left_0_4_clk;
    logic [31:0] left_0_4_out;
    logic left_0_4_done;
    logic [31:0] pe_0_5_top;
    logic [31:0] pe_0_5_left;
    logic [31:0] pe_0_5_out;
    logic pe_0_5_go;
    logic pe_0_5_clk;
    logic pe_0_5_done;
    logic [31:0] top_0_5_in;
    logic top_0_5_write_en;
    logic top_0_5_clk;
    logic [31:0] top_0_5_out;
    logic top_0_5_done;
    logic [31:0] left_0_5_in;
    logic left_0_5_write_en;
    logic left_0_5_clk;
    logic [31:0] left_0_5_out;
    logic left_0_5_done;
    logic [31:0] pe_0_6_top;
    logic [31:0] pe_0_6_left;
    logic [31:0] pe_0_6_out;
    logic pe_0_6_go;
    logic pe_0_6_clk;
    logic pe_0_6_done;
    logic [31:0] top_0_6_in;
    logic top_0_6_write_en;
    logic top_0_6_clk;
    logic [31:0] top_0_6_out;
    logic top_0_6_done;
    logic [31:0] left_0_6_in;
    logic left_0_6_write_en;
    logic left_0_6_clk;
    logic [31:0] left_0_6_out;
    logic left_0_6_done;
    logic [31:0] pe_0_7_top;
    logic [31:0] pe_0_7_left;
    logic [31:0] pe_0_7_out;
    logic pe_0_7_go;
    logic pe_0_7_clk;
    logic pe_0_7_done;
    logic [31:0] top_0_7_in;
    logic top_0_7_write_en;
    logic top_0_7_clk;
    logic [31:0] top_0_7_out;
    logic top_0_7_done;
    logic [31:0] left_0_7_in;
    logic left_0_7_write_en;
    logic left_0_7_clk;
    logic [31:0] left_0_7_out;
    logic left_0_7_done;
    logic [31:0] pe_1_0_top;
    logic [31:0] pe_1_0_left;
    logic [31:0] pe_1_0_out;
    logic pe_1_0_go;
    logic pe_1_0_clk;
    logic pe_1_0_done;
    logic [31:0] top_1_0_in;
    logic top_1_0_write_en;
    logic top_1_0_clk;
    logic [31:0] top_1_0_out;
    logic top_1_0_done;
    logic [31:0] left_1_0_in;
    logic left_1_0_write_en;
    logic left_1_0_clk;
    logic [31:0] left_1_0_out;
    logic left_1_0_done;
    logic [31:0] pe_1_1_top;
    logic [31:0] pe_1_1_left;
    logic [31:0] pe_1_1_out;
    logic pe_1_1_go;
    logic pe_1_1_clk;
    logic pe_1_1_done;
    logic [31:0] top_1_1_in;
    logic top_1_1_write_en;
    logic top_1_1_clk;
    logic [31:0] top_1_1_out;
    logic top_1_1_done;
    logic [31:0] left_1_1_in;
    logic left_1_1_write_en;
    logic left_1_1_clk;
    logic [31:0] left_1_1_out;
    logic left_1_1_done;
    logic [31:0] pe_1_2_top;
    logic [31:0] pe_1_2_left;
    logic [31:0] pe_1_2_out;
    logic pe_1_2_go;
    logic pe_1_2_clk;
    logic pe_1_2_done;
    logic [31:0] top_1_2_in;
    logic top_1_2_write_en;
    logic top_1_2_clk;
    logic [31:0] top_1_2_out;
    logic top_1_2_done;
    logic [31:0] left_1_2_in;
    logic left_1_2_write_en;
    logic left_1_2_clk;
    logic [31:0] left_1_2_out;
    logic left_1_2_done;
    logic [31:0] pe_1_3_top;
    logic [31:0] pe_1_3_left;
    logic [31:0] pe_1_3_out;
    logic pe_1_3_go;
    logic pe_1_3_clk;
    logic pe_1_3_done;
    logic [31:0] top_1_3_in;
    logic top_1_3_write_en;
    logic top_1_3_clk;
    logic [31:0] top_1_3_out;
    logic top_1_3_done;
    logic [31:0] left_1_3_in;
    logic left_1_3_write_en;
    logic left_1_3_clk;
    logic [31:0] left_1_3_out;
    logic left_1_3_done;
    logic [31:0] pe_1_4_top;
    logic [31:0] pe_1_4_left;
    logic [31:0] pe_1_4_out;
    logic pe_1_4_go;
    logic pe_1_4_clk;
    logic pe_1_4_done;
    logic [31:0] top_1_4_in;
    logic top_1_4_write_en;
    logic top_1_4_clk;
    logic [31:0] top_1_4_out;
    logic top_1_4_done;
    logic [31:0] left_1_4_in;
    logic left_1_4_write_en;
    logic left_1_4_clk;
    logic [31:0] left_1_4_out;
    logic left_1_4_done;
    logic [31:0] pe_1_5_top;
    logic [31:0] pe_1_5_left;
    logic [31:0] pe_1_5_out;
    logic pe_1_5_go;
    logic pe_1_5_clk;
    logic pe_1_5_done;
    logic [31:0] top_1_5_in;
    logic top_1_5_write_en;
    logic top_1_5_clk;
    logic [31:0] top_1_5_out;
    logic top_1_5_done;
    logic [31:0] left_1_5_in;
    logic left_1_5_write_en;
    logic left_1_5_clk;
    logic [31:0] left_1_5_out;
    logic left_1_5_done;
    logic [31:0] pe_1_6_top;
    logic [31:0] pe_1_6_left;
    logic [31:0] pe_1_6_out;
    logic pe_1_6_go;
    logic pe_1_6_clk;
    logic pe_1_6_done;
    logic [31:0] top_1_6_in;
    logic top_1_6_write_en;
    logic top_1_6_clk;
    logic [31:0] top_1_6_out;
    logic top_1_6_done;
    logic [31:0] left_1_6_in;
    logic left_1_6_write_en;
    logic left_1_6_clk;
    logic [31:0] left_1_6_out;
    logic left_1_6_done;
    logic [31:0] pe_1_7_top;
    logic [31:0] pe_1_7_left;
    logic [31:0] pe_1_7_out;
    logic pe_1_7_go;
    logic pe_1_7_clk;
    logic pe_1_7_done;
    logic [31:0] top_1_7_in;
    logic top_1_7_write_en;
    logic top_1_7_clk;
    logic [31:0] top_1_7_out;
    logic top_1_7_done;
    logic [31:0] left_1_7_in;
    logic left_1_7_write_en;
    logic left_1_7_clk;
    logic [31:0] left_1_7_out;
    logic left_1_7_done;
    logic [31:0] pe_2_0_top;
    logic [31:0] pe_2_0_left;
    logic [31:0] pe_2_0_out;
    logic pe_2_0_go;
    logic pe_2_0_clk;
    logic pe_2_0_done;
    logic [31:0] top_2_0_in;
    logic top_2_0_write_en;
    logic top_2_0_clk;
    logic [31:0] top_2_0_out;
    logic top_2_0_done;
    logic [31:0] left_2_0_in;
    logic left_2_0_write_en;
    logic left_2_0_clk;
    logic [31:0] left_2_0_out;
    logic left_2_0_done;
    logic [31:0] pe_2_1_top;
    logic [31:0] pe_2_1_left;
    logic [31:0] pe_2_1_out;
    logic pe_2_1_go;
    logic pe_2_1_clk;
    logic pe_2_1_done;
    logic [31:0] top_2_1_in;
    logic top_2_1_write_en;
    logic top_2_1_clk;
    logic [31:0] top_2_1_out;
    logic top_2_1_done;
    logic [31:0] left_2_1_in;
    logic left_2_1_write_en;
    logic left_2_1_clk;
    logic [31:0] left_2_1_out;
    logic left_2_1_done;
    logic [31:0] pe_2_2_top;
    logic [31:0] pe_2_2_left;
    logic [31:0] pe_2_2_out;
    logic pe_2_2_go;
    logic pe_2_2_clk;
    logic pe_2_2_done;
    logic [31:0] top_2_2_in;
    logic top_2_2_write_en;
    logic top_2_2_clk;
    logic [31:0] top_2_2_out;
    logic top_2_2_done;
    logic [31:0] left_2_2_in;
    logic left_2_2_write_en;
    logic left_2_2_clk;
    logic [31:0] left_2_2_out;
    logic left_2_2_done;
    logic [31:0] pe_2_3_top;
    logic [31:0] pe_2_3_left;
    logic [31:0] pe_2_3_out;
    logic pe_2_3_go;
    logic pe_2_3_clk;
    logic pe_2_3_done;
    logic [31:0] top_2_3_in;
    logic top_2_3_write_en;
    logic top_2_3_clk;
    logic [31:0] top_2_3_out;
    logic top_2_3_done;
    logic [31:0] left_2_3_in;
    logic left_2_3_write_en;
    logic left_2_3_clk;
    logic [31:0] left_2_3_out;
    logic left_2_3_done;
    logic [31:0] pe_2_4_top;
    logic [31:0] pe_2_4_left;
    logic [31:0] pe_2_4_out;
    logic pe_2_4_go;
    logic pe_2_4_clk;
    logic pe_2_4_done;
    logic [31:0] top_2_4_in;
    logic top_2_4_write_en;
    logic top_2_4_clk;
    logic [31:0] top_2_4_out;
    logic top_2_4_done;
    logic [31:0] left_2_4_in;
    logic left_2_4_write_en;
    logic left_2_4_clk;
    logic [31:0] left_2_4_out;
    logic left_2_4_done;
    logic [31:0] pe_2_5_top;
    logic [31:0] pe_2_5_left;
    logic [31:0] pe_2_5_out;
    logic pe_2_5_go;
    logic pe_2_5_clk;
    logic pe_2_5_done;
    logic [31:0] top_2_5_in;
    logic top_2_5_write_en;
    logic top_2_5_clk;
    logic [31:0] top_2_5_out;
    logic top_2_5_done;
    logic [31:0] left_2_5_in;
    logic left_2_5_write_en;
    logic left_2_5_clk;
    logic [31:0] left_2_5_out;
    logic left_2_5_done;
    logic [31:0] pe_2_6_top;
    logic [31:0] pe_2_6_left;
    logic [31:0] pe_2_6_out;
    logic pe_2_6_go;
    logic pe_2_6_clk;
    logic pe_2_6_done;
    logic [31:0] top_2_6_in;
    logic top_2_6_write_en;
    logic top_2_6_clk;
    logic [31:0] top_2_6_out;
    logic top_2_6_done;
    logic [31:0] left_2_6_in;
    logic left_2_6_write_en;
    logic left_2_6_clk;
    logic [31:0] left_2_6_out;
    logic left_2_6_done;
    logic [31:0] pe_2_7_top;
    logic [31:0] pe_2_7_left;
    logic [31:0] pe_2_7_out;
    logic pe_2_7_go;
    logic pe_2_7_clk;
    logic pe_2_7_done;
    logic [31:0] top_2_7_in;
    logic top_2_7_write_en;
    logic top_2_7_clk;
    logic [31:0] top_2_7_out;
    logic top_2_7_done;
    logic [31:0] left_2_7_in;
    logic left_2_7_write_en;
    logic left_2_7_clk;
    logic [31:0] left_2_7_out;
    logic left_2_7_done;
    logic [31:0] pe_3_0_top;
    logic [31:0] pe_3_0_left;
    logic [31:0] pe_3_0_out;
    logic pe_3_0_go;
    logic pe_3_0_clk;
    logic pe_3_0_done;
    logic [31:0] top_3_0_in;
    logic top_3_0_write_en;
    logic top_3_0_clk;
    logic [31:0] top_3_0_out;
    logic top_3_0_done;
    logic [31:0] left_3_0_in;
    logic left_3_0_write_en;
    logic left_3_0_clk;
    logic [31:0] left_3_0_out;
    logic left_3_0_done;
    logic [31:0] pe_3_1_top;
    logic [31:0] pe_3_1_left;
    logic [31:0] pe_3_1_out;
    logic pe_3_1_go;
    logic pe_3_1_clk;
    logic pe_3_1_done;
    logic [31:0] top_3_1_in;
    logic top_3_1_write_en;
    logic top_3_1_clk;
    logic [31:0] top_3_1_out;
    logic top_3_1_done;
    logic [31:0] left_3_1_in;
    logic left_3_1_write_en;
    logic left_3_1_clk;
    logic [31:0] left_3_1_out;
    logic left_3_1_done;
    logic [31:0] pe_3_2_top;
    logic [31:0] pe_3_2_left;
    logic [31:0] pe_3_2_out;
    logic pe_3_2_go;
    logic pe_3_2_clk;
    logic pe_3_2_done;
    logic [31:0] top_3_2_in;
    logic top_3_2_write_en;
    logic top_3_2_clk;
    logic [31:0] top_3_2_out;
    logic top_3_2_done;
    logic [31:0] left_3_2_in;
    logic left_3_2_write_en;
    logic left_3_2_clk;
    logic [31:0] left_3_2_out;
    logic left_3_2_done;
    logic [31:0] pe_3_3_top;
    logic [31:0] pe_3_3_left;
    logic [31:0] pe_3_3_out;
    logic pe_3_3_go;
    logic pe_3_3_clk;
    logic pe_3_3_done;
    logic [31:0] top_3_3_in;
    logic top_3_3_write_en;
    logic top_3_3_clk;
    logic [31:0] top_3_3_out;
    logic top_3_3_done;
    logic [31:0] left_3_3_in;
    logic left_3_3_write_en;
    logic left_3_3_clk;
    logic [31:0] left_3_3_out;
    logic left_3_3_done;
    logic [31:0] pe_3_4_top;
    logic [31:0] pe_3_4_left;
    logic [31:0] pe_3_4_out;
    logic pe_3_4_go;
    logic pe_3_4_clk;
    logic pe_3_4_done;
    logic [31:0] top_3_4_in;
    logic top_3_4_write_en;
    logic top_3_4_clk;
    logic [31:0] top_3_4_out;
    logic top_3_4_done;
    logic [31:0] left_3_4_in;
    logic left_3_4_write_en;
    logic left_3_4_clk;
    logic [31:0] left_3_4_out;
    logic left_3_4_done;
    logic [31:0] pe_3_5_top;
    logic [31:0] pe_3_5_left;
    logic [31:0] pe_3_5_out;
    logic pe_3_5_go;
    logic pe_3_5_clk;
    logic pe_3_5_done;
    logic [31:0] top_3_5_in;
    logic top_3_5_write_en;
    logic top_3_5_clk;
    logic [31:0] top_3_5_out;
    logic top_3_5_done;
    logic [31:0] left_3_5_in;
    logic left_3_5_write_en;
    logic left_3_5_clk;
    logic [31:0] left_3_5_out;
    logic left_3_5_done;
    logic [31:0] pe_3_6_top;
    logic [31:0] pe_3_6_left;
    logic [31:0] pe_3_6_out;
    logic pe_3_6_go;
    logic pe_3_6_clk;
    logic pe_3_6_done;
    logic [31:0] top_3_6_in;
    logic top_3_6_write_en;
    logic top_3_6_clk;
    logic [31:0] top_3_6_out;
    logic top_3_6_done;
    logic [31:0] left_3_6_in;
    logic left_3_6_write_en;
    logic left_3_6_clk;
    logic [31:0] left_3_6_out;
    logic left_3_6_done;
    logic [31:0] pe_3_7_top;
    logic [31:0] pe_3_7_left;
    logic [31:0] pe_3_7_out;
    logic pe_3_7_go;
    logic pe_3_7_clk;
    logic pe_3_7_done;
    logic [31:0] top_3_7_in;
    logic top_3_7_write_en;
    logic top_3_7_clk;
    logic [31:0] top_3_7_out;
    logic top_3_7_done;
    logic [31:0] left_3_7_in;
    logic left_3_7_write_en;
    logic left_3_7_clk;
    logic [31:0] left_3_7_out;
    logic left_3_7_done;
    logic [31:0] pe_4_0_top;
    logic [31:0] pe_4_0_left;
    logic [31:0] pe_4_0_out;
    logic pe_4_0_go;
    logic pe_4_0_clk;
    logic pe_4_0_done;
    logic [31:0] top_4_0_in;
    logic top_4_0_write_en;
    logic top_4_0_clk;
    logic [31:0] top_4_0_out;
    logic top_4_0_done;
    logic [31:0] left_4_0_in;
    logic left_4_0_write_en;
    logic left_4_0_clk;
    logic [31:0] left_4_0_out;
    logic left_4_0_done;
    logic [31:0] pe_4_1_top;
    logic [31:0] pe_4_1_left;
    logic [31:0] pe_4_1_out;
    logic pe_4_1_go;
    logic pe_4_1_clk;
    logic pe_4_1_done;
    logic [31:0] top_4_1_in;
    logic top_4_1_write_en;
    logic top_4_1_clk;
    logic [31:0] top_4_1_out;
    logic top_4_1_done;
    logic [31:0] left_4_1_in;
    logic left_4_1_write_en;
    logic left_4_1_clk;
    logic [31:0] left_4_1_out;
    logic left_4_1_done;
    logic [31:0] pe_4_2_top;
    logic [31:0] pe_4_2_left;
    logic [31:0] pe_4_2_out;
    logic pe_4_2_go;
    logic pe_4_2_clk;
    logic pe_4_2_done;
    logic [31:0] top_4_2_in;
    logic top_4_2_write_en;
    logic top_4_2_clk;
    logic [31:0] top_4_2_out;
    logic top_4_2_done;
    logic [31:0] left_4_2_in;
    logic left_4_2_write_en;
    logic left_4_2_clk;
    logic [31:0] left_4_2_out;
    logic left_4_2_done;
    logic [31:0] pe_4_3_top;
    logic [31:0] pe_4_3_left;
    logic [31:0] pe_4_3_out;
    logic pe_4_3_go;
    logic pe_4_3_clk;
    logic pe_4_3_done;
    logic [31:0] top_4_3_in;
    logic top_4_3_write_en;
    logic top_4_3_clk;
    logic [31:0] top_4_3_out;
    logic top_4_3_done;
    logic [31:0] left_4_3_in;
    logic left_4_3_write_en;
    logic left_4_3_clk;
    logic [31:0] left_4_3_out;
    logic left_4_3_done;
    logic [31:0] pe_4_4_top;
    logic [31:0] pe_4_4_left;
    logic [31:0] pe_4_4_out;
    logic pe_4_4_go;
    logic pe_4_4_clk;
    logic pe_4_4_done;
    logic [31:0] top_4_4_in;
    logic top_4_4_write_en;
    logic top_4_4_clk;
    logic [31:0] top_4_4_out;
    logic top_4_4_done;
    logic [31:0] left_4_4_in;
    logic left_4_4_write_en;
    logic left_4_4_clk;
    logic [31:0] left_4_4_out;
    logic left_4_4_done;
    logic [31:0] pe_4_5_top;
    logic [31:0] pe_4_5_left;
    logic [31:0] pe_4_5_out;
    logic pe_4_5_go;
    logic pe_4_5_clk;
    logic pe_4_5_done;
    logic [31:0] top_4_5_in;
    logic top_4_5_write_en;
    logic top_4_5_clk;
    logic [31:0] top_4_5_out;
    logic top_4_5_done;
    logic [31:0] left_4_5_in;
    logic left_4_5_write_en;
    logic left_4_5_clk;
    logic [31:0] left_4_5_out;
    logic left_4_5_done;
    logic [31:0] pe_4_6_top;
    logic [31:0] pe_4_6_left;
    logic [31:0] pe_4_6_out;
    logic pe_4_6_go;
    logic pe_4_6_clk;
    logic pe_4_6_done;
    logic [31:0] top_4_6_in;
    logic top_4_6_write_en;
    logic top_4_6_clk;
    logic [31:0] top_4_6_out;
    logic top_4_6_done;
    logic [31:0] left_4_6_in;
    logic left_4_6_write_en;
    logic left_4_6_clk;
    logic [31:0] left_4_6_out;
    logic left_4_6_done;
    logic [31:0] pe_4_7_top;
    logic [31:0] pe_4_7_left;
    logic [31:0] pe_4_7_out;
    logic pe_4_7_go;
    logic pe_4_7_clk;
    logic pe_4_7_done;
    logic [31:0] top_4_7_in;
    logic top_4_7_write_en;
    logic top_4_7_clk;
    logic [31:0] top_4_7_out;
    logic top_4_7_done;
    logic [31:0] left_4_7_in;
    logic left_4_7_write_en;
    logic left_4_7_clk;
    logic [31:0] left_4_7_out;
    logic left_4_7_done;
    logic [31:0] pe_5_0_top;
    logic [31:0] pe_5_0_left;
    logic [31:0] pe_5_0_out;
    logic pe_5_0_go;
    logic pe_5_0_clk;
    logic pe_5_0_done;
    logic [31:0] top_5_0_in;
    logic top_5_0_write_en;
    logic top_5_0_clk;
    logic [31:0] top_5_0_out;
    logic top_5_0_done;
    logic [31:0] left_5_0_in;
    logic left_5_0_write_en;
    logic left_5_0_clk;
    logic [31:0] left_5_0_out;
    logic left_5_0_done;
    logic [31:0] pe_5_1_top;
    logic [31:0] pe_5_1_left;
    logic [31:0] pe_5_1_out;
    logic pe_5_1_go;
    logic pe_5_1_clk;
    logic pe_5_1_done;
    logic [31:0] top_5_1_in;
    logic top_5_1_write_en;
    logic top_5_1_clk;
    logic [31:0] top_5_1_out;
    logic top_5_1_done;
    logic [31:0] left_5_1_in;
    logic left_5_1_write_en;
    logic left_5_1_clk;
    logic [31:0] left_5_1_out;
    logic left_5_1_done;
    logic [31:0] pe_5_2_top;
    logic [31:0] pe_5_2_left;
    logic [31:0] pe_5_2_out;
    logic pe_5_2_go;
    logic pe_5_2_clk;
    logic pe_5_2_done;
    logic [31:0] top_5_2_in;
    logic top_5_2_write_en;
    logic top_5_2_clk;
    logic [31:0] top_5_2_out;
    logic top_5_2_done;
    logic [31:0] left_5_2_in;
    logic left_5_2_write_en;
    logic left_5_2_clk;
    logic [31:0] left_5_2_out;
    logic left_5_2_done;
    logic [31:0] pe_5_3_top;
    logic [31:0] pe_5_3_left;
    logic [31:0] pe_5_3_out;
    logic pe_5_3_go;
    logic pe_5_3_clk;
    logic pe_5_3_done;
    logic [31:0] top_5_3_in;
    logic top_5_3_write_en;
    logic top_5_3_clk;
    logic [31:0] top_5_3_out;
    logic top_5_3_done;
    logic [31:0] left_5_3_in;
    logic left_5_3_write_en;
    logic left_5_3_clk;
    logic [31:0] left_5_3_out;
    logic left_5_3_done;
    logic [31:0] pe_5_4_top;
    logic [31:0] pe_5_4_left;
    logic [31:0] pe_5_4_out;
    logic pe_5_4_go;
    logic pe_5_4_clk;
    logic pe_5_4_done;
    logic [31:0] top_5_4_in;
    logic top_5_4_write_en;
    logic top_5_4_clk;
    logic [31:0] top_5_4_out;
    logic top_5_4_done;
    logic [31:0] left_5_4_in;
    logic left_5_4_write_en;
    logic left_5_4_clk;
    logic [31:0] left_5_4_out;
    logic left_5_4_done;
    logic [31:0] pe_5_5_top;
    logic [31:0] pe_5_5_left;
    logic [31:0] pe_5_5_out;
    logic pe_5_5_go;
    logic pe_5_5_clk;
    logic pe_5_5_done;
    logic [31:0] top_5_5_in;
    logic top_5_5_write_en;
    logic top_5_5_clk;
    logic [31:0] top_5_5_out;
    logic top_5_5_done;
    logic [31:0] left_5_5_in;
    logic left_5_5_write_en;
    logic left_5_5_clk;
    logic [31:0] left_5_5_out;
    logic left_5_5_done;
    logic [31:0] pe_5_6_top;
    logic [31:0] pe_5_6_left;
    logic [31:0] pe_5_6_out;
    logic pe_5_6_go;
    logic pe_5_6_clk;
    logic pe_5_6_done;
    logic [31:0] top_5_6_in;
    logic top_5_6_write_en;
    logic top_5_6_clk;
    logic [31:0] top_5_6_out;
    logic top_5_6_done;
    logic [31:0] left_5_6_in;
    logic left_5_6_write_en;
    logic left_5_6_clk;
    logic [31:0] left_5_6_out;
    logic left_5_6_done;
    logic [31:0] pe_5_7_top;
    logic [31:0] pe_5_7_left;
    logic [31:0] pe_5_7_out;
    logic pe_5_7_go;
    logic pe_5_7_clk;
    logic pe_5_7_done;
    logic [31:0] top_5_7_in;
    logic top_5_7_write_en;
    logic top_5_7_clk;
    logic [31:0] top_5_7_out;
    logic top_5_7_done;
    logic [31:0] left_5_7_in;
    logic left_5_7_write_en;
    logic left_5_7_clk;
    logic [31:0] left_5_7_out;
    logic left_5_7_done;
    logic [31:0] pe_6_0_top;
    logic [31:0] pe_6_0_left;
    logic [31:0] pe_6_0_out;
    logic pe_6_0_go;
    logic pe_6_0_clk;
    logic pe_6_0_done;
    logic [31:0] top_6_0_in;
    logic top_6_0_write_en;
    logic top_6_0_clk;
    logic [31:0] top_6_0_out;
    logic top_6_0_done;
    logic [31:0] left_6_0_in;
    logic left_6_0_write_en;
    logic left_6_0_clk;
    logic [31:0] left_6_0_out;
    logic left_6_0_done;
    logic [31:0] pe_6_1_top;
    logic [31:0] pe_6_1_left;
    logic [31:0] pe_6_1_out;
    logic pe_6_1_go;
    logic pe_6_1_clk;
    logic pe_6_1_done;
    logic [31:0] top_6_1_in;
    logic top_6_1_write_en;
    logic top_6_1_clk;
    logic [31:0] top_6_1_out;
    logic top_6_1_done;
    logic [31:0] left_6_1_in;
    logic left_6_1_write_en;
    logic left_6_1_clk;
    logic [31:0] left_6_1_out;
    logic left_6_1_done;
    logic [31:0] pe_6_2_top;
    logic [31:0] pe_6_2_left;
    logic [31:0] pe_6_2_out;
    logic pe_6_2_go;
    logic pe_6_2_clk;
    logic pe_6_2_done;
    logic [31:0] top_6_2_in;
    logic top_6_2_write_en;
    logic top_6_2_clk;
    logic [31:0] top_6_2_out;
    logic top_6_2_done;
    logic [31:0] left_6_2_in;
    logic left_6_2_write_en;
    logic left_6_2_clk;
    logic [31:0] left_6_2_out;
    logic left_6_2_done;
    logic [31:0] pe_6_3_top;
    logic [31:0] pe_6_3_left;
    logic [31:0] pe_6_3_out;
    logic pe_6_3_go;
    logic pe_6_3_clk;
    logic pe_6_3_done;
    logic [31:0] top_6_3_in;
    logic top_6_3_write_en;
    logic top_6_3_clk;
    logic [31:0] top_6_3_out;
    logic top_6_3_done;
    logic [31:0] left_6_3_in;
    logic left_6_3_write_en;
    logic left_6_3_clk;
    logic [31:0] left_6_3_out;
    logic left_6_3_done;
    logic [31:0] pe_6_4_top;
    logic [31:0] pe_6_4_left;
    logic [31:0] pe_6_4_out;
    logic pe_6_4_go;
    logic pe_6_4_clk;
    logic pe_6_4_done;
    logic [31:0] top_6_4_in;
    logic top_6_4_write_en;
    logic top_6_4_clk;
    logic [31:0] top_6_4_out;
    logic top_6_4_done;
    logic [31:0] left_6_4_in;
    logic left_6_4_write_en;
    logic left_6_4_clk;
    logic [31:0] left_6_4_out;
    logic left_6_4_done;
    logic [31:0] pe_6_5_top;
    logic [31:0] pe_6_5_left;
    logic [31:0] pe_6_5_out;
    logic pe_6_5_go;
    logic pe_6_5_clk;
    logic pe_6_5_done;
    logic [31:0] top_6_5_in;
    logic top_6_5_write_en;
    logic top_6_5_clk;
    logic [31:0] top_6_5_out;
    logic top_6_5_done;
    logic [31:0] left_6_5_in;
    logic left_6_5_write_en;
    logic left_6_5_clk;
    logic [31:0] left_6_5_out;
    logic left_6_5_done;
    logic [31:0] pe_6_6_top;
    logic [31:0] pe_6_6_left;
    logic [31:0] pe_6_6_out;
    logic pe_6_6_go;
    logic pe_6_6_clk;
    logic pe_6_6_done;
    logic [31:0] top_6_6_in;
    logic top_6_6_write_en;
    logic top_6_6_clk;
    logic [31:0] top_6_6_out;
    logic top_6_6_done;
    logic [31:0] left_6_6_in;
    logic left_6_6_write_en;
    logic left_6_6_clk;
    logic [31:0] left_6_6_out;
    logic left_6_6_done;
    logic [31:0] pe_6_7_top;
    logic [31:0] pe_6_7_left;
    logic [31:0] pe_6_7_out;
    logic pe_6_7_go;
    logic pe_6_7_clk;
    logic pe_6_7_done;
    logic [31:0] top_6_7_in;
    logic top_6_7_write_en;
    logic top_6_7_clk;
    logic [31:0] top_6_7_out;
    logic top_6_7_done;
    logic [31:0] left_6_7_in;
    logic left_6_7_write_en;
    logic left_6_7_clk;
    logic [31:0] left_6_7_out;
    logic left_6_7_done;
    logic [31:0] pe_7_0_top;
    logic [31:0] pe_7_0_left;
    logic [31:0] pe_7_0_out;
    logic pe_7_0_go;
    logic pe_7_0_clk;
    logic pe_7_0_done;
    logic [31:0] top_7_0_in;
    logic top_7_0_write_en;
    logic top_7_0_clk;
    logic [31:0] top_7_0_out;
    logic top_7_0_done;
    logic [31:0] left_7_0_in;
    logic left_7_0_write_en;
    logic left_7_0_clk;
    logic [31:0] left_7_0_out;
    logic left_7_0_done;
    logic [31:0] pe_7_1_top;
    logic [31:0] pe_7_1_left;
    logic [31:0] pe_7_1_out;
    logic pe_7_1_go;
    logic pe_7_1_clk;
    logic pe_7_1_done;
    logic [31:0] top_7_1_in;
    logic top_7_1_write_en;
    logic top_7_1_clk;
    logic [31:0] top_7_1_out;
    logic top_7_1_done;
    logic [31:0] left_7_1_in;
    logic left_7_1_write_en;
    logic left_7_1_clk;
    logic [31:0] left_7_1_out;
    logic left_7_1_done;
    logic [31:0] pe_7_2_top;
    logic [31:0] pe_7_2_left;
    logic [31:0] pe_7_2_out;
    logic pe_7_2_go;
    logic pe_7_2_clk;
    logic pe_7_2_done;
    logic [31:0] top_7_2_in;
    logic top_7_2_write_en;
    logic top_7_2_clk;
    logic [31:0] top_7_2_out;
    logic top_7_2_done;
    logic [31:0] left_7_2_in;
    logic left_7_2_write_en;
    logic left_7_2_clk;
    logic [31:0] left_7_2_out;
    logic left_7_2_done;
    logic [31:0] pe_7_3_top;
    logic [31:0] pe_7_3_left;
    logic [31:0] pe_7_3_out;
    logic pe_7_3_go;
    logic pe_7_3_clk;
    logic pe_7_3_done;
    logic [31:0] top_7_3_in;
    logic top_7_3_write_en;
    logic top_7_3_clk;
    logic [31:0] top_7_3_out;
    logic top_7_3_done;
    logic [31:0] left_7_3_in;
    logic left_7_3_write_en;
    logic left_7_3_clk;
    logic [31:0] left_7_3_out;
    logic left_7_3_done;
    logic [31:0] pe_7_4_top;
    logic [31:0] pe_7_4_left;
    logic [31:0] pe_7_4_out;
    logic pe_7_4_go;
    logic pe_7_4_clk;
    logic pe_7_4_done;
    logic [31:0] top_7_4_in;
    logic top_7_4_write_en;
    logic top_7_4_clk;
    logic [31:0] top_7_4_out;
    logic top_7_4_done;
    logic [31:0] left_7_4_in;
    logic left_7_4_write_en;
    logic left_7_4_clk;
    logic [31:0] left_7_4_out;
    logic left_7_4_done;
    logic [31:0] pe_7_5_top;
    logic [31:0] pe_7_5_left;
    logic [31:0] pe_7_5_out;
    logic pe_7_5_go;
    logic pe_7_5_clk;
    logic pe_7_5_done;
    logic [31:0] top_7_5_in;
    logic top_7_5_write_en;
    logic top_7_5_clk;
    logic [31:0] top_7_5_out;
    logic top_7_5_done;
    logic [31:0] left_7_5_in;
    logic left_7_5_write_en;
    logic left_7_5_clk;
    logic [31:0] left_7_5_out;
    logic left_7_5_done;
    logic [31:0] pe_7_6_top;
    logic [31:0] pe_7_6_left;
    logic [31:0] pe_7_6_out;
    logic pe_7_6_go;
    logic pe_7_6_clk;
    logic pe_7_6_done;
    logic [31:0] top_7_6_in;
    logic top_7_6_write_en;
    logic top_7_6_clk;
    logic [31:0] top_7_6_out;
    logic top_7_6_done;
    logic [31:0] left_7_6_in;
    logic left_7_6_write_en;
    logic left_7_6_clk;
    logic [31:0] left_7_6_out;
    logic left_7_6_done;
    logic [31:0] pe_7_7_top;
    logic [31:0] pe_7_7_left;
    logic [31:0] pe_7_7_out;
    logic pe_7_7_go;
    logic pe_7_7_clk;
    logic pe_7_7_done;
    logic [31:0] top_7_7_in;
    logic top_7_7_write_en;
    logic top_7_7_clk;
    logic [31:0] top_7_7_out;
    logic top_7_7_done;
    logic [31:0] left_7_7_in;
    logic left_7_7_write_en;
    logic left_7_7_clk;
    logic [31:0] left_7_7_out;
    logic left_7_7_done;
    logic fsm_in;
    logic fsm_write_en;
    logic fsm_clk;
    logic fsm_out;
    logic fsm_done;
    logic incr_left;
    logic incr_right;
    logic incr_out;
    logic fsm0_in;
    logic fsm0_write_en;
    logic fsm0_clk;
    logic fsm0_out;
    logic fsm0_done;
    logic incr0_left;
    logic incr0_right;
    logic incr0_out;
    logic fsm1_in;
    logic fsm1_write_en;
    logic fsm1_clk;
    logic fsm1_out;
    logic fsm1_done;
    logic incr1_left;
    logic incr1_right;
    logic incr1_out;
    logic [2:0] fsm2_in;
    logic fsm2_write_en;
    logic fsm2_clk;
    logic [2:0] fsm2_out;
    logic fsm2_done;
    logic [2:0] incr2_left;
    logic [2:0] incr2_right;
    logic [2:0] incr2_out;
    logic fsm3_in;
    logic fsm3_write_en;
    logic fsm3_clk;
    logic fsm3_out;
    logic fsm3_done;
    logic incr3_left;
    logic incr3_right;
    logic incr3_out;
    logic [2:0] fsm4_in;
    logic fsm4_write_en;
    logic fsm4_clk;
    logic [2:0] fsm4_out;
    logic fsm4_done;
    logic [2:0] incr4_left;
    logic [2:0] incr4_right;
    logic [2:0] incr4_out;
    logic fsm5_in;
    logic fsm5_write_en;
    logic fsm5_clk;
    logic fsm5_out;
    logic fsm5_done;
    logic incr5_left;
    logic incr5_right;
    logic incr5_out;
    logic [2:0] fsm6_in;
    logic fsm6_write_en;
    logic fsm6_clk;
    logic [2:0] fsm6_out;
    logic fsm6_done;
    logic [2:0] incr6_left;
    logic [2:0] incr6_right;
    logic [2:0] incr6_out;
    logic fsm7_in;
    logic fsm7_write_en;
    logic fsm7_clk;
    logic fsm7_out;
    logic fsm7_done;
    logic incr7_left;
    logic incr7_right;
    logic incr7_out;
    logic [2:0] fsm8_in;
    logic fsm8_write_en;
    logic fsm8_clk;
    logic [2:0] fsm8_out;
    logic fsm8_done;
    logic [2:0] incr8_left;
    logic [2:0] incr8_right;
    logic [2:0] incr8_out;
    logic fsm9_in;
    logic fsm9_write_en;
    logic fsm9_clk;
    logic fsm9_out;
    logic fsm9_done;
    logic incr9_left;
    logic incr9_right;
    logic incr9_out;
    logic [2:0] fsm10_in;
    logic fsm10_write_en;
    logic fsm10_clk;
    logic [2:0] fsm10_out;
    logic fsm10_done;
    logic [2:0] incr10_left;
    logic [2:0] incr10_right;
    logic [2:0] incr10_out;
    logic fsm11_in;
    logic fsm11_write_en;
    logic fsm11_clk;
    logic fsm11_out;
    logic fsm11_done;
    logic incr11_left;
    logic incr11_right;
    logic incr11_out;
    logic [2:0] fsm12_in;
    logic fsm12_write_en;
    logic fsm12_clk;
    logic [2:0] fsm12_out;
    logic fsm12_done;
    logic [2:0] incr12_left;
    logic [2:0] incr12_right;
    logic [2:0] incr12_out;
    logic fsm13_in;
    logic fsm13_write_en;
    logic fsm13_clk;
    logic fsm13_out;
    logic fsm13_done;
    logic incr13_left;
    logic incr13_right;
    logic incr13_out;
    logic [2:0] fsm14_in;
    logic fsm14_write_en;
    logic fsm14_clk;
    logic [2:0] fsm14_out;
    logic fsm14_done;
    logic [2:0] incr14_left;
    logic [2:0] incr14_right;
    logic [2:0] incr14_out;
    logic fsm15_in;
    logic fsm15_write_en;
    logic fsm15_clk;
    logic fsm15_out;
    logic fsm15_done;
    logic incr15_left;
    logic incr15_right;
    logic incr15_out;
    logic [2:0] fsm16_in;
    logic fsm16_write_en;
    logic fsm16_clk;
    logic [2:0] fsm16_out;
    logic fsm16_done;
    logic [2:0] incr16_left;
    logic [2:0] incr16_right;
    logic [2:0] incr16_out;
    logic fsm17_in;
    logic fsm17_write_en;
    logic fsm17_clk;
    logic fsm17_out;
    logic fsm17_done;
    logic incr17_left;
    logic incr17_right;
    logic incr17_out;
    logic [2:0] fsm18_in;
    logic fsm18_write_en;
    logic fsm18_clk;
    logic [2:0] fsm18_out;
    logic fsm18_done;
    logic [2:0] incr18_left;
    logic [2:0] incr18_right;
    logic [2:0] incr18_out;
    logic fsm19_in;
    logic fsm19_write_en;
    logic fsm19_clk;
    logic fsm19_out;
    logic fsm19_done;
    logic incr19_left;
    logic incr19_right;
    logic incr19_out;
    logic [2:0] fsm20_in;
    logic fsm20_write_en;
    logic fsm20_clk;
    logic [2:0] fsm20_out;
    logic fsm20_done;
    logic [2:0] incr20_left;
    logic [2:0] incr20_right;
    logic [2:0] incr20_out;
    logic fsm21_in;
    logic fsm21_write_en;
    logic fsm21_clk;
    logic fsm21_out;
    logic fsm21_done;
    logic incr21_left;
    logic incr21_right;
    logic incr21_out;
    logic [2:0] fsm22_in;
    logic fsm22_write_en;
    logic fsm22_clk;
    logic [2:0] fsm22_out;
    logic fsm22_done;
    logic [2:0] incr22_left;
    logic [2:0] incr22_right;
    logic [2:0] incr22_out;
    logic fsm23_in;
    logic fsm23_write_en;
    logic fsm23_clk;
    logic fsm23_out;
    logic fsm23_done;
    logic incr23_left;
    logic incr23_right;
    logic incr23_out;
    logic [2:0] fsm24_in;
    logic fsm24_write_en;
    logic fsm24_clk;
    logic [2:0] fsm24_out;
    logic fsm24_done;
    logic [2:0] incr24_left;
    logic [2:0] incr24_right;
    logic [2:0] incr24_out;
    logic fsm25_in;
    logic fsm25_write_en;
    logic fsm25_clk;
    logic fsm25_out;
    logic fsm25_done;
    logic incr25_left;
    logic incr25_right;
    logic incr25_out;
    logic [2:0] fsm26_in;
    logic fsm26_write_en;
    logic fsm26_clk;
    logic [2:0] fsm26_out;
    logic fsm26_done;
    logic [2:0] incr26_left;
    logic [2:0] incr26_right;
    logic [2:0] incr26_out;
    logic fsm27_in;
    logic fsm27_write_en;
    logic fsm27_clk;
    logic fsm27_out;
    logic fsm27_done;
    logic incr27_left;
    logic incr27_right;
    logic incr27_out;
    logic [2:0] fsm28_in;
    logic fsm28_write_en;
    logic fsm28_clk;
    logic [2:0] fsm28_out;
    logic fsm28_done;
    logic [2:0] incr28_left;
    logic [2:0] incr28_right;
    logic [2:0] incr28_out;
    logic fsm29_in;
    logic fsm29_write_en;
    logic fsm29_clk;
    logic fsm29_out;
    logic fsm29_done;
    logic incr29_left;
    logic incr29_right;
    logic incr29_out;
    logic [2:0] fsm30_in;
    logic fsm30_write_en;
    logic fsm30_clk;
    logic [2:0] fsm30_out;
    logic fsm30_done;
    logic [2:0] incr30_left;
    logic [2:0] incr30_right;
    logic [2:0] incr30_out;
    logic fsm31_in;
    logic fsm31_write_en;
    logic fsm31_clk;
    logic fsm31_out;
    logic fsm31_done;
    logic incr31_left;
    logic incr31_right;
    logic incr31_out;
    logic [2:0] fsm32_in;
    logic fsm32_write_en;
    logic fsm32_clk;
    logic [2:0] fsm32_out;
    logic fsm32_done;
    logic [2:0] incr32_left;
    logic [2:0] incr32_right;
    logic [2:0] incr32_out;
    logic fsm33_in;
    logic fsm33_write_en;
    logic fsm33_clk;
    logic fsm33_out;
    logic fsm33_done;
    logic incr33_left;
    logic incr33_right;
    logic incr33_out;
    logic [2:0] fsm34_in;
    logic fsm34_write_en;
    logic fsm34_clk;
    logic [2:0] fsm34_out;
    logic fsm34_done;
    logic [2:0] incr34_left;
    logic [2:0] incr34_right;
    logic [2:0] incr34_out;
    logic fsm35_in;
    logic fsm35_write_en;
    logic fsm35_clk;
    logic fsm35_out;
    logic fsm35_done;
    logic incr35_left;
    logic incr35_right;
    logic incr35_out;
    logic [2:0] fsm36_in;
    logic fsm36_write_en;
    logic fsm36_clk;
    logic [2:0] fsm36_out;
    logic fsm36_done;
    logic [2:0] incr36_left;
    logic [2:0] incr36_right;
    logic [2:0] incr36_out;
    logic fsm37_in;
    logic fsm37_write_en;
    logic fsm37_clk;
    logic fsm37_out;
    logic fsm37_done;
    logic incr37_left;
    logic incr37_right;
    logic incr37_out;
    logic [2:0] fsm38_in;
    logic fsm38_write_en;
    logic fsm38_clk;
    logic [2:0] fsm38_out;
    logic fsm38_done;
    logic [2:0] incr38_left;
    logic [2:0] incr38_right;
    logic [2:0] incr38_out;
    logic fsm39_in;
    logic fsm39_write_en;
    logic fsm39_clk;
    logic fsm39_out;
    logic fsm39_done;
    logic incr39_left;
    logic incr39_right;
    logic incr39_out;
    logic [2:0] fsm40_in;
    logic fsm40_write_en;
    logic fsm40_clk;
    logic [2:0] fsm40_out;
    logic fsm40_done;
    logic [2:0] incr40_left;
    logic [2:0] incr40_right;
    logic [2:0] incr40_out;
    logic fsm41_in;
    logic fsm41_write_en;
    logic fsm41_clk;
    logic fsm41_out;
    logic fsm41_done;
    logic incr41_left;
    logic incr41_right;
    logic incr41_out;
    logic [2:0] fsm42_in;
    logic fsm42_write_en;
    logic fsm42_clk;
    logic [2:0] fsm42_out;
    logic fsm42_done;
    logic [2:0] incr42_left;
    logic [2:0] incr42_right;
    logic [2:0] incr42_out;
    logic fsm43_in;
    logic fsm43_write_en;
    logic fsm43_clk;
    logic fsm43_out;
    logic fsm43_done;
    logic incr43_left;
    logic incr43_right;
    logic incr43_out;
    logic [7:0] fsm44_in;
    logic fsm44_write_en;
    logic fsm44_clk;
    logic [7:0] fsm44_out;
    logic fsm44_done;
    logic [7:0] incr44_left;
    logic [7:0] incr44_right;
    logic [7:0] incr44_out;
    initial begin
        t0_idx_in = 4'd0;
        t0_idx_write_en = 1'd0;
        t0_idx_clk = 1'd0;
        t0_add_left = 4'd0;
        t0_add_right = 4'd0;
        t1_idx_in = 4'd0;
        t1_idx_write_en = 1'd0;
        t1_idx_clk = 1'd0;
        t1_add_left = 4'd0;
        t1_add_right = 4'd0;
        t2_idx_in = 4'd0;
        t2_idx_write_en = 1'd0;
        t2_idx_clk = 1'd0;
        t2_add_left = 4'd0;
        t2_add_right = 4'd0;
        t3_idx_in = 4'd0;
        t3_idx_write_en = 1'd0;
        t3_idx_clk = 1'd0;
        t3_add_left = 4'd0;
        t3_add_right = 4'd0;
        t4_idx_in = 4'd0;
        t4_idx_write_en = 1'd0;
        t4_idx_clk = 1'd0;
        t4_add_left = 4'd0;
        t4_add_right = 4'd0;
        t5_idx_in = 4'd0;
        t5_idx_write_en = 1'd0;
        t5_idx_clk = 1'd0;
        t5_add_left = 4'd0;
        t5_add_right = 4'd0;
        t6_idx_in = 4'd0;
        t6_idx_write_en = 1'd0;
        t6_idx_clk = 1'd0;
        t6_add_left = 4'd0;
        t6_add_right = 4'd0;
        t7_idx_in = 4'd0;
        t7_idx_write_en = 1'd0;
        t7_idx_clk = 1'd0;
        t7_add_left = 4'd0;
        t7_add_right = 4'd0;
        l0_idx_in = 4'd0;
        l0_idx_write_en = 1'd0;
        l0_idx_clk = 1'd0;
        l0_add_left = 4'd0;
        l0_add_right = 4'd0;
        l1_idx_in = 4'd0;
        l1_idx_write_en = 1'd0;
        l1_idx_clk = 1'd0;
        l1_add_left = 4'd0;
        l1_add_right = 4'd0;
        l2_idx_in = 4'd0;
        l2_idx_write_en = 1'd0;
        l2_idx_clk = 1'd0;
        l2_add_left = 4'd0;
        l2_add_right = 4'd0;
        l3_idx_in = 4'd0;
        l3_idx_write_en = 1'd0;
        l3_idx_clk = 1'd0;
        l3_add_left = 4'd0;
        l3_add_right = 4'd0;
        l4_idx_in = 4'd0;
        l4_idx_write_en = 1'd0;
        l4_idx_clk = 1'd0;
        l4_add_left = 4'd0;
        l4_add_right = 4'd0;
        l5_idx_in = 4'd0;
        l5_idx_write_en = 1'd0;
        l5_idx_clk = 1'd0;
        l5_add_left = 4'd0;
        l5_add_right = 4'd0;
        l6_idx_in = 4'd0;
        l6_idx_write_en = 1'd0;
        l6_idx_clk = 1'd0;
        l6_add_left = 4'd0;
        l6_add_right = 4'd0;
        l7_idx_in = 4'd0;
        l7_idx_write_en = 1'd0;
        l7_idx_clk = 1'd0;
        l7_add_left = 4'd0;
        l7_add_right = 4'd0;
        pe_0_0_top = 32'd0;
        pe_0_0_left = 32'd0;
        pe_0_0_go = 1'd0;
        pe_0_0_clk = 1'd0;
        top_0_0_in = 32'd0;
        top_0_0_write_en = 1'd0;
        top_0_0_clk = 1'd0;
        left_0_0_in = 32'd0;
        left_0_0_write_en = 1'd0;
        left_0_0_clk = 1'd0;
        pe_0_1_top = 32'd0;
        pe_0_1_left = 32'd0;
        pe_0_1_go = 1'd0;
        pe_0_1_clk = 1'd0;
        top_0_1_in = 32'd0;
        top_0_1_write_en = 1'd0;
        top_0_1_clk = 1'd0;
        left_0_1_in = 32'd0;
        left_0_1_write_en = 1'd0;
        left_0_1_clk = 1'd0;
        pe_0_2_top = 32'd0;
        pe_0_2_left = 32'd0;
        pe_0_2_go = 1'd0;
        pe_0_2_clk = 1'd0;
        top_0_2_in = 32'd0;
        top_0_2_write_en = 1'd0;
        top_0_2_clk = 1'd0;
        left_0_2_in = 32'd0;
        left_0_2_write_en = 1'd0;
        left_0_2_clk = 1'd0;
        pe_0_3_top = 32'd0;
        pe_0_3_left = 32'd0;
        pe_0_3_go = 1'd0;
        pe_0_3_clk = 1'd0;
        top_0_3_in = 32'd0;
        top_0_3_write_en = 1'd0;
        top_0_3_clk = 1'd0;
        left_0_3_in = 32'd0;
        left_0_3_write_en = 1'd0;
        left_0_3_clk = 1'd0;
        pe_0_4_top = 32'd0;
        pe_0_4_left = 32'd0;
        pe_0_4_go = 1'd0;
        pe_0_4_clk = 1'd0;
        top_0_4_in = 32'd0;
        top_0_4_write_en = 1'd0;
        top_0_4_clk = 1'd0;
        left_0_4_in = 32'd0;
        left_0_4_write_en = 1'd0;
        left_0_4_clk = 1'd0;
        pe_0_5_top = 32'd0;
        pe_0_5_left = 32'd0;
        pe_0_5_go = 1'd0;
        pe_0_5_clk = 1'd0;
        top_0_5_in = 32'd0;
        top_0_5_write_en = 1'd0;
        top_0_5_clk = 1'd0;
        left_0_5_in = 32'd0;
        left_0_5_write_en = 1'd0;
        left_0_5_clk = 1'd0;
        pe_0_6_top = 32'd0;
        pe_0_6_left = 32'd0;
        pe_0_6_go = 1'd0;
        pe_0_6_clk = 1'd0;
        top_0_6_in = 32'd0;
        top_0_6_write_en = 1'd0;
        top_0_6_clk = 1'd0;
        left_0_6_in = 32'd0;
        left_0_6_write_en = 1'd0;
        left_0_6_clk = 1'd0;
        pe_0_7_top = 32'd0;
        pe_0_7_left = 32'd0;
        pe_0_7_go = 1'd0;
        pe_0_7_clk = 1'd0;
        top_0_7_in = 32'd0;
        top_0_7_write_en = 1'd0;
        top_0_7_clk = 1'd0;
        left_0_7_in = 32'd0;
        left_0_7_write_en = 1'd0;
        left_0_7_clk = 1'd0;
        pe_1_0_top = 32'd0;
        pe_1_0_left = 32'd0;
        pe_1_0_go = 1'd0;
        pe_1_0_clk = 1'd0;
        top_1_0_in = 32'd0;
        top_1_0_write_en = 1'd0;
        top_1_0_clk = 1'd0;
        left_1_0_in = 32'd0;
        left_1_0_write_en = 1'd0;
        left_1_0_clk = 1'd0;
        pe_1_1_top = 32'd0;
        pe_1_1_left = 32'd0;
        pe_1_1_go = 1'd0;
        pe_1_1_clk = 1'd0;
        top_1_1_in = 32'd0;
        top_1_1_write_en = 1'd0;
        top_1_1_clk = 1'd0;
        left_1_1_in = 32'd0;
        left_1_1_write_en = 1'd0;
        left_1_1_clk = 1'd0;
        pe_1_2_top = 32'd0;
        pe_1_2_left = 32'd0;
        pe_1_2_go = 1'd0;
        pe_1_2_clk = 1'd0;
        top_1_2_in = 32'd0;
        top_1_2_write_en = 1'd0;
        top_1_2_clk = 1'd0;
        left_1_2_in = 32'd0;
        left_1_2_write_en = 1'd0;
        left_1_2_clk = 1'd0;
        pe_1_3_top = 32'd0;
        pe_1_3_left = 32'd0;
        pe_1_3_go = 1'd0;
        pe_1_3_clk = 1'd0;
        top_1_3_in = 32'd0;
        top_1_3_write_en = 1'd0;
        top_1_3_clk = 1'd0;
        left_1_3_in = 32'd0;
        left_1_3_write_en = 1'd0;
        left_1_3_clk = 1'd0;
        pe_1_4_top = 32'd0;
        pe_1_4_left = 32'd0;
        pe_1_4_go = 1'd0;
        pe_1_4_clk = 1'd0;
        top_1_4_in = 32'd0;
        top_1_4_write_en = 1'd0;
        top_1_4_clk = 1'd0;
        left_1_4_in = 32'd0;
        left_1_4_write_en = 1'd0;
        left_1_4_clk = 1'd0;
        pe_1_5_top = 32'd0;
        pe_1_5_left = 32'd0;
        pe_1_5_go = 1'd0;
        pe_1_5_clk = 1'd0;
        top_1_5_in = 32'd0;
        top_1_5_write_en = 1'd0;
        top_1_5_clk = 1'd0;
        left_1_5_in = 32'd0;
        left_1_5_write_en = 1'd0;
        left_1_5_clk = 1'd0;
        pe_1_6_top = 32'd0;
        pe_1_6_left = 32'd0;
        pe_1_6_go = 1'd0;
        pe_1_6_clk = 1'd0;
        top_1_6_in = 32'd0;
        top_1_6_write_en = 1'd0;
        top_1_6_clk = 1'd0;
        left_1_6_in = 32'd0;
        left_1_6_write_en = 1'd0;
        left_1_6_clk = 1'd0;
        pe_1_7_top = 32'd0;
        pe_1_7_left = 32'd0;
        pe_1_7_go = 1'd0;
        pe_1_7_clk = 1'd0;
        top_1_7_in = 32'd0;
        top_1_7_write_en = 1'd0;
        top_1_7_clk = 1'd0;
        left_1_7_in = 32'd0;
        left_1_7_write_en = 1'd0;
        left_1_7_clk = 1'd0;
        pe_2_0_top = 32'd0;
        pe_2_0_left = 32'd0;
        pe_2_0_go = 1'd0;
        pe_2_0_clk = 1'd0;
        top_2_0_in = 32'd0;
        top_2_0_write_en = 1'd0;
        top_2_0_clk = 1'd0;
        left_2_0_in = 32'd0;
        left_2_0_write_en = 1'd0;
        left_2_0_clk = 1'd0;
        pe_2_1_top = 32'd0;
        pe_2_1_left = 32'd0;
        pe_2_1_go = 1'd0;
        pe_2_1_clk = 1'd0;
        top_2_1_in = 32'd0;
        top_2_1_write_en = 1'd0;
        top_2_1_clk = 1'd0;
        left_2_1_in = 32'd0;
        left_2_1_write_en = 1'd0;
        left_2_1_clk = 1'd0;
        pe_2_2_top = 32'd0;
        pe_2_2_left = 32'd0;
        pe_2_2_go = 1'd0;
        pe_2_2_clk = 1'd0;
        top_2_2_in = 32'd0;
        top_2_2_write_en = 1'd0;
        top_2_2_clk = 1'd0;
        left_2_2_in = 32'd0;
        left_2_2_write_en = 1'd0;
        left_2_2_clk = 1'd0;
        pe_2_3_top = 32'd0;
        pe_2_3_left = 32'd0;
        pe_2_3_go = 1'd0;
        pe_2_3_clk = 1'd0;
        top_2_3_in = 32'd0;
        top_2_3_write_en = 1'd0;
        top_2_3_clk = 1'd0;
        left_2_3_in = 32'd0;
        left_2_3_write_en = 1'd0;
        left_2_3_clk = 1'd0;
        pe_2_4_top = 32'd0;
        pe_2_4_left = 32'd0;
        pe_2_4_go = 1'd0;
        pe_2_4_clk = 1'd0;
        top_2_4_in = 32'd0;
        top_2_4_write_en = 1'd0;
        top_2_4_clk = 1'd0;
        left_2_4_in = 32'd0;
        left_2_4_write_en = 1'd0;
        left_2_4_clk = 1'd0;
        pe_2_5_top = 32'd0;
        pe_2_5_left = 32'd0;
        pe_2_5_go = 1'd0;
        pe_2_5_clk = 1'd0;
        top_2_5_in = 32'd0;
        top_2_5_write_en = 1'd0;
        top_2_5_clk = 1'd0;
        left_2_5_in = 32'd0;
        left_2_5_write_en = 1'd0;
        left_2_5_clk = 1'd0;
        pe_2_6_top = 32'd0;
        pe_2_6_left = 32'd0;
        pe_2_6_go = 1'd0;
        pe_2_6_clk = 1'd0;
        top_2_6_in = 32'd0;
        top_2_6_write_en = 1'd0;
        top_2_6_clk = 1'd0;
        left_2_6_in = 32'd0;
        left_2_6_write_en = 1'd0;
        left_2_6_clk = 1'd0;
        pe_2_7_top = 32'd0;
        pe_2_7_left = 32'd0;
        pe_2_7_go = 1'd0;
        pe_2_7_clk = 1'd0;
        top_2_7_in = 32'd0;
        top_2_7_write_en = 1'd0;
        top_2_7_clk = 1'd0;
        left_2_7_in = 32'd0;
        left_2_7_write_en = 1'd0;
        left_2_7_clk = 1'd0;
        pe_3_0_top = 32'd0;
        pe_3_0_left = 32'd0;
        pe_3_0_go = 1'd0;
        pe_3_0_clk = 1'd0;
        top_3_0_in = 32'd0;
        top_3_0_write_en = 1'd0;
        top_3_0_clk = 1'd0;
        left_3_0_in = 32'd0;
        left_3_0_write_en = 1'd0;
        left_3_0_clk = 1'd0;
        pe_3_1_top = 32'd0;
        pe_3_1_left = 32'd0;
        pe_3_1_go = 1'd0;
        pe_3_1_clk = 1'd0;
        top_3_1_in = 32'd0;
        top_3_1_write_en = 1'd0;
        top_3_1_clk = 1'd0;
        left_3_1_in = 32'd0;
        left_3_1_write_en = 1'd0;
        left_3_1_clk = 1'd0;
        pe_3_2_top = 32'd0;
        pe_3_2_left = 32'd0;
        pe_3_2_go = 1'd0;
        pe_3_2_clk = 1'd0;
        top_3_2_in = 32'd0;
        top_3_2_write_en = 1'd0;
        top_3_2_clk = 1'd0;
        left_3_2_in = 32'd0;
        left_3_2_write_en = 1'd0;
        left_3_2_clk = 1'd0;
        pe_3_3_top = 32'd0;
        pe_3_3_left = 32'd0;
        pe_3_3_go = 1'd0;
        pe_3_3_clk = 1'd0;
        top_3_3_in = 32'd0;
        top_3_3_write_en = 1'd0;
        top_3_3_clk = 1'd0;
        left_3_3_in = 32'd0;
        left_3_3_write_en = 1'd0;
        left_3_3_clk = 1'd0;
        pe_3_4_top = 32'd0;
        pe_3_4_left = 32'd0;
        pe_3_4_go = 1'd0;
        pe_3_4_clk = 1'd0;
        top_3_4_in = 32'd0;
        top_3_4_write_en = 1'd0;
        top_3_4_clk = 1'd0;
        left_3_4_in = 32'd0;
        left_3_4_write_en = 1'd0;
        left_3_4_clk = 1'd0;
        pe_3_5_top = 32'd0;
        pe_3_5_left = 32'd0;
        pe_3_5_go = 1'd0;
        pe_3_5_clk = 1'd0;
        top_3_5_in = 32'd0;
        top_3_5_write_en = 1'd0;
        top_3_5_clk = 1'd0;
        left_3_5_in = 32'd0;
        left_3_5_write_en = 1'd0;
        left_3_5_clk = 1'd0;
        pe_3_6_top = 32'd0;
        pe_3_6_left = 32'd0;
        pe_3_6_go = 1'd0;
        pe_3_6_clk = 1'd0;
        top_3_6_in = 32'd0;
        top_3_6_write_en = 1'd0;
        top_3_6_clk = 1'd0;
        left_3_6_in = 32'd0;
        left_3_6_write_en = 1'd0;
        left_3_6_clk = 1'd0;
        pe_3_7_top = 32'd0;
        pe_3_7_left = 32'd0;
        pe_3_7_go = 1'd0;
        pe_3_7_clk = 1'd0;
        top_3_7_in = 32'd0;
        top_3_7_write_en = 1'd0;
        top_3_7_clk = 1'd0;
        left_3_7_in = 32'd0;
        left_3_7_write_en = 1'd0;
        left_3_7_clk = 1'd0;
        pe_4_0_top = 32'd0;
        pe_4_0_left = 32'd0;
        pe_4_0_go = 1'd0;
        pe_4_0_clk = 1'd0;
        top_4_0_in = 32'd0;
        top_4_0_write_en = 1'd0;
        top_4_0_clk = 1'd0;
        left_4_0_in = 32'd0;
        left_4_0_write_en = 1'd0;
        left_4_0_clk = 1'd0;
        pe_4_1_top = 32'd0;
        pe_4_1_left = 32'd0;
        pe_4_1_go = 1'd0;
        pe_4_1_clk = 1'd0;
        top_4_1_in = 32'd0;
        top_4_1_write_en = 1'd0;
        top_4_1_clk = 1'd0;
        left_4_1_in = 32'd0;
        left_4_1_write_en = 1'd0;
        left_4_1_clk = 1'd0;
        pe_4_2_top = 32'd0;
        pe_4_2_left = 32'd0;
        pe_4_2_go = 1'd0;
        pe_4_2_clk = 1'd0;
        top_4_2_in = 32'd0;
        top_4_2_write_en = 1'd0;
        top_4_2_clk = 1'd0;
        left_4_2_in = 32'd0;
        left_4_2_write_en = 1'd0;
        left_4_2_clk = 1'd0;
        pe_4_3_top = 32'd0;
        pe_4_3_left = 32'd0;
        pe_4_3_go = 1'd0;
        pe_4_3_clk = 1'd0;
        top_4_3_in = 32'd0;
        top_4_3_write_en = 1'd0;
        top_4_3_clk = 1'd0;
        left_4_3_in = 32'd0;
        left_4_3_write_en = 1'd0;
        left_4_3_clk = 1'd0;
        pe_4_4_top = 32'd0;
        pe_4_4_left = 32'd0;
        pe_4_4_go = 1'd0;
        pe_4_4_clk = 1'd0;
        top_4_4_in = 32'd0;
        top_4_4_write_en = 1'd0;
        top_4_4_clk = 1'd0;
        left_4_4_in = 32'd0;
        left_4_4_write_en = 1'd0;
        left_4_4_clk = 1'd0;
        pe_4_5_top = 32'd0;
        pe_4_5_left = 32'd0;
        pe_4_5_go = 1'd0;
        pe_4_5_clk = 1'd0;
        top_4_5_in = 32'd0;
        top_4_5_write_en = 1'd0;
        top_4_5_clk = 1'd0;
        left_4_5_in = 32'd0;
        left_4_5_write_en = 1'd0;
        left_4_5_clk = 1'd0;
        pe_4_6_top = 32'd0;
        pe_4_6_left = 32'd0;
        pe_4_6_go = 1'd0;
        pe_4_6_clk = 1'd0;
        top_4_6_in = 32'd0;
        top_4_6_write_en = 1'd0;
        top_4_6_clk = 1'd0;
        left_4_6_in = 32'd0;
        left_4_6_write_en = 1'd0;
        left_4_6_clk = 1'd0;
        pe_4_7_top = 32'd0;
        pe_4_7_left = 32'd0;
        pe_4_7_go = 1'd0;
        pe_4_7_clk = 1'd0;
        top_4_7_in = 32'd0;
        top_4_7_write_en = 1'd0;
        top_4_7_clk = 1'd0;
        left_4_7_in = 32'd0;
        left_4_7_write_en = 1'd0;
        left_4_7_clk = 1'd0;
        pe_5_0_top = 32'd0;
        pe_5_0_left = 32'd0;
        pe_5_0_go = 1'd0;
        pe_5_0_clk = 1'd0;
        top_5_0_in = 32'd0;
        top_5_0_write_en = 1'd0;
        top_5_0_clk = 1'd0;
        left_5_0_in = 32'd0;
        left_5_0_write_en = 1'd0;
        left_5_0_clk = 1'd0;
        pe_5_1_top = 32'd0;
        pe_5_1_left = 32'd0;
        pe_5_1_go = 1'd0;
        pe_5_1_clk = 1'd0;
        top_5_1_in = 32'd0;
        top_5_1_write_en = 1'd0;
        top_5_1_clk = 1'd0;
        left_5_1_in = 32'd0;
        left_5_1_write_en = 1'd0;
        left_5_1_clk = 1'd0;
        pe_5_2_top = 32'd0;
        pe_5_2_left = 32'd0;
        pe_5_2_go = 1'd0;
        pe_5_2_clk = 1'd0;
        top_5_2_in = 32'd0;
        top_5_2_write_en = 1'd0;
        top_5_2_clk = 1'd0;
        left_5_2_in = 32'd0;
        left_5_2_write_en = 1'd0;
        left_5_2_clk = 1'd0;
        pe_5_3_top = 32'd0;
        pe_5_3_left = 32'd0;
        pe_5_3_go = 1'd0;
        pe_5_3_clk = 1'd0;
        top_5_3_in = 32'd0;
        top_5_3_write_en = 1'd0;
        top_5_3_clk = 1'd0;
        left_5_3_in = 32'd0;
        left_5_3_write_en = 1'd0;
        left_5_3_clk = 1'd0;
        pe_5_4_top = 32'd0;
        pe_5_4_left = 32'd0;
        pe_5_4_go = 1'd0;
        pe_5_4_clk = 1'd0;
        top_5_4_in = 32'd0;
        top_5_4_write_en = 1'd0;
        top_5_4_clk = 1'd0;
        left_5_4_in = 32'd0;
        left_5_4_write_en = 1'd0;
        left_5_4_clk = 1'd0;
        pe_5_5_top = 32'd0;
        pe_5_5_left = 32'd0;
        pe_5_5_go = 1'd0;
        pe_5_5_clk = 1'd0;
        top_5_5_in = 32'd0;
        top_5_5_write_en = 1'd0;
        top_5_5_clk = 1'd0;
        left_5_5_in = 32'd0;
        left_5_5_write_en = 1'd0;
        left_5_5_clk = 1'd0;
        pe_5_6_top = 32'd0;
        pe_5_6_left = 32'd0;
        pe_5_6_go = 1'd0;
        pe_5_6_clk = 1'd0;
        top_5_6_in = 32'd0;
        top_5_6_write_en = 1'd0;
        top_5_6_clk = 1'd0;
        left_5_6_in = 32'd0;
        left_5_6_write_en = 1'd0;
        left_5_6_clk = 1'd0;
        pe_5_7_top = 32'd0;
        pe_5_7_left = 32'd0;
        pe_5_7_go = 1'd0;
        pe_5_7_clk = 1'd0;
        top_5_7_in = 32'd0;
        top_5_7_write_en = 1'd0;
        top_5_7_clk = 1'd0;
        left_5_7_in = 32'd0;
        left_5_7_write_en = 1'd0;
        left_5_7_clk = 1'd0;
        pe_6_0_top = 32'd0;
        pe_6_0_left = 32'd0;
        pe_6_0_go = 1'd0;
        pe_6_0_clk = 1'd0;
        top_6_0_in = 32'd0;
        top_6_0_write_en = 1'd0;
        top_6_0_clk = 1'd0;
        left_6_0_in = 32'd0;
        left_6_0_write_en = 1'd0;
        left_6_0_clk = 1'd0;
        pe_6_1_top = 32'd0;
        pe_6_1_left = 32'd0;
        pe_6_1_go = 1'd0;
        pe_6_1_clk = 1'd0;
        top_6_1_in = 32'd0;
        top_6_1_write_en = 1'd0;
        top_6_1_clk = 1'd0;
        left_6_1_in = 32'd0;
        left_6_1_write_en = 1'd0;
        left_6_1_clk = 1'd0;
        pe_6_2_top = 32'd0;
        pe_6_2_left = 32'd0;
        pe_6_2_go = 1'd0;
        pe_6_2_clk = 1'd0;
        top_6_2_in = 32'd0;
        top_6_2_write_en = 1'd0;
        top_6_2_clk = 1'd0;
        left_6_2_in = 32'd0;
        left_6_2_write_en = 1'd0;
        left_6_2_clk = 1'd0;
        pe_6_3_top = 32'd0;
        pe_6_3_left = 32'd0;
        pe_6_3_go = 1'd0;
        pe_6_3_clk = 1'd0;
        top_6_3_in = 32'd0;
        top_6_3_write_en = 1'd0;
        top_6_3_clk = 1'd0;
        left_6_3_in = 32'd0;
        left_6_3_write_en = 1'd0;
        left_6_3_clk = 1'd0;
        pe_6_4_top = 32'd0;
        pe_6_4_left = 32'd0;
        pe_6_4_go = 1'd0;
        pe_6_4_clk = 1'd0;
        top_6_4_in = 32'd0;
        top_6_4_write_en = 1'd0;
        top_6_4_clk = 1'd0;
        left_6_4_in = 32'd0;
        left_6_4_write_en = 1'd0;
        left_6_4_clk = 1'd0;
        pe_6_5_top = 32'd0;
        pe_6_5_left = 32'd0;
        pe_6_5_go = 1'd0;
        pe_6_5_clk = 1'd0;
        top_6_5_in = 32'd0;
        top_6_5_write_en = 1'd0;
        top_6_5_clk = 1'd0;
        left_6_5_in = 32'd0;
        left_6_5_write_en = 1'd0;
        left_6_5_clk = 1'd0;
        pe_6_6_top = 32'd0;
        pe_6_6_left = 32'd0;
        pe_6_6_go = 1'd0;
        pe_6_6_clk = 1'd0;
        top_6_6_in = 32'd0;
        top_6_6_write_en = 1'd0;
        top_6_6_clk = 1'd0;
        left_6_6_in = 32'd0;
        left_6_6_write_en = 1'd0;
        left_6_6_clk = 1'd0;
        pe_6_7_top = 32'd0;
        pe_6_7_left = 32'd0;
        pe_6_7_go = 1'd0;
        pe_6_7_clk = 1'd0;
        top_6_7_in = 32'd0;
        top_6_7_write_en = 1'd0;
        top_6_7_clk = 1'd0;
        left_6_7_in = 32'd0;
        left_6_7_write_en = 1'd0;
        left_6_7_clk = 1'd0;
        pe_7_0_top = 32'd0;
        pe_7_0_left = 32'd0;
        pe_7_0_go = 1'd0;
        pe_7_0_clk = 1'd0;
        top_7_0_in = 32'd0;
        top_7_0_write_en = 1'd0;
        top_7_0_clk = 1'd0;
        left_7_0_in = 32'd0;
        left_7_0_write_en = 1'd0;
        left_7_0_clk = 1'd0;
        pe_7_1_top = 32'd0;
        pe_7_1_left = 32'd0;
        pe_7_1_go = 1'd0;
        pe_7_1_clk = 1'd0;
        top_7_1_in = 32'd0;
        top_7_1_write_en = 1'd0;
        top_7_1_clk = 1'd0;
        left_7_1_in = 32'd0;
        left_7_1_write_en = 1'd0;
        left_7_1_clk = 1'd0;
        pe_7_2_top = 32'd0;
        pe_7_2_left = 32'd0;
        pe_7_2_go = 1'd0;
        pe_7_2_clk = 1'd0;
        top_7_2_in = 32'd0;
        top_7_2_write_en = 1'd0;
        top_7_2_clk = 1'd0;
        left_7_2_in = 32'd0;
        left_7_2_write_en = 1'd0;
        left_7_2_clk = 1'd0;
        pe_7_3_top = 32'd0;
        pe_7_3_left = 32'd0;
        pe_7_3_go = 1'd0;
        pe_7_3_clk = 1'd0;
        top_7_3_in = 32'd0;
        top_7_3_write_en = 1'd0;
        top_7_3_clk = 1'd0;
        left_7_3_in = 32'd0;
        left_7_3_write_en = 1'd0;
        left_7_3_clk = 1'd0;
        pe_7_4_top = 32'd0;
        pe_7_4_left = 32'd0;
        pe_7_4_go = 1'd0;
        pe_7_4_clk = 1'd0;
        top_7_4_in = 32'd0;
        top_7_4_write_en = 1'd0;
        top_7_4_clk = 1'd0;
        left_7_4_in = 32'd0;
        left_7_4_write_en = 1'd0;
        left_7_4_clk = 1'd0;
        pe_7_5_top = 32'd0;
        pe_7_5_left = 32'd0;
        pe_7_5_go = 1'd0;
        pe_7_5_clk = 1'd0;
        top_7_5_in = 32'd0;
        top_7_5_write_en = 1'd0;
        top_7_5_clk = 1'd0;
        left_7_5_in = 32'd0;
        left_7_5_write_en = 1'd0;
        left_7_5_clk = 1'd0;
        pe_7_6_top = 32'd0;
        pe_7_6_left = 32'd0;
        pe_7_6_go = 1'd0;
        pe_7_6_clk = 1'd0;
        top_7_6_in = 32'd0;
        top_7_6_write_en = 1'd0;
        top_7_6_clk = 1'd0;
        left_7_6_in = 32'd0;
        left_7_6_write_en = 1'd0;
        left_7_6_clk = 1'd0;
        pe_7_7_top = 32'd0;
        pe_7_7_left = 32'd0;
        pe_7_7_go = 1'd0;
        pe_7_7_clk = 1'd0;
        top_7_7_in = 32'd0;
        top_7_7_write_en = 1'd0;
        top_7_7_clk = 1'd0;
        left_7_7_in = 32'd0;
        left_7_7_write_en = 1'd0;
        left_7_7_clk = 1'd0;
        fsm_in = 1'd0;
        fsm_write_en = 1'd0;
        fsm_clk = 1'd0;
        incr_left = 1'd0;
        incr_right = 1'd0;
        fsm0_in = 1'd0;
        fsm0_write_en = 1'd0;
        fsm0_clk = 1'd0;
        incr0_left = 1'd0;
        incr0_right = 1'd0;
        fsm1_in = 1'd0;
        fsm1_write_en = 1'd0;
        fsm1_clk = 1'd0;
        incr1_left = 1'd0;
        incr1_right = 1'd0;
        fsm2_in = 3'd0;
        fsm2_write_en = 1'd0;
        fsm2_clk = 1'd0;
        incr2_left = 3'd0;
        incr2_right = 3'd0;
        fsm3_in = 1'd0;
        fsm3_write_en = 1'd0;
        fsm3_clk = 1'd0;
        incr3_left = 1'd0;
        incr3_right = 1'd0;
        fsm4_in = 3'd0;
        fsm4_write_en = 1'd0;
        fsm4_clk = 1'd0;
        incr4_left = 3'd0;
        incr4_right = 3'd0;
        fsm5_in = 1'd0;
        fsm5_write_en = 1'd0;
        fsm5_clk = 1'd0;
        incr5_left = 1'd0;
        incr5_right = 1'd0;
        fsm6_in = 3'd0;
        fsm6_write_en = 1'd0;
        fsm6_clk = 1'd0;
        incr6_left = 3'd0;
        incr6_right = 3'd0;
        fsm7_in = 1'd0;
        fsm7_write_en = 1'd0;
        fsm7_clk = 1'd0;
        incr7_left = 1'd0;
        incr7_right = 1'd0;
        fsm8_in = 3'd0;
        fsm8_write_en = 1'd0;
        fsm8_clk = 1'd0;
        incr8_left = 3'd0;
        incr8_right = 3'd0;
        fsm9_in = 1'd0;
        fsm9_write_en = 1'd0;
        fsm9_clk = 1'd0;
        incr9_left = 1'd0;
        incr9_right = 1'd0;
        fsm10_in = 3'd0;
        fsm10_write_en = 1'd0;
        fsm10_clk = 1'd0;
        incr10_left = 3'd0;
        incr10_right = 3'd0;
        fsm11_in = 1'd0;
        fsm11_write_en = 1'd0;
        fsm11_clk = 1'd0;
        incr11_left = 1'd0;
        incr11_right = 1'd0;
        fsm12_in = 3'd0;
        fsm12_write_en = 1'd0;
        fsm12_clk = 1'd0;
        incr12_left = 3'd0;
        incr12_right = 3'd0;
        fsm13_in = 1'd0;
        fsm13_write_en = 1'd0;
        fsm13_clk = 1'd0;
        incr13_left = 1'd0;
        incr13_right = 1'd0;
        fsm14_in = 3'd0;
        fsm14_write_en = 1'd0;
        fsm14_clk = 1'd0;
        incr14_left = 3'd0;
        incr14_right = 3'd0;
        fsm15_in = 1'd0;
        fsm15_write_en = 1'd0;
        fsm15_clk = 1'd0;
        incr15_left = 1'd0;
        incr15_right = 1'd0;
        fsm16_in = 3'd0;
        fsm16_write_en = 1'd0;
        fsm16_clk = 1'd0;
        incr16_left = 3'd0;
        incr16_right = 3'd0;
        fsm17_in = 1'd0;
        fsm17_write_en = 1'd0;
        fsm17_clk = 1'd0;
        incr17_left = 1'd0;
        incr17_right = 1'd0;
        fsm18_in = 3'd0;
        fsm18_write_en = 1'd0;
        fsm18_clk = 1'd0;
        incr18_left = 3'd0;
        incr18_right = 3'd0;
        fsm19_in = 1'd0;
        fsm19_write_en = 1'd0;
        fsm19_clk = 1'd0;
        incr19_left = 1'd0;
        incr19_right = 1'd0;
        fsm20_in = 3'd0;
        fsm20_write_en = 1'd0;
        fsm20_clk = 1'd0;
        incr20_left = 3'd0;
        incr20_right = 3'd0;
        fsm21_in = 1'd0;
        fsm21_write_en = 1'd0;
        fsm21_clk = 1'd0;
        incr21_left = 1'd0;
        incr21_right = 1'd0;
        fsm22_in = 3'd0;
        fsm22_write_en = 1'd0;
        fsm22_clk = 1'd0;
        incr22_left = 3'd0;
        incr22_right = 3'd0;
        fsm23_in = 1'd0;
        fsm23_write_en = 1'd0;
        fsm23_clk = 1'd0;
        incr23_left = 1'd0;
        incr23_right = 1'd0;
        fsm24_in = 3'd0;
        fsm24_write_en = 1'd0;
        fsm24_clk = 1'd0;
        incr24_left = 3'd0;
        incr24_right = 3'd0;
        fsm25_in = 1'd0;
        fsm25_write_en = 1'd0;
        fsm25_clk = 1'd0;
        incr25_left = 1'd0;
        incr25_right = 1'd0;
        fsm26_in = 3'd0;
        fsm26_write_en = 1'd0;
        fsm26_clk = 1'd0;
        incr26_left = 3'd0;
        incr26_right = 3'd0;
        fsm27_in = 1'd0;
        fsm27_write_en = 1'd0;
        fsm27_clk = 1'd0;
        incr27_left = 1'd0;
        incr27_right = 1'd0;
        fsm28_in = 3'd0;
        fsm28_write_en = 1'd0;
        fsm28_clk = 1'd0;
        incr28_left = 3'd0;
        incr28_right = 3'd0;
        fsm29_in = 1'd0;
        fsm29_write_en = 1'd0;
        fsm29_clk = 1'd0;
        incr29_left = 1'd0;
        incr29_right = 1'd0;
        fsm30_in = 3'd0;
        fsm30_write_en = 1'd0;
        fsm30_clk = 1'd0;
        incr30_left = 3'd0;
        incr30_right = 3'd0;
        fsm31_in = 1'd0;
        fsm31_write_en = 1'd0;
        fsm31_clk = 1'd0;
        incr31_left = 1'd0;
        incr31_right = 1'd0;
        fsm32_in = 3'd0;
        fsm32_write_en = 1'd0;
        fsm32_clk = 1'd0;
        incr32_left = 3'd0;
        incr32_right = 3'd0;
        fsm33_in = 1'd0;
        fsm33_write_en = 1'd0;
        fsm33_clk = 1'd0;
        incr33_left = 1'd0;
        incr33_right = 1'd0;
        fsm34_in = 3'd0;
        fsm34_write_en = 1'd0;
        fsm34_clk = 1'd0;
        incr34_left = 3'd0;
        incr34_right = 3'd0;
        fsm35_in = 1'd0;
        fsm35_write_en = 1'd0;
        fsm35_clk = 1'd0;
        incr35_left = 1'd0;
        incr35_right = 1'd0;
        fsm36_in = 3'd0;
        fsm36_write_en = 1'd0;
        fsm36_clk = 1'd0;
        incr36_left = 3'd0;
        incr36_right = 3'd0;
        fsm37_in = 1'd0;
        fsm37_write_en = 1'd0;
        fsm37_clk = 1'd0;
        incr37_left = 1'd0;
        incr37_right = 1'd0;
        fsm38_in = 3'd0;
        fsm38_write_en = 1'd0;
        fsm38_clk = 1'd0;
        incr38_left = 3'd0;
        incr38_right = 3'd0;
        fsm39_in = 1'd0;
        fsm39_write_en = 1'd0;
        fsm39_clk = 1'd0;
        incr39_left = 1'd0;
        incr39_right = 1'd0;
        fsm40_in = 3'd0;
        fsm40_write_en = 1'd0;
        fsm40_clk = 1'd0;
        incr40_left = 3'd0;
        incr40_right = 3'd0;
        fsm41_in = 1'd0;
        fsm41_write_en = 1'd0;
        fsm41_clk = 1'd0;
        incr41_left = 1'd0;
        incr41_right = 1'd0;
        fsm42_in = 3'd0;
        fsm42_write_en = 1'd0;
        fsm42_clk = 1'd0;
        incr42_left = 3'd0;
        incr42_right = 3'd0;
        fsm43_in = 1'd0;
        fsm43_write_en = 1'd0;
        fsm43_clk = 1'd0;
        incr43_left = 1'd0;
        incr43_right = 1'd0;
        fsm44_in = 8'd0;
        fsm44_write_en = 1'd0;
        fsm44_clk = 1'd0;
        incr44_left = 8'd0;
        incr44_right = 8'd0;
    end
    std_reg # (
        .width(4)
    ) t0_idx (
        .clk(t0_idx_clk),
        .done(t0_idx_done),
        .in(t0_idx_in),
        .out(t0_idx_out),
        .write_en(t0_idx_write_en)
    );
    std_add # (
        .width(4)
    ) t0_add (
        .left(t0_add_left),
        .out(t0_add_out),
        .right(t0_add_right)
    );
    std_reg # (
        .width(4)
    ) t1_idx (
        .clk(t1_idx_clk),
        .done(t1_idx_done),
        .in(t1_idx_in),
        .out(t1_idx_out),
        .write_en(t1_idx_write_en)
    );
    std_add # (
        .width(4)
    ) t1_add (
        .left(t1_add_left),
        .out(t1_add_out),
        .right(t1_add_right)
    );
    std_reg # (
        .width(4)
    ) t2_idx (
        .clk(t2_idx_clk),
        .done(t2_idx_done),
        .in(t2_idx_in),
        .out(t2_idx_out),
        .write_en(t2_idx_write_en)
    );
    std_add # (
        .width(4)
    ) t2_add (
        .left(t2_add_left),
        .out(t2_add_out),
        .right(t2_add_right)
    );
    std_reg # (
        .width(4)
    ) t3_idx (
        .clk(t3_idx_clk),
        .done(t3_idx_done),
        .in(t3_idx_in),
        .out(t3_idx_out),
        .write_en(t3_idx_write_en)
    );
    std_add # (
        .width(4)
    ) t3_add (
        .left(t3_add_left),
        .out(t3_add_out),
        .right(t3_add_right)
    );
    std_reg # (
        .width(4)
    ) t4_idx (
        .clk(t4_idx_clk),
        .done(t4_idx_done),
        .in(t4_idx_in),
        .out(t4_idx_out),
        .write_en(t4_idx_write_en)
    );
    std_add # (
        .width(4)
    ) t4_add (
        .left(t4_add_left),
        .out(t4_add_out),
        .right(t4_add_right)
    );
    std_reg # (
        .width(4)
    ) t5_idx (
        .clk(t5_idx_clk),
        .done(t5_idx_done),
        .in(t5_idx_in),
        .out(t5_idx_out),
        .write_en(t5_idx_write_en)
    );
    std_add # (
        .width(4)
    ) t5_add (
        .left(t5_add_left),
        .out(t5_add_out),
        .right(t5_add_right)
    );
    std_reg # (
        .width(4)
    ) t6_idx (
        .clk(t6_idx_clk),
        .done(t6_idx_done),
        .in(t6_idx_in),
        .out(t6_idx_out),
        .write_en(t6_idx_write_en)
    );
    std_add # (
        .width(4)
    ) t6_add (
        .left(t6_add_left),
        .out(t6_add_out),
        .right(t6_add_right)
    );
    std_reg # (
        .width(4)
    ) t7_idx (
        .clk(t7_idx_clk),
        .done(t7_idx_done),
        .in(t7_idx_in),
        .out(t7_idx_out),
        .write_en(t7_idx_write_en)
    );
    std_add # (
        .width(4)
    ) t7_add (
        .left(t7_add_left),
        .out(t7_add_out),
        .right(t7_add_right)
    );
    std_reg # (
        .width(4)
    ) l0_idx (
        .clk(l0_idx_clk),
        .done(l0_idx_done),
        .in(l0_idx_in),
        .out(l0_idx_out),
        .write_en(l0_idx_write_en)
    );
    std_add # (
        .width(4)
    ) l0_add (
        .left(l0_add_left),
        .out(l0_add_out),
        .right(l0_add_right)
    );
    std_reg # (
        .width(4)
    ) l1_idx (
        .clk(l1_idx_clk),
        .done(l1_idx_done),
        .in(l1_idx_in),
        .out(l1_idx_out),
        .write_en(l1_idx_write_en)
    );
    std_add # (
        .width(4)
    ) l1_add (
        .left(l1_add_left),
        .out(l1_add_out),
        .right(l1_add_right)
    );
    std_reg # (
        .width(4)
    ) l2_idx (
        .clk(l2_idx_clk),
        .done(l2_idx_done),
        .in(l2_idx_in),
        .out(l2_idx_out),
        .write_en(l2_idx_write_en)
    );
    std_add # (
        .width(4)
    ) l2_add (
        .left(l2_add_left),
        .out(l2_add_out),
        .right(l2_add_right)
    );
    std_reg # (
        .width(4)
    ) l3_idx (
        .clk(l3_idx_clk),
        .done(l3_idx_done),
        .in(l3_idx_in),
        .out(l3_idx_out),
        .write_en(l3_idx_write_en)
    );
    std_add # (
        .width(4)
    ) l3_add (
        .left(l3_add_left),
        .out(l3_add_out),
        .right(l3_add_right)
    );
    std_reg # (
        .width(4)
    ) l4_idx (
        .clk(l4_idx_clk),
        .done(l4_idx_done),
        .in(l4_idx_in),
        .out(l4_idx_out),
        .write_en(l4_idx_write_en)
    );
    std_add # (
        .width(4)
    ) l4_add (
        .left(l4_add_left),
        .out(l4_add_out),
        .right(l4_add_right)
    );
    std_reg # (
        .width(4)
    ) l5_idx (
        .clk(l5_idx_clk),
        .done(l5_idx_done),
        .in(l5_idx_in),
        .out(l5_idx_out),
        .write_en(l5_idx_write_en)
    );
    std_add # (
        .width(4)
    ) l5_add (
        .left(l5_add_left),
        .out(l5_add_out),
        .right(l5_add_right)
    );
    std_reg # (
        .width(4)
    ) l6_idx (
        .clk(l6_idx_clk),
        .done(l6_idx_done),
        .in(l6_idx_in),
        .out(l6_idx_out),
        .write_en(l6_idx_write_en)
    );
    std_add # (
        .width(4)
    ) l6_add (
        .left(l6_add_left),
        .out(l6_add_out),
        .right(l6_add_right)
    );
    std_reg # (
        .width(4)
    ) l7_idx (
        .clk(l7_idx_clk),
        .done(l7_idx_done),
        .in(l7_idx_in),
        .out(l7_idx_out),
        .write_en(l7_idx_write_en)
    );
    std_add # (
        .width(4)
    ) l7_add (
        .left(l7_add_left),
        .out(l7_add_out),
        .right(l7_add_right)
    );
    mac_pe pe_0_0 (
        .clk(pe_0_0_clk),
        .done(pe_0_0_done),
        .go(pe_0_0_go),
        .left(pe_0_0_left),
        .out(pe_0_0_out),
        .top(pe_0_0_top)
    );
    std_reg # (
        .width(32)
    ) top_0_0 (
        .clk(top_0_0_clk),
        .done(top_0_0_done),
        .in(top_0_0_in),
        .out(top_0_0_out),
        .write_en(top_0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_0 (
        .clk(left_0_0_clk),
        .done(left_0_0_done),
        .in(left_0_0_in),
        .out(left_0_0_out),
        .write_en(left_0_0_write_en)
    );
    mac_pe pe_0_1 (
        .clk(pe_0_1_clk),
        .done(pe_0_1_done),
        .go(pe_0_1_go),
        .left(pe_0_1_left),
        .out(pe_0_1_out),
        .top(pe_0_1_top)
    );
    std_reg # (
        .width(32)
    ) top_0_1 (
        .clk(top_0_1_clk),
        .done(top_0_1_done),
        .in(top_0_1_in),
        .out(top_0_1_out),
        .write_en(top_0_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_1 (
        .clk(left_0_1_clk),
        .done(left_0_1_done),
        .in(left_0_1_in),
        .out(left_0_1_out),
        .write_en(left_0_1_write_en)
    );
    mac_pe pe_0_2 (
        .clk(pe_0_2_clk),
        .done(pe_0_2_done),
        .go(pe_0_2_go),
        .left(pe_0_2_left),
        .out(pe_0_2_out),
        .top(pe_0_2_top)
    );
    std_reg # (
        .width(32)
    ) top_0_2 (
        .clk(top_0_2_clk),
        .done(top_0_2_done),
        .in(top_0_2_in),
        .out(top_0_2_out),
        .write_en(top_0_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_2 (
        .clk(left_0_2_clk),
        .done(left_0_2_done),
        .in(left_0_2_in),
        .out(left_0_2_out),
        .write_en(left_0_2_write_en)
    );
    mac_pe pe_0_3 (
        .clk(pe_0_3_clk),
        .done(pe_0_3_done),
        .go(pe_0_3_go),
        .left(pe_0_3_left),
        .out(pe_0_3_out),
        .top(pe_0_3_top)
    );
    std_reg # (
        .width(32)
    ) top_0_3 (
        .clk(top_0_3_clk),
        .done(top_0_3_done),
        .in(top_0_3_in),
        .out(top_0_3_out),
        .write_en(top_0_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_3 (
        .clk(left_0_3_clk),
        .done(left_0_3_done),
        .in(left_0_3_in),
        .out(left_0_3_out),
        .write_en(left_0_3_write_en)
    );
    mac_pe pe_0_4 (
        .clk(pe_0_4_clk),
        .done(pe_0_4_done),
        .go(pe_0_4_go),
        .left(pe_0_4_left),
        .out(pe_0_4_out),
        .top(pe_0_4_top)
    );
    std_reg # (
        .width(32)
    ) top_0_4 (
        .clk(top_0_4_clk),
        .done(top_0_4_done),
        .in(top_0_4_in),
        .out(top_0_4_out),
        .write_en(top_0_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_4 (
        .clk(left_0_4_clk),
        .done(left_0_4_done),
        .in(left_0_4_in),
        .out(left_0_4_out),
        .write_en(left_0_4_write_en)
    );
    mac_pe pe_0_5 (
        .clk(pe_0_5_clk),
        .done(pe_0_5_done),
        .go(pe_0_5_go),
        .left(pe_0_5_left),
        .out(pe_0_5_out),
        .top(pe_0_5_top)
    );
    std_reg # (
        .width(32)
    ) top_0_5 (
        .clk(top_0_5_clk),
        .done(top_0_5_done),
        .in(top_0_5_in),
        .out(top_0_5_out),
        .write_en(top_0_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_5 (
        .clk(left_0_5_clk),
        .done(left_0_5_done),
        .in(left_0_5_in),
        .out(left_0_5_out),
        .write_en(left_0_5_write_en)
    );
    mac_pe pe_0_6 (
        .clk(pe_0_6_clk),
        .done(pe_0_6_done),
        .go(pe_0_6_go),
        .left(pe_0_6_left),
        .out(pe_0_6_out),
        .top(pe_0_6_top)
    );
    std_reg # (
        .width(32)
    ) top_0_6 (
        .clk(top_0_6_clk),
        .done(top_0_6_done),
        .in(top_0_6_in),
        .out(top_0_6_out),
        .write_en(top_0_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_6 (
        .clk(left_0_6_clk),
        .done(left_0_6_done),
        .in(left_0_6_in),
        .out(left_0_6_out),
        .write_en(left_0_6_write_en)
    );
    mac_pe pe_0_7 (
        .clk(pe_0_7_clk),
        .done(pe_0_7_done),
        .go(pe_0_7_go),
        .left(pe_0_7_left),
        .out(pe_0_7_out),
        .top(pe_0_7_top)
    );
    std_reg # (
        .width(32)
    ) top_0_7 (
        .clk(top_0_7_clk),
        .done(top_0_7_done),
        .in(top_0_7_in),
        .out(top_0_7_out),
        .write_en(top_0_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_7 (
        .clk(left_0_7_clk),
        .done(left_0_7_done),
        .in(left_0_7_in),
        .out(left_0_7_out),
        .write_en(left_0_7_write_en)
    );
    mac_pe pe_1_0 (
        .clk(pe_1_0_clk),
        .done(pe_1_0_done),
        .go(pe_1_0_go),
        .left(pe_1_0_left),
        .out(pe_1_0_out),
        .top(pe_1_0_top)
    );
    std_reg # (
        .width(32)
    ) top_1_0 (
        .clk(top_1_0_clk),
        .done(top_1_0_done),
        .in(top_1_0_in),
        .out(top_1_0_out),
        .write_en(top_1_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_0 (
        .clk(left_1_0_clk),
        .done(left_1_0_done),
        .in(left_1_0_in),
        .out(left_1_0_out),
        .write_en(left_1_0_write_en)
    );
    mac_pe pe_1_1 (
        .clk(pe_1_1_clk),
        .done(pe_1_1_done),
        .go(pe_1_1_go),
        .left(pe_1_1_left),
        .out(pe_1_1_out),
        .top(pe_1_1_top)
    );
    std_reg # (
        .width(32)
    ) top_1_1 (
        .clk(top_1_1_clk),
        .done(top_1_1_done),
        .in(top_1_1_in),
        .out(top_1_1_out),
        .write_en(top_1_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_1 (
        .clk(left_1_1_clk),
        .done(left_1_1_done),
        .in(left_1_1_in),
        .out(left_1_1_out),
        .write_en(left_1_1_write_en)
    );
    mac_pe pe_1_2 (
        .clk(pe_1_2_clk),
        .done(pe_1_2_done),
        .go(pe_1_2_go),
        .left(pe_1_2_left),
        .out(pe_1_2_out),
        .top(pe_1_2_top)
    );
    std_reg # (
        .width(32)
    ) top_1_2 (
        .clk(top_1_2_clk),
        .done(top_1_2_done),
        .in(top_1_2_in),
        .out(top_1_2_out),
        .write_en(top_1_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_2 (
        .clk(left_1_2_clk),
        .done(left_1_2_done),
        .in(left_1_2_in),
        .out(left_1_2_out),
        .write_en(left_1_2_write_en)
    );
    mac_pe pe_1_3 (
        .clk(pe_1_3_clk),
        .done(pe_1_3_done),
        .go(pe_1_3_go),
        .left(pe_1_3_left),
        .out(pe_1_3_out),
        .top(pe_1_3_top)
    );
    std_reg # (
        .width(32)
    ) top_1_3 (
        .clk(top_1_3_clk),
        .done(top_1_3_done),
        .in(top_1_3_in),
        .out(top_1_3_out),
        .write_en(top_1_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_3 (
        .clk(left_1_3_clk),
        .done(left_1_3_done),
        .in(left_1_3_in),
        .out(left_1_3_out),
        .write_en(left_1_3_write_en)
    );
    mac_pe pe_1_4 (
        .clk(pe_1_4_clk),
        .done(pe_1_4_done),
        .go(pe_1_4_go),
        .left(pe_1_4_left),
        .out(pe_1_4_out),
        .top(pe_1_4_top)
    );
    std_reg # (
        .width(32)
    ) top_1_4 (
        .clk(top_1_4_clk),
        .done(top_1_4_done),
        .in(top_1_4_in),
        .out(top_1_4_out),
        .write_en(top_1_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_4 (
        .clk(left_1_4_clk),
        .done(left_1_4_done),
        .in(left_1_4_in),
        .out(left_1_4_out),
        .write_en(left_1_4_write_en)
    );
    mac_pe pe_1_5 (
        .clk(pe_1_5_clk),
        .done(pe_1_5_done),
        .go(pe_1_5_go),
        .left(pe_1_5_left),
        .out(pe_1_5_out),
        .top(pe_1_5_top)
    );
    std_reg # (
        .width(32)
    ) top_1_5 (
        .clk(top_1_5_clk),
        .done(top_1_5_done),
        .in(top_1_5_in),
        .out(top_1_5_out),
        .write_en(top_1_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_5 (
        .clk(left_1_5_clk),
        .done(left_1_5_done),
        .in(left_1_5_in),
        .out(left_1_5_out),
        .write_en(left_1_5_write_en)
    );
    mac_pe pe_1_6 (
        .clk(pe_1_6_clk),
        .done(pe_1_6_done),
        .go(pe_1_6_go),
        .left(pe_1_6_left),
        .out(pe_1_6_out),
        .top(pe_1_6_top)
    );
    std_reg # (
        .width(32)
    ) top_1_6 (
        .clk(top_1_6_clk),
        .done(top_1_6_done),
        .in(top_1_6_in),
        .out(top_1_6_out),
        .write_en(top_1_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_6 (
        .clk(left_1_6_clk),
        .done(left_1_6_done),
        .in(left_1_6_in),
        .out(left_1_6_out),
        .write_en(left_1_6_write_en)
    );
    mac_pe pe_1_7 (
        .clk(pe_1_7_clk),
        .done(pe_1_7_done),
        .go(pe_1_7_go),
        .left(pe_1_7_left),
        .out(pe_1_7_out),
        .top(pe_1_7_top)
    );
    std_reg # (
        .width(32)
    ) top_1_7 (
        .clk(top_1_7_clk),
        .done(top_1_7_done),
        .in(top_1_7_in),
        .out(top_1_7_out),
        .write_en(top_1_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_7 (
        .clk(left_1_7_clk),
        .done(left_1_7_done),
        .in(left_1_7_in),
        .out(left_1_7_out),
        .write_en(left_1_7_write_en)
    );
    mac_pe pe_2_0 (
        .clk(pe_2_0_clk),
        .done(pe_2_0_done),
        .go(pe_2_0_go),
        .left(pe_2_0_left),
        .out(pe_2_0_out),
        .top(pe_2_0_top)
    );
    std_reg # (
        .width(32)
    ) top_2_0 (
        .clk(top_2_0_clk),
        .done(top_2_0_done),
        .in(top_2_0_in),
        .out(top_2_0_out),
        .write_en(top_2_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_0 (
        .clk(left_2_0_clk),
        .done(left_2_0_done),
        .in(left_2_0_in),
        .out(left_2_0_out),
        .write_en(left_2_0_write_en)
    );
    mac_pe pe_2_1 (
        .clk(pe_2_1_clk),
        .done(pe_2_1_done),
        .go(pe_2_1_go),
        .left(pe_2_1_left),
        .out(pe_2_1_out),
        .top(pe_2_1_top)
    );
    std_reg # (
        .width(32)
    ) top_2_1 (
        .clk(top_2_1_clk),
        .done(top_2_1_done),
        .in(top_2_1_in),
        .out(top_2_1_out),
        .write_en(top_2_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_1 (
        .clk(left_2_1_clk),
        .done(left_2_1_done),
        .in(left_2_1_in),
        .out(left_2_1_out),
        .write_en(left_2_1_write_en)
    );
    mac_pe pe_2_2 (
        .clk(pe_2_2_clk),
        .done(pe_2_2_done),
        .go(pe_2_2_go),
        .left(pe_2_2_left),
        .out(pe_2_2_out),
        .top(pe_2_2_top)
    );
    std_reg # (
        .width(32)
    ) top_2_2 (
        .clk(top_2_2_clk),
        .done(top_2_2_done),
        .in(top_2_2_in),
        .out(top_2_2_out),
        .write_en(top_2_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_2 (
        .clk(left_2_2_clk),
        .done(left_2_2_done),
        .in(left_2_2_in),
        .out(left_2_2_out),
        .write_en(left_2_2_write_en)
    );
    mac_pe pe_2_3 (
        .clk(pe_2_3_clk),
        .done(pe_2_3_done),
        .go(pe_2_3_go),
        .left(pe_2_3_left),
        .out(pe_2_3_out),
        .top(pe_2_3_top)
    );
    std_reg # (
        .width(32)
    ) top_2_3 (
        .clk(top_2_3_clk),
        .done(top_2_3_done),
        .in(top_2_3_in),
        .out(top_2_3_out),
        .write_en(top_2_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_3 (
        .clk(left_2_3_clk),
        .done(left_2_3_done),
        .in(left_2_3_in),
        .out(left_2_3_out),
        .write_en(left_2_3_write_en)
    );
    mac_pe pe_2_4 (
        .clk(pe_2_4_clk),
        .done(pe_2_4_done),
        .go(pe_2_4_go),
        .left(pe_2_4_left),
        .out(pe_2_4_out),
        .top(pe_2_4_top)
    );
    std_reg # (
        .width(32)
    ) top_2_4 (
        .clk(top_2_4_clk),
        .done(top_2_4_done),
        .in(top_2_4_in),
        .out(top_2_4_out),
        .write_en(top_2_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_4 (
        .clk(left_2_4_clk),
        .done(left_2_4_done),
        .in(left_2_4_in),
        .out(left_2_4_out),
        .write_en(left_2_4_write_en)
    );
    mac_pe pe_2_5 (
        .clk(pe_2_5_clk),
        .done(pe_2_5_done),
        .go(pe_2_5_go),
        .left(pe_2_5_left),
        .out(pe_2_5_out),
        .top(pe_2_5_top)
    );
    std_reg # (
        .width(32)
    ) top_2_5 (
        .clk(top_2_5_clk),
        .done(top_2_5_done),
        .in(top_2_5_in),
        .out(top_2_5_out),
        .write_en(top_2_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_5 (
        .clk(left_2_5_clk),
        .done(left_2_5_done),
        .in(left_2_5_in),
        .out(left_2_5_out),
        .write_en(left_2_5_write_en)
    );
    mac_pe pe_2_6 (
        .clk(pe_2_6_clk),
        .done(pe_2_6_done),
        .go(pe_2_6_go),
        .left(pe_2_6_left),
        .out(pe_2_6_out),
        .top(pe_2_6_top)
    );
    std_reg # (
        .width(32)
    ) top_2_6 (
        .clk(top_2_6_clk),
        .done(top_2_6_done),
        .in(top_2_6_in),
        .out(top_2_6_out),
        .write_en(top_2_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_6 (
        .clk(left_2_6_clk),
        .done(left_2_6_done),
        .in(left_2_6_in),
        .out(left_2_6_out),
        .write_en(left_2_6_write_en)
    );
    mac_pe pe_2_7 (
        .clk(pe_2_7_clk),
        .done(pe_2_7_done),
        .go(pe_2_7_go),
        .left(pe_2_7_left),
        .out(pe_2_7_out),
        .top(pe_2_7_top)
    );
    std_reg # (
        .width(32)
    ) top_2_7 (
        .clk(top_2_7_clk),
        .done(top_2_7_done),
        .in(top_2_7_in),
        .out(top_2_7_out),
        .write_en(top_2_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_7 (
        .clk(left_2_7_clk),
        .done(left_2_7_done),
        .in(left_2_7_in),
        .out(left_2_7_out),
        .write_en(left_2_7_write_en)
    );
    mac_pe pe_3_0 (
        .clk(pe_3_0_clk),
        .done(pe_3_0_done),
        .go(pe_3_0_go),
        .left(pe_3_0_left),
        .out(pe_3_0_out),
        .top(pe_3_0_top)
    );
    std_reg # (
        .width(32)
    ) top_3_0 (
        .clk(top_3_0_clk),
        .done(top_3_0_done),
        .in(top_3_0_in),
        .out(top_3_0_out),
        .write_en(top_3_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_0 (
        .clk(left_3_0_clk),
        .done(left_3_0_done),
        .in(left_3_0_in),
        .out(left_3_0_out),
        .write_en(left_3_0_write_en)
    );
    mac_pe pe_3_1 (
        .clk(pe_3_1_clk),
        .done(pe_3_1_done),
        .go(pe_3_1_go),
        .left(pe_3_1_left),
        .out(pe_3_1_out),
        .top(pe_3_1_top)
    );
    std_reg # (
        .width(32)
    ) top_3_1 (
        .clk(top_3_1_clk),
        .done(top_3_1_done),
        .in(top_3_1_in),
        .out(top_3_1_out),
        .write_en(top_3_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_1 (
        .clk(left_3_1_clk),
        .done(left_3_1_done),
        .in(left_3_1_in),
        .out(left_3_1_out),
        .write_en(left_3_1_write_en)
    );
    mac_pe pe_3_2 (
        .clk(pe_3_2_clk),
        .done(pe_3_2_done),
        .go(pe_3_2_go),
        .left(pe_3_2_left),
        .out(pe_3_2_out),
        .top(pe_3_2_top)
    );
    std_reg # (
        .width(32)
    ) top_3_2 (
        .clk(top_3_2_clk),
        .done(top_3_2_done),
        .in(top_3_2_in),
        .out(top_3_2_out),
        .write_en(top_3_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_2 (
        .clk(left_3_2_clk),
        .done(left_3_2_done),
        .in(left_3_2_in),
        .out(left_3_2_out),
        .write_en(left_3_2_write_en)
    );
    mac_pe pe_3_3 (
        .clk(pe_3_3_clk),
        .done(pe_3_3_done),
        .go(pe_3_3_go),
        .left(pe_3_3_left),
        .out(pe_3_3_out),
        .top(pe_3_3_top)
    );
    std_reg # (
        .width(32)
    ) top_3_3 (
        .clk(top_3_3_clk),
        .done(top_3_3_done),
        .in(top_3_3_in),
        .out(top_3_3_out),
        .write_en(top_3_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_3 (
        .clk(left_3_3_clk),
        .done(left_3_3_done),
        .in(left_3_3_in),
        .out(left_3_3_out),
        .write_en(left_3_3_write_en)
    );
    mac_pe pe_3_4 (
        .clk(pe_3_4_clk),
        .done(pe_3_4_done),
        .go(pe_3_4_go),
        .left(pe_3_4_left),
        .out(pe_3_4_out),
        .top(pe_3_4_top)
    );
    std_reg # (
        .width(32)
    ) top_3_4 (
        .clk(top_3_4_clk),
        .done(top_3_4_done),
        .in(top_3_4_in),
        .out(top_3_4_out),
        .write_en(top_3_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_4 (
        .clk(left_3_4_clk),
        .done(left_3_4_done),
        .in(left_3_4_in),
        .out(left_3_4_out),
        .write_en(left_3_4_write_en)
    );
    mac_pe pe_3_5 (
        .clk(pe_3_5_clk),
        .done(pe_3_5_done),
        .go(pe_3_5_go),
        .left(pe_3_5_left),
        .out(pe_3_5_out),
        .top(pe_3_5_top)
    );
    std_reg # (
        .width(32)
    ) top_3_5 (
        .clk(top_3_5_clk),
        .done(top_3_5_done),
        .in(top_3_5_in),
        .out(top_3_5_out),
        .write_en(top_3_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_5 (
        .clk(left_3_5_clk),
        .done(left_3_5_done),
        .in(left_3_5_in),
        .out(left_3_5_out),
        .write_en(left_3_5_write_en)
    );
    mac_pe pe_3_6 (
        .clk(pe_3_6_clk),
        .done(pe_3_6_done),
        .go(pe_3_6_go),
        .left(pe_3_6_left),
        .out(pe_3_6_out),
        .top(pe_3_6_top)
    );
    std_reg # (
        .width(32)
    ) top_3_6 (
        .clk(top_3_6_clk),
        .done(top_3_6_done),
        .in(top_3_6_in),
        .out(top_3_6_out),
        .write_en(top_3_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_6 (
        .clk(left_3_6_clk),
        .done(left_3_6_done),
        .in(left_3_6_in),
        .out(left_3_6_out),
        .write_en(left_3_6_write_en)
    );
    mac_pe pe_3_7 (
        .clk(pe_3_7_clk),
        .done(pe_3_7_done),
        .go(pe_3_7_go),
        .left(pe_3_7_left),
        .out(pe_3_7_out),
        .top(pe_3_7_top)
    );
    std_reg # (
        .width(32)
    ) top_3_7 (
        .clk(top_3_7_clk),
        .done(top_3_7_done),
        .in(top_3_7_in),
        .out(top_3_7_out),
        .write_en(top_3_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_7 (
        .clk(left_3_7_clk),
        .done(left_3_7_done),
        .in(left_3_7_in),
        .out(left_3_7_out),
        .write_en(left_3_7_write_en)
    );
    mac_pe pe_4_0 (
        .clk(pe_4_0_clk),
        .done(pe_4_0_done),
        .go(pe_4_0_go),
        .left(pe_4_0_left),
        .out(pe_4_0_out),
        .top(pe_4_0_top)
    );
    std_reg # (
        .width(32)
    ) top_4_0 (
        .clk(top_4_0_clk),
        .done(top_4_0_done),
        .in(top_4_0_in),
        .out(top_4_0_out),
        .write_en(top_4_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_0 (
        .clk(left_4_0_clk),
        .done(left_4_0_done),
        .in(left_4_0_in),
        .out(left_4_0_out),
        .write_en(left_4_0_write_en)
    );
    mac_pe pe_4_1 (
        .clk(pe_4_1_clk),
        .done(pe_4_1_done),
        .go(pe_4_1_go),
        .left(pe_4_1_left),
        .out(pe_4_1_out),
        .top(pe_4_1_top)
    );
    std_reg # (
        .width(32)
    ) top_4_1 (
        .clk(top_4_1_clk),
        .done(top_4_1_done),
        .in(top_4_1_in),
        .out(top_4_1_out),
        .write_en(top_4_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_1 (
        .clk(left_4_1_clk),
        .done(left_4_1_done),
        .in(left_4_1_in),
        .out(left_4_1_out),
        .write_en(left_4_1_write_en)
    );
    mac_pe pe_4_2 (
        .clk(pe_4_2_clk),
        .done(pe_4_2_done),
        .go(pe_4_2_go),
        .left(pe_4_2_left),
        .out(pe_4_2_out),
        .top(pe_4_2_top)
    );
    std_reg # (
        .width(32)
    ) top_4_2 (
        .clk(top_4_2_clk),
        .done(top_4_2_done),
        .in(top_4_2_in),
        .out(top_4_2_out),
        .write_en(top_4_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_2 (
        .clk(left_4_2_clk),
        .done(left_4_2_done),
        .in(left_4_2_in),
        .out(left_4_2_out),
        .write_en(left_4_2_write_en)
    );
    mac_pe pe_4_3 (
        .clk(pe_4_3_clk),
        .done(pe_4_3_done),
        .go(pe_4_3_go),
        .left(pe_4_3_left),
        .out(pe_4_3_out),
        .top(pe_4_3_top)
    );
    std_reg # (
        .width(32)
    ) top_4_3 (
        .clk(top_4_3_clk),
        .done(top_4_3_done),
        .in(top_4_3_in),
        .out(top_4_3_out),
        .write_en(top_4_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_3 (
        .clk(left_4_3_clk),
        .done(left_4_3_done),
        .in(left_4_3_in),
        .out(left_4_3_out),
        .write_en(left_4_3_write_en)
    );
    mac_pe pe_4_4 (
        .clk(pe_4_4_clk),
        .done(pe_4_4_done),
        .go(pe_4_4_go),
        .left(pe_4_4_left),
        .out(pe_4_4_out),
        .top(pe_4_4_top)
    );
    std_reg # (
        .width(32)
    ) top_4_4 (
        .clk(top_4_4_clk),
        .done(top_4_4_done),
        .in(top_4_4_in),
        .out(top_4_4_out),
        .write_en(top_4_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_4 (
        .clk(left_4_4_clk),
        .done(left_4_4_done),
        .in(left_4_4_in),
        .out(left_4_4_out),
        .write_en(left_4_4_write_en)
    );
    mac_pe pe_4_5 (
        .clk(pe_4_5_clk),
        .done(pe_4_5_done),
        .go(pe_4_5_go),
        .left(pe_4_5_left),
        .out(pe_4_5_out),
        .top(pe_4_5_top)
    );
    std_reg # (
        .width(32)
    ) top_4_5 (
        .clk(top_4_5_clk),
        .done(top_4_5_done),
        .in(top_4_5_in),
        .out(top_4_5_out),
        .write_en(top_4_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_5 (
        .clk(left_4_5_clk),
        .done(left_4_5_done),
        .in(left_4_5_in),
        .out(left_4_5_out),
        .write_en(left_4_5_write_en)
    );
    mac_pe pe_4_6 (
        .clk(pe_4_6_clk),
        .done(pe_4_6_done),
        .go(pe_4_6_go),
        .left(pe_4_6_left),
        .out(pe_4_6_out),
        .top(pe_4_6_top)
    );
    std_reg # (
        .width(32)
    ) top_4_6 (
        .clk(top_4_6_clk),
        .done(top_4_6_done),
        .in(top_4_6_in),
        .out(top_4_6_out),
        .write_en(top_4_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_6 (
        .clk(left_4_6_clk),
        .done(left_4_6_done),
        .in(left_4_6_in),
        .out(left_4_6_out),
        .write_en(left_4_6_write_en)
    );
    mac_pe pe_4_7 (
        .clk(pe_4_7_clk),
        .done(pe_4_7_done),
        .go(pe_4_7_go),
        .left(pe_4_7_left),
        .out(pe_4_7_out),
        .top(pe_4_7_top)
    );
    std_reg # (
        .width(32)
    ) top_4_7 (
        .clk(top_4_7_clk),
        .done(top_4_7_done),
        .in(top_4_7_in),
        .out(top_4_7_out),
        .write_en(top_4_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_7 (
        .clk(left_4_7_clk),
        .done(left_4_7_done),
        .in(left_4_7_in),
        .out(left_4_7_out),
        .write_en(left_4_7_write_en)
    );
    mac_pe pe_5_0 (
        .clk(pe_5_0_clk),
        .done(pe_5_0_done),
        .go(pe_5_0_go),
        .left(pe_5_0_left),
        .out(pe_5_0_out),
        .top(pe_5_0_top)
    );
    std_reg # (
        .width(32)
    ) top_5_0 (
        .clk(top_5_0_clk),
        .done(top_5_0_done),
        .in(top_5_0_in),
        .out(top_5_0_out),
        .write_en(top_5_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_0 (
        .clk(left_5_0_clk),
        .done(left_5_0_done),
        .in(left_5_0_in),
        .out(left_5_0_out),
        .write_en(left_5_0_write_en)
    );
    mac_pe pe_5_1 (
        .clk(pe_5_1_clk),
        .done(pe_5_1_done),
        .go(pe_5_1_go),
        .left(pe_5_1_left),
        .out(pe_5_1_out),
        .top(pe_5_1_top)
    );
    std_reg # (
        .width(32)
    ) top_5_1 (
        .clk(top_5_1_clk),
        .done(top_5_1_done),
        .in(top_5_1_in),
        .out(top_5_1_out),
        .write_en(top_5_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_1 (
        .clk(left_5_1_clk),
        .done(left_5_1_done),
        .in(left_5_1_in),
        .out(left_5_1_out),
        .write_en(left_5_1_write_en)
    );
    mac_pe pe_5_2 (
        .clk(pe_5_2_clk),
        .done(pe_5_2_done),
        .go(pe_5_2_go),
        .left(pe_5_2_left),
        .out(pe_5_2_out),
        .top(pe_5_2_top)
    );
    std_reg # (
        .width(32)
    ) top_5_2 (
        .clk(top_5_2_clk),
        .done(top_5_2_done),
        .in(top_5_2_in),
        .out(top_5_2_out),
        .write_en(top_5_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_2 (
        .clk(left_5_2_clk),
        .done(left_5_2_done),
        .in(left_5_2_in),
        .out(left_5_2_out),
        .write_en(left_5_2_write_en)
    );
    mac_pe pe_5_3 (
        .clk(pe_5_3_clk),
        .done(pe_5_3_done),
        .go(pe_5_3_go),
        .left(pe_5_3_left),
        .out(pe_5_3_out),
        .top(pe_5_3_top)
    );
    std_reg # (
        .width(32)
    ) top_5_3 (
        .clk(top_5_3_clk),
        .done(top_5_3_done),
        .in(top_5_3_in),
        .out(top_5_3_out),
        .write_en(top_5_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_3 (
        .clk(left_5_3_clk),
        .done(left_5_3_done),
        .in(left_5_3_in),
        .out(left_5_3_out),
        .write_en(left_5_3_write_en)
    );
    mac_pe pe_5_4 (
        .clk(pe_5_4_clk),
        .done(pe_5_4_done),
        .go(pe_5_4_go),
        .left(pe_5_4_left),
        .out(pe_5_4_out),
        .top(pe_5_4_top)
    );
    std_reg # (
        .width(32)
    ) top_5_4 (
        .clk(top_5_4_clk),
        .done(top_5_4_done),
        .in(top_5_4_in),
        .out(top_5_4_out),
        .write_en(top_5_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_4 (
        .clk(left_5_4_clk),
        .done(left_5_4_done),
        .in(left_5_4_in),
        .out(left_5_4_out),
        .write_en(left_5_4_write_en)
    );
    mac_pe pe_5_5 (
        .clk(pe_5_5_clk),
        .done(pe_5_5_done),
        .go(pe_5_5_go),
        .left(pe_5_5_left),
        .out(pe_5_5_out),
        .top(pe_5_5_top)
    );
    std_reg # (
        .width(32)
    ) top_5_5 (
        .clk(top_5_5_clk),
        .done(top_5_5_done),
        .in(top_5_5_in),
        .out(top_5_5_out),
        .write_en(top_5_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_5 (
        .clk(left_5_5_clk),
        .done(left_5_5_done),
        .in(left_5_5_in),
        .out(left_5_5_out),
        .write_en(left_5_5_write_en)
    );
    mac_pe pe_5_6 (
        .clk(pe_5_6_clk),
        .done(pe_5_6_done),
        .go(pe_5_6_go),
        .left(pe_5_6_left),
        .out(pe_5_6_out),
        .top(pe_5_6_top)
    );
    std_reg # (
        .width(32)
    ) top_5_6 (
        .clk(top_5_6_clk),
        .done(top_5_6_done),
        .in(top_5_6_in),
        .out(top_5_6_out),
        .write_en(top_5_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_6 (
        .clk(left_5_6_clk),
        .done(left_5_6_done),
        .in(left_5_6_in),
        .out(left_5_6_out),
        .write_en(left_5_6_write_en)
    );
    mac_pe pe_5_7 (
        .clk(pe_5_7_clk),
        .done(pe_5_7_done),
        .go(pe_5_7_go),
        .left(pe_5_7_left),
        .out(pe_5_7_out),
        .top(pe_5_7_top)
    );
    std_reg # (
        .width(32)
    ) top_5_7 (
        .clk(top_5_7_clk),
        .done(top_5_7_done),
        .in(top_5_7_in),
        .out(top_5_7_out),
        .write_en(top_5_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_7 (
        .clk(left_5_7_clk),
        .done(left_5_7_done),
        .in(left_5_7_in),
        .out(left_5_7_out),
        .write_en(left_5_7_write_en)
    );
    mac_pe pe_6_0 (
        .clk(pe_6_0_clk),
        .done(pe_6_0_done),
        .go(pe_6_0_go),
        .left(pe_6_0_left),
        .out(pe_6_0_out),
        .top(pe_6_0_top)
    );
    std_reg # (
        .width(32)
    ) top_6_0 (
        .clk(top_6_0_clk),
        .done(top_6_0_done),
        .in(top_6_0_in),
        .out(top_6_0_out),
        .write_en(top_6_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_0 (
        .clk(left_6_0_clk),
        .done(left_6_0_done),
        .in(left_6_0_in),
        .out(left_6_0_out),
        .write_en(left_6_0_write_en)
    );
    mac_pe pe_6_1 (
        .clk(pe_6_1_clk),
        .done(pe_6_1_done),
        .go(pe_6_1_go),
        .left(pe_6_1_left),
        .out(pe_6_1_out),
        .top(pe_6_1_top)
    );
    std_reg # (
        .width(32)
    ) top_6_1 (
        .clk(top_6_1_clk),
        .done(top_6_1_done),
        .in(top_6_1_in),
        .out(top_6_1_out),
        .write_en(top_6_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_1 (
        .clk(left_6_1_clk),
        .done(left_6_1_done),
        .in(left_6_1_in),
        .out(left_6_1_out),
        .write_en(left_6_1_write_en)
    );
    mac_pe pe_6_2 (
        .clk(pe_6_2_clk),
        .done(pe_6_2_done),
        .go(pe_6_2_go),
        .left(pe_6_2_left),
        .out(pe_6_2_out),
        .top(pe_6_2_top)
    );
    std_reg # (
        .width(32)
    ) top_6_2 (
        .clk(top_6_2_clk),
        .done(top_6_2_done),
        .in(top_6_2_in),
        .out(top_6_2_out),
        .write_en(top_6_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_2 (
        .clk(left_6_2_clk),
        .done(left_6_2_done),
        .in(left_6_2_in),
        .out(left_6_2_out),
        .write_en(left_6_2_write_en)
    );
    mac_pe pe_6_3 (
        .clk(pe_6_3_clk),
        .done(pe_6_3_done),
        .go(pe_6_3_go),
        .left(pe_6_3_left),
        .out(pe_6_3_out),
        .top(pe_6_3_top)
    );
    std_reg # (
        .width(32)
    ) top_6_3 (
        .clk(top_6_3_clk),
        .done(top_6_3_done),
        .in(top_6_3_in),
        .out(top_6_3_out),
        .write_en(top_6_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_3 (
        .clk(left_6_3_clk),
        .done(left_6_3_done),
        .in(left_6_3_in),
        .out(left_6_3_out),
        .write_en(left_6_3_write_en)
    );
    mac_pe pe_6_4 (
        .clk(pe_6_4_clk),
        .done(pe_6_4_done),
        .go(pe_6_4_go),
        .left(pe_6_4_left),
        .out(pe_6_4_out),
        .top(pe_6_4_top)
    );
    std_reg # (
        .width(32)
    ) top_6_4 (
        .clk(top_6_4_clk),
        .done(top_6_4_done),
        .in(top_6_4_in),
        .out(top_6_4_out),
        .write_en(top_6_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_4 (
        .clk(left_6_4_clk),
        .done(left_6_4_done),
        .in(left_6_4_in),
        .out(left_6_4_out),
        .write_en(left_6_4_write_en)
    );
    mac_pe pe_6_5 (
        .clk(pe_6_5_clk),
        .done(pe_6_5_done),
        .go(pe_6_5_go),
        .left(pe_6_5_left),
        .out(pe_6_5_out),
        .top(pe_6_5_top)
    );
    std_reg # (
        .width(32)
    ) top_6_5 (
        .clk(top_6_5_clk),
        .done(top_6_5_done),
        .in(top_6_5_in),
        .out(top_6_5_out),
        .write_en(top_6_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_5 (
        .clk(left_6_5_clk),
        .done(left_6_5_done),
        .in(left_6_5_in),
        .out(left_6_5_out),
        .write_en(left_6_5_write_en)
    );
    mac_pe pe_6_6 (
        .clk(pe_6_6_clk),
        .done(pe_6_6_done),
        .go(pe_6_6_go),
        .left(pe_6_6_left),
        .out(pe_6_6_out),
        .top(pe_6_6_top)
    );
    std_reg # (
        .width(32)
    ) top_6_6 (
        .clk(top_6_6_clk),
        .done(top_6_6_done),
        .in(top_6_6_in),
        .out(top_6_6_out),
        .write_en(top_6_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_6 (
        .clk(left_6_6_clk),
        .done(left_6_6_done),
        .in(left_6_6_in),
        .out(left_6_6_out),
        .write_en(left_6_6_write_en)
    );
    mac_pe pe_6_7 (
        .clk(pe_6_7_clk),
        .done(pe_6_7_done),
        .go(pe_6_7_go),
        .left(pe_6_7_left),
        .out(pe_6_7_out),
        .top(pe_6_7_top)
    );
    std_reg # (
        .width(32)
    ) top_6_7 (
        .clk(top_6_7_clk),
        .done(top_6_7_done),
        .in(top_6_7_in),
        .out(top_6_7_out),
        .write_en(top_6_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_7 (
        .clk(left_6_7_clk),
        .done(left_6_7_done),
        .in(left_6_7_in),
        .out(left_6_7_out),
        .write_en(left_6_7_write_en)
    );
    mac_pe pe_7_0 (
        .clk(pe_7_0_clk),
        .done(pe_7_0_done),
        .go(pe_7_0_go),
        .left(pe_7_0_left),
        .out(pe_7_0_out),
        .top(pe_7_0_top)
    );
    std_reg # (
        .width(32)
    ) top_7_0 (
        .clk(top_7_0_clk),
        .done(top_7_0_done),
        .in(top_7_0_in),
        .out(top_7_0_out),
        .write_en(top_7_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_0 (
        .clk(left_7_0_clk),
        .done(left_7_0_done),
        .in(left_7_0_in),
        .out(left_7_0_out),
        .write_en(left_7_0_write_en)
    );
    mac_pe pe_7_1 (
        .clk(pe_7_1_clk),
        .done(pe_7_1_done),
        .go(pe_7_1_go),
        .left(pe_7_1_left),
        .out(pe_7_1_out),
        .top(pe_7_1_top)
    );
    std_reg # (
        .width(32)
    ) top_7_1 (
        .clk(top_7_1_clk),
        .done(top_7_1_done),
        .in(top_7_1_in),
        .out(top_7_1_out),
        .write_en(top_7_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_1 (
        .clk(left_7_1_clk),
        .done(left_7_1_done),
        .in(left_7_1_in),
        .out(left_7_1_out),
        .write_en(left_7_1_write_en)
    );
    mac_pe pe_7_2 (
        .clk(pe_7_2_clk),
        .done(pe_7_2_done),
        .go(pe_7_2_go),
        .left(pe_7_2_left),
        .out(pe_7_2_out),
        .top(pe_7_2_top)
    );
    std_reg # (
        .width(32)
    ) top_7_2 (
        .clk(top_7_2_clk),
        .done(top_7_2_done),
        .in(top_7_2_in),
        .out(top_7_2_out),
        .write_en(top_7_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_2 (
        .clk(left_7_2_clk),
        .done(left_7_2_done),
        .in(left_7_2_in),
        .out(left_7_2_out),
        .write_en(left_7_2_write_en)
    );
    mac_pe pe_7_3 (
        .clk(pe_7_3_clk),
        .done(pe_7_3_done),
        .go(pe_7_3_go),
        .left(pe_7_3_left),
        .out(pe_7_3_out),
        .top(pe_7_3_top)
    );
    std_reg # (
        .width(32)
    ) top_7_3 (
        .clk(top_7_3_clk),
        .done(top_7_3_done),
        .in(top_7_3_in),
        .out(top_7_3_out),
        .write_en(top_7_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_3 (
        .clk(left_7_3_clk),
        .done(left_7_3_done),
        .in(left_7_3_in),
        .out(left_7_3_out),
        .write_en(left_7_3_write_en)
    );
    mac_pe pe_7_4 (
        .clk(pe_7_4_clk),
        .done(pe_7_4_done),
        .go(pe_7_4_go),
        .left(pe_7_4_left),
        .out(pe_7_4_out),
        .top(pe_7_4_top)
    );
    std_reg # (
        .width(32)
    ) top_7_4 (
        .clk(top_7_4_clk),
        .done(top_7_4_done),
        .in(top_7_4_in),
        .out(top_7_4_out),
        .write_en(top_7_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_4 (
        .clk(left_7_4_clk),
        .done(left_7_4_done),
        .in(left_7_4_in),
        .out(left_7_4_out),
        .write_en(left_7_4_write_en)
    );
    mac_pe pe_7_5 (
        .clk(pe_7_5_clk),
        .done(pe_7_5_done),
        .go(pe_7_5_go),
        .left(pe_7_5_left),
        .out(pe_7_5_out),
        .top(pe_7_5_top)
    );
    std_reg # (
        .width(32)
    ) top_7_5 (
        .clk(top_7_5_clk),
        .done(top_7_5_done),
        .in(top_7_5_in),
        .out(top_7_5_out),
        .write_en(top_7_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_5 (
        .clk(left_7_5_clk),
        .done(left_7_5_done),
        .in(left_7_5_in),
        .out(left_7_5_out),
        .write_en(left_7_5_write_en)
    );
    mac_pe pe_7_6 (
        .clk(pe_7_6_clk),
        .done(pe_7_6_done),
        .go(pe_7_6_go),
        .left(pe_7_6_left),
        .out(pe_7_6_out),
        .top(pe_7_6_top)
    );
    std_reg # (
        .width(32)
    ) top_7_6 (
        .clk(top_7_6_clk),
        .done(top_7_6_done),
        .in(top_7_6_in),
        .out(top_7_6_out),
        .write_en(top_7_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_6 (
        .clk(left_7_6_clk),
        .done(left_7_6_done),
        .in(left_7_6_in),
        .out(left_7_6_out),
        .write_en(left_7_6_write_en)
    );
    mac_pe pe_7_7 (
        .clk(pe_7_7_clk),
        .done(pe_7_7_done),
        .go(pe_7_7_go),
        .left(pe_7_7_left),
        .out(pe_7_7_out),
        .top(pe_7_7_top)
    );
    std_reg # (
        .width(32)
    ) top_7_7 (
        .clk(top_7_7_clk),
        .done(top_7_7_done),
        .in(top_7_7_in),
        .out(top_7_7_out),
        .write_en(top_7_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_7 (
        .clk(left_7_7_clk),
        .done(left_7_7_done),
        .in(left_7_7_in),
        .out(left_7_7_out),
        .write_en(left_7_7_write_en)
    );
    std_reg # (
        .width(1)
    ) fsm (
        .clk(fsm_clk),
        .done(fsm_done),
        .in(fsm_in),
        .out(fsm_out),
        .write_en(fsm_write_en)
    );
    std_add # (
        .width(1)
    ) incr (
        .left(incr_left),
        .out(incr_out),
        .right(incr_right)
    );
    std_reg # (
        .width(1)
    ) fsm0 (
        .clk(fsm0_clk),
        .done(fsm0_done),
        .in(fsm0_in),
        .out(fsm0_out),
        .write_en(fsm0_write_en)
    );
    std_add # (
        .width(1)
    ) incr0 (
        .left(incr0_left),
        .out(incr0_out),
        .right(incr0_right)
    );
    std_reg # (
        .width(1)
    ) fsm1 (
        .clk(fsm1_clk),
        .done(fsm1_done),
        .in(fsm1_in),
        .out(fsm1_out),
        .write_en(fsm1_write_en)
    );
    std_add # (
        .width(1)
    ) incr1 (
        .left(incr1_left),
        .out(incr1_out),
        .right(incr1_right)
    );
    std_reg # (
        .width(3)
    ) fsm2 (
        .clk(fsm2_clk),
        .done(fsm2_done),
        .in(fsm2_in),
        .out(fsm2_out),
        .write_en(fsm2_write_en)
    );
    std_add # (
        .width(3)
    ) incr2 (
        .left(incr2_left),
        .out(incr2_out),
        .right(incr2_right)
    );
    std_reg # (
        .width(1)
    ) fsm3 (
        .clk(fsm3_clk),
        .done(fsm3_done),
        .in(fsm3_in),
        .out(fsm3_out),
        .write_en(fsm3_write_en)
    );
    std_add # (
        .width(1)
    ) incr3 (
        .left(incr3_left),
        .out(incr3_out),
        .right(incr3_right)
    );
    std_reg # (
        .width(3)
    ) fsm4 (
        .clk(fsm4_clk),
        .done(fsm4_done),
        .in(fsm4_in),
        .out(fsm4_out),
        .write_en(fsm4_write_en)
    );
    std_add # (
        .width(3)
    ) incr4 (
        .left(incr4_left),
        .out(incr4_out),
        .right(incr4_right)
    );
    std_reg # (
        .width(1)
    ) fsm5 (
        .clk(fsm5_clk),
        .done(fsm5_done),
        .in(fsm5_in),
        .out(fsm5_out),
        .write_en(fsm5_write_en)
    );
    std_add # (
        .width(1)
    ) incr5 (
        .left(incr5_left),
        .out(incr5_out),
        .right(incr5_right)
    );
    std_reg # (
        .width(3)
    ) fsm6 (
        .clk(fsm6_clk),
        .done(fsm6_done),
        .in(fsm6_in),
        .out(fsm6_out),
        .write_en(fsm6_write_en)
    );
    std_add # (
        .width(3)
    ) incr6 (
        .left(incr6_left),
        .out(incr6_out),
        .right(incr6_right)
    );
    std_reg # (
        .width(1)
    ) fsm7 (
        .clk(fsm7_clk),
        .done(fsm7_done),
        .in(fsm7_in),
        .out(fsm7_out),
        .write_en(fsm7_write_en)
    );
    std_add # (
        .width(1)
    ) incr7 (
        .left(incr7_left),
        .out(incr7_out),
        .right(incr7_right)
    );
    std_reg # (
        .width(3)
    ) fsm8 (
        .clk(fsm8_clk),
        .done(fsm8_done),
        .in(fsm8_in),
        .out(fsm8_out),
        .write_en(fsm8_write_en)
    );
    std_add # (
        .width(3)
    ) incr8 (
        .left(incr8_left),
        .out(incr8_out),
        .right(incr8_right)
    );
    std_reg # (
        .width(1)
    ) fsm9 (
        .clk(fsm9_clk),
        .done(fsm9_done),
        .in(fsm9_in),
        .out(fsm9_out),
        .write_en(fsm9_write_en)
    );
    std_add # (
        .width(1)
    ) incr9 (
        .left(incr9_left),
        .out(incr9_out),
        .right(incr9_right)
    );
    std_reg # (
        .width(3)
    ) fsm10 (
        .clk(fsm10_clk),
        .done(fsm10_done),
        .in(fsm10_in),
        .out(fsm10_out),
        .write_en(fsm10_write_en)
    );
    std_add # (
        .width(3)
    ) incr10 (
        .left(incr10_left),
        .out(incr10_out),
        .right(incr10_right)
    );
    std_reg # (
        .width(1)
    ) fsm11 (
        .clk(fsm11_clk),
        .done(fsm11_done),
        .in(fsm11_in),
        .out(fsm11_out),
        .write_en(fsm11_write_en)
    );
    std_add # (
        .width(1)
    ) incr11 (
        .left(incr11_left),
        .out(incr11_out),
        .right(incr11_right)
    );
    std_reg # (
        .width(3)
    ) fsm12 (
        .clk(fsm12_clk),
        .done(fsm12_done),
        .in(fsm12_in),
        .out(fsm12_out),
        .write_en(fsm12_write_en)
    );
    std_add # (
        .width(3)
    ) incr12 (
        .left(incr12_left),
        .out(incr12_out),
        .right(incr12_right)
    );
    std_reg # (
        .width(1)
    ) fsm13 (
        .clk(fsm13_clk),
        .done(fsm13_done),
        .in(fsm13_in),
        .out(fsm13_out),
        .write_en(fsm13_write_en)
    );
    std_add # (
        .width(1)
    ) incr13 (
        .left(incr13_left),
        .out(incr13_out),
        .right(incr13_right)
    );
    std_reg # (
        .width(3)
    ) fsm14 (
        .clk(fsm14_clk),
        .done(fsm14_done),
        .in(fsm14_in),
        .out(fsm14_out),
        .write_en(fsm14_write_en)
    );
    std_add # (
        .width(3)
    ) incr14 (
        .left(incr14_left),
        .out(incr14_out),
        .right(incr14_right)
    );
    std_reg # (
        .width(1)
    ) fsm15 (
        .clk(fsm15_clk),
        .done(fsm15_done),
        .in(fsm15_in),
        .out(fsm15_out),
        .write_en(fsm15_write_en)
    );
    std_add # (
        .width(1)
    ) incr15 (
        .left(incr15_left),
        .out(incr15_out),
        .right(incr15_right)
    );
    std_reg # (
        .width(3)
    ) fsm16 (
        .clk(fsm16_clk),
        .done(fsm16_done),
        .in(fsm16_in),
        .out(fsm16_out),
        .write_en(fsm16_write_en)
    );
    std_add # (
        .width(3)
    ) incr16 (
        .left(incr16_left),
        .out(incr16_out),
        .right(incr16_right)
    );
    std_reg # (
        .width(1)
    ) fsm17 (
        .clk(fsm17_clk),
        .done(fsm17_done),
        .in(fsm17_in),
        .out(fsm17_out),
        .write_en(fsm17_write_en)
    );
    std_add # (
        .width(1)
    ) incr17 (
        .left(incr17_left),
        .out(incr17_out),
        .right(incr17_right)
    );
    std_reg # (
        .width(3)
    ) fsm18 (
        .clk(fsm18_clk),
        .done(fsm18_done),
        .in(fsm18_in),
        .out(fsm18_out),
        .write_en(fsm18_write_en)
    );
    std_add # (
        .width(3)
    ) incr18 (
        .left(incr18_left),
        .out(incr18_out),
        .right(incr18_right)
    );
    std_reg # (
        .width(1)
    ) fsm19 (
        .clk(fsm19_clk),
        .done(fsm19_done),
        .in(fsm19_in),
        .out(fsm19_out),
        .write_en(fsm19_write_en)
    );
    std_add # (
        .width(1)
    ) incr19 (
        .left(incr19_left),
        .out(incr19_out),
        .right(incr19_right)
    );
    std_reg # (
        .width(3)
    ) fsm20 (
        .clk(fsm20_clk),
        .done(fsm20_done),
        .in(fsm20_in),
        .out(fsm20_out),
        .write_en(fsm20_write_en)
    );
    std_add # (
        .width(3)
    ) incr20 (
        .left(incr20_left),
        .out(incr20_out),
        .right(incr20_right)
    );
    std_reg # (
        .width(1)
    ) fsm21 (
        .clk(fsm21_clk),
        .done(fsm21_done),
        .in(fsm21_in),
        .out(fsm21_out),
        .write_en(fsm21_write_en)
    );
    std_add # (
        .width(1)
    ) incr21 (
        .left(incr21_left),
        .out(incr21_out),
        .right(incr21_right)
    );
    std_reg # (
        .width(3)
    ) fsm22 (
        .clk(fsm22_clk),
        .done(fsm22_done),
        .in(fsm22_in),
        .out(fsm22_out),
        .write_en(fsm22_write_en)
    );
    std_add # (
        .width(3)
    ) incr22 (
        .left(incr22_left),
        .out(incr22_out),
        .right(incr22_right)
    );
    std_reg # (
        .width(1)
    ) fsm23 (
        .clk(fsm23_clk),
        .done(fsm23_done),
        .in(fsm23_in),
        .out(fsm23_out),
        .write_en(fsm23_write_en)
    );
    std_add # (
        .width(1)
    ) incr23 (
        .left(incr23_left),
        .out(incr23_out),
        .right(incr23_right)
    );
    std_reg # (
        .width(3)
    ) fsm24 (
        .clk(fsm24_clk),
        .done(fsm24_done),
        .in(fsm24_in),
        .out(fsm24_out),
        .write_en(fsm24_write_en)
    );
    std_add # (
        .width(3)
    ) incr24 (
        .left(incr24_left),
        .out(incr24_out),
        .right(incr24_right)
    );
    std_reg # (
        .width(1)
    ) fsm25 (
        .clk(fsm25_clk),
        .done(fsm25_done),
        .in(fsm25_in),
        .out(fsm25_out),
        .write_en(fsm25_write_en)
    );
    std_add # (
        .width(1)
    ) incr25 (
        .left(incr25_left),
        .out(incr25_out),
        .right(incr25_right)
    );
    std_reg # (
        .width(3)
    ) fsm26 (
        .clk(fsm26_clk),
        .done(fsm26_done),
        .in(fsm26_in),
        .out(fsm26_out),
        .write_en(fsm26_write_en)
    );
    std_add # (
        .width(3)
    ) incr26 (
        .left(incr26_left),
        .out(incr26_out),
        .right(incr26_right)
    );
    std_reg # (
        .width(1)
    ) fsm27 (
        .clk(fsm27_clk),
        .done(fsm27_done),
        .in(fsm27_in),
        .out(fsm27_out),
        .write_en(fsm27_write_en)
    );
    std_add # (
        .width(1)
    ) incr27 (
        .left(incr27_left),
        .out(incr27_out),
        .right(incr27_right)
    );
    std_reg # (
        .width(3)
    ) fsm28 (
        .clk(fsm28_clk),
        .done(fsm28_done),
        .in(fsm28_in),
        .out(fsm28_out),
        .write_en(fsm28_write_en)
    );
    std_add # (
        .width(3)
    ) incr28 (
        .left(incr28_left),
        .out(incr28_out),
        .right(incr28_right)
    );
    std_reg # (
        .width(1)
    ) fsm29 (
        .clk(fsm29_clk),
        .done(fsm29_done),
        .in(fsm29_in),
        .out(fsm29_out),
        .write_en(fsm29_write_en)
    );
    std_add # (
        .width(1)
    ) incr29 (
        .left(incr29_left),
        .out(incr29_out),
        .right(incr29_right)
    );
    std_reg # (
        .width(3)
    ) fsm30 (
        .clk(fsm30_clk),
        .done(fsm30_done),
        .in(fsm30_in),
        .out(fsm30_out),
        .write_en(fsm30_write_en)
    );
    std_add # (
        .width(3)
    ) incr30 (
        .left(incr30_left),
        .out(incr30_out),
        .right(incr30_right)
    );
    std_reg # (
        .width(1)
    ) fsm31 (
        .clk(fsm31_clk),
        .done(fsm31_done),
        .in(fsm31_in),
        .out(fsm31_out),
        .write_en(fsm31_write_en)
    );
    std_add # (
        .width(1)
    ) incr31 (
        .left(incr31_left),
        .out(incr31_out),
        .right(incr31_right)
    );
    std_reg # (
        .width(3)
    ) fsm32 (
        .clk(fsm32_clk),
        .done(fsm32_done),
        .in(fsm32_in),
        .out(fsm32_out),
        .write_en(fsm32_write_en)
    );
    std_add # (
        .width(3)
    ) incr32 (
        .left(incr32_left),
        .out(incr32_out),
        .right(incr32_right)
    );
    std_reg # (
        .width(1)
    ) fsm33 (
        .clk(fsm33_clk),
        .done(fsm33_done),
        .in(fsm33_in),
        .out(fsm33_out),
        .write_en(fsm33_write_en)
    );
    std_add # (
        .width(1)
    ) incr33 (
        .left(incr33_left),
        .out(incr33_out),
        .right(incr33_right)
    );
    std_reg # (
        .width(3)
    ) fsm34 (
        .clk(fsm34_clk),
        .done(fsm34_done),
        .in(fsm34_in),
        .out(fsm34_out),
        .write_en(fsm34_write_en)
    );
    std_add # (
        .width(3)
    ) incr34 (
        .left(incr34_left),
        .out(incr34_out),
        .right(incr34_right)
    );
    std_reg # (
        .width(1)
    ) fsm35 (
        .clk(fsm35_clk),
        .done(fsm35_done),
        .in(fsm35_in),
        .out(fsm35_out),
        .write_en(fsm35_write_en)
    );
    std_add # (
        .width(1)
    ) incr35 (
        .left(incr35_left),
        .out(incr35_out),
        .right(incr35_right)
    );
    std_reg # (
        .width(3)
    ) fsm36 (
        .clk(fsm36_clk),
        .done(fsm36_done),
        .in(fsm36_in),
        .out(fsm36_out),
        .write_en(fsm36_write_en)
    );
    std_add # (
        .width(3)
    ) incr36 (
        .left(incr36_left),
        .out(incr36_out),
        .right(incr36_right)
    );
    std_reg # (
        .width(1)
    ) fsm37 (
        .clk(fsm37_clk),
        .done(fsm37_done),
        .in(fsm37_in),
        .out(fsm37_out),
        .write_en(fsm37_write_en)
    );
    std_add # (
        .width(1)
    ) incr37 (
        .left(incr37_left),
        .out(incr37_out),
        .right(incr37_right)
    );
    std_reg # (
        .width(3)
    ) fsm38 (
        .clk(fsm38_clk),
        .done(fsm38_done),
        .in(fsm38_in),
        .out(fsm38_out),
        .write_en(fsm38_write_en)
    );
    std_add # (
        .width(3)
    ) incr38 (
        .left(incr38_left),
        .out(incr38_out),
        .right(incr38_right)
    );
    std_reg # (
        .width(1)
    ) fsm39 (
        .clk(fsm39_clk),
        .done(fsm39_done),
        .in(fsm39_in),
        .out(fsm39_out),
        .write_en(fsm39_write_en)
    );
    std_add # (
        .width(1)
    ) incr39 (
        .left(incr39_left),
        .out(incr39_out),
        .right(incr39_right)
    );
    std_reg # (
        .width(3)
    ) fsm40 (
        .clk(fsm40_clk),
        .done(fsm40_done),
        .in(fsm40_in),
        .out(fsm40_out),
        .write_en(fsm40_write_en)
    );
    std_add # (
        .width(3)
    ) incr40 (
        .left(incr40_left),
        .out(incr40_out),
        .right(incr40_right)
    );
    std_reg # (
        .width(1)
    ) fsm41 (
        .clk(fsm41_clk),
        .done(fsm41_done),
        .in(fsm41_in),
        .out(fsm41_out),
        .write_en(fsm41_write_en)
    );
    std_add # (
        .width(1)
    ) incr41 (
        .left(incr41_left),
        .out(incr41_out),
        .right(incr41_right)
    );
    std_reg # (
        .width(3)
    ) fsm42 (
        .clk(fsm42_clk),
        .done(fsm42_done),
        .in(fsm42_in),
        .out(fsm42_out),
        .write_en(fsm42_write_en)
    );
    std_add # (
        .width(3)
    ) incr42 (
        .left(incr42_left),
        .out(incr42_out),
        .right(incr42_right)
    );
    std_reg # (
        .width(1)
    ) fsm43 (
        .clk(fsm43_clk),
        .done(fsm43_done),
        .in(fsm43_in),
        .out(fsm43_out),
        .write_en(fsm43_write_en)
    );
    std_add # (
        .width(1)
    ) incr43 (
        .left(incr43_left),
        .out(incr43_out),
        .right(incr43_right)
    );
    std_reg # (
        .width(8)
    ) fsm44 (
        .clk(fsm44_clk),
        .done(fsm44_done),
        .in(fsm44_in),
        .out(fsm44_out),
        .write_en(fsm44_write_en)
    );
    std_add # (
        .width(8)
    ) incr44 (
        .left(incr44_left),
        .out(incr44_out),
        .right(incr44_right)
    );
    assign done =
     fsm44_out == 8'd134 ? 1'd1 : 1'd0;
    assign l0_addr0 =
     fsm1_out < 1'd1 & fsm44_out == 8'd2 & go | fsm3_out < 1'd1 & fsm44_out == 8'd8 & go | fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go ? l0_idx_out : 4'd0;
    assign l0_clk =
     1'b1 ? clk : 1'd0;
    assign l1_addr0 =
     fsm3_out < 1'd1 & fsm44_out == 8'd8 & go | fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go ? l1_idx_out : 4'd0;
    assign l1_clk =
     1'b1 ? clk : 1'd0;
    assign l2_addr0 =
     fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go ? l2_idx_out : 4'd0;
    assign l2_clk =
     1'b1 ? clk : 1'd0;
    assign l3_addr0 =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? l3_idx_out : 4'd0;
    assign l3_clk =
     1'b1 ? clk : 1'd0;
    assign l4_addr0 =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? l4_idx_out : 4'd0;
    assign l4_clk =
     1'b1 ? clk : 1'd0;
    assign l5_addr0 =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? l5_idx_out : 4'd0;
    assign l5_clk =
     1'b1 ? clk : 1'd0;
    assign l6_addr0 =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? l6_idx_out : 4'd0;
    assign l6_clk =
     1'b1 ? clk : 1'd0;
    assign l7_addr0 =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? l7_idx_out : 4'd0;
    assign l7_clk =
     1'b1 ? clk : 1'd0;
    assign t0_addr0 =
     fsm1_out < 1'd1 & fsm44_out == 8'd2 & go | fsm3_out < 1'd1 & fsm44_out == 8'd8 & go | fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go ? t0_idx_out : 4'd0;
    assign t0_clk =
     1'b1 ? clk : 1'd0;
    assign t1_addr0 =
     fsm3_out < 1'd1 & fsm44_out == 8'd8 & go | fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go ? t1_idx_out : 4'd0;
    assign t1_clk =
     1'b1 ? clk : 1'd0;
    assign t2_addr0 =
     fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go ? t2_idx_out : 4'd0;
    assign t2_clk =
     1'b1 ? clk : 1'd0;
    assign t3_addr0 =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? t3_idx_out : 4'd0;
    assign t3_clk =
     1'b1 ? clk : 1'd0;
    assign t4_addr0 =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? t4_idx_out : 4'd0;
    assign t4_clk =
     1'b1 ? clk : 1'd0;
    assign t5_addr0 =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? t5_idx_out : 4'd0;
    assign t5_clk =
     1'b1 ? clk : 1'd0;
    assign t6_addr0 =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? t6_idx_out : 4'd0;
    assign t6_clk =
     1'b1 ? clk : 1'd0;
    assign t7_addr0 =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? t7_idx_out : 4'd0;
    assign t7_clk =
     1'b1 ? clk : 1'd0;
    assign fsm_clk =
     1'b1 ? clk : 1'd0;
    assign fsm_in =
     fsm_out == 1'd1 ? 1'd0 :
     fsm_out != 1'd1 & fsm44_out == 8'd0 & go ? incr_out : 1'd0;
    assign fsm_write_en =
     fsm_out != 1'd1 & fsm44_out == 8'd0 & go | fsm_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm0_clk =
     1'b1 ? clk : 1'd0;
    assign fsm0_in =
     fsm0_out == 1'd1 ? 1'd0 :
     fsm0_out != 1'd1 & fsm44_out == 8'd1 & go ? incr0_out : 1'd0;
    assign fsm0_write_en =
     fsm0_out != 1'd1 & fsm44_out == 8'd1 & go | fsm0_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm1_clk =
     1'b1 ? clk : 1'd0;
    assign fsm1_in =
     fsm1_out == 1'd1 ? 1'd0 :
     fsm1_out != 1'd1 & fsm44_out == 8'd2 & go ? incr1_out : 1'd0;
    assign fsm1_write_en =
     fsm1_out != 1'd1 & fsm44_out == 8'd2 & go | fsm1_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm10_clk =
     1'b1 ? clk : 1'd0;
    assign fsm10_in =
     fsm10_out == 3'd5 ? 3'd0 :
     fsm10_out != 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go ? incr10_out : 3'd0;
    assign fsm10_write_en =
     fsm10_out != 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm10_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm11_clk =
     1'b1 ? clk : 1'd0;
    assign fsm11_in =
     fsm11_out == 1'd1 ? 1'd0 :
     fsm11_out != 1'd1 & fsm44_out == 8'd32 & go ? incr11_out : 1'd0;
    assign fsm11_write_en =
     fsm11_out != 1'd1 & fsm44_out == 8'd32 & go | fsm11_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm12_clk =
     1'b1 ? clk : 1'd0;
    assign fsm12_in =
     fsm12_out == 3'd5 ? 3'd0 :
     fsm12_out != 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go ? incr12_out : 3'd0;
    assign fsm12_write_en =
     fsm12_out != 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm12_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm13_clk =
     1'b1 ? clk : 1'd0;
    assign fsm13_in =
     fsm13_out == 1'd1 ? 1'd0 :
     fsm13_out != 1'd1 & fsm44_out == 8'd38 & go ? incr13_out : 1'd0;
    assign fsm13_write_en =
     fsm13_out != 1'd1 & fsm44_out == 8'd38 & go | fsm13_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm14_clk =
     1'b1 ? clk : 1'd0;
    assign fsm14_in =
     fsm14_out == 3'd5 ? 3'd0 :
     fsm14_out != 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go ? incr14_out : 3'd0;
    assign fsm14_write_en =
     fsm14_out != 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm14_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm15_clk =
     1'b1 ? clk : 1'd0;
    assign fsm15_in =
     fsm15_out == 1'd1 ? 1'd0 :
     fsm15_out != 1'd1 & fsm44_out == 8'd44 & go ? incr15_out : 1'd0;
    assign fsm15_write_en =
     fsm15_out != 1'd1 & fsm44_out == 8'd44 & go | fsm15_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm16_clk =
     1'b1 ? clk : 1'd0;
    assign fsm16_in =
     fsm16_out == 3'd5 ? 3'd0 :
     fsm16_out != 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go ? incr16_out : 3'd0;
    assign fsm16_write_en =
     fsm16_out != 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm16_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm17_clk =
     1'b1 ? clk : 1'd0;
    assign fsm17_in =
     fsm17_out == 1'd1 ? 1'd0 :
     fsm17_out != 1'd1 & fsm44_out == 8'd50 & go ? incr17_out : 1'd0;
    assign fsm17_write_en =
     fsm17_out != 1'd1 & fsm44_out == 8'd50 & go | fsm17_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm18_clk =
     1'b1 ? clk : 1'd0;
    assign fsm18_in =
     fsm18_out == 3'd5 ? 3'd0 :
     fsm18_out != 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? incr18_out : 3'd0;
    assign fsm18_write_en =
     fsm18_out != 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm18_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm19_clk =
     1'b1 ? clk : 1'd0;
    assign fsm19_in =
     fsm19_out == 1'd1 ? 1'd0 :
     fsm19_out != 1'd1 & fsm44_out == 8'd56 & go ? incr19_out : 1'd0;
    assign fsm19_write_en =
     fsm19_out != 1'd1 & fsm44_out == 8'd56 & go | fsm19_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm2_clk =
     1'b1 ? clk : 1'd0;
    assign fsm2_in =
     fsm2_out == 3'd5 ? 3'd0 :
     fsm2_out != 3'd5 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go ? incr2_out : 3'd0;
    assign fsm2_write_en =
     fsm2_out != 3'd5 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm2_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm20_clk =
     1'b1 ? clk : 1'd0;
    assign fsm20_in =
     fsm20_out == 3'd5 ? 3'd0 :
     fsm20_out != 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? incr20_out : 3'd0;
    assign fsm20_write_en =
     fsm20_out != 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm20_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm21_clk =
     1'b1 ? clk : 1'd0;
    assign fsm21_in =
     fsm21_out == 1'd1 ? 1'd0 :
     fsm21_out != 1'd1 & fsm44_out == 8'd62 & go ? incr21_out : 1'd0;
    assign fsm21_write_en =
     fsm21_out != 1'd1 & fsm44_out == 8'd62 & go | fsm21_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm22_clk =
     1'b1 ? clk : 1'd0;
    assign fsm22_in =
     fsm22_out == 3'd5 ? 3'd0 :
     fsm22_out != 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? incr22_out : 3'd0;
    assign fsm22_write_en =
     fsm22_out != 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm22_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm23_clk =
     1'b1 ? clk : 1'd0;
    assign fsm23_in =
     fsm23_out == 1'd1 ? 1'd0 :
     fsm23_out != 1'd1 & fsm44_out == 8'd68 & go ? incr23_out : 1'd0;
    assign fsm23_write_en =
     fsm23_out != 1'd1 & fsm44_out == 8'd68 & go | fsm23_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm24_clk =
     1'b1 ? clk : 1'd0;
    assign fsm24_in =
     fsm24_out == 3'd5 ? 3'd0 :
     fsm24_out != 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? incr24_out : 3'd0;
    assign fsm24_write_en =
     fsm24_out != 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm24_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm25_clk =
     1'b1 ? clk : 1'd0;
    assign fsm25_in =
     fsm25_out == 1'd1 ? 1'd0 :
     fsm25_out != 1'd1 & fsm44_out == 8'd74 & go ? incr25_out : 1'd0;
    assign fsm25_write_en =
     fsm25_out != 1'd1 & fsm44_out == 8'd74 & go | fsm25_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm26_clk =
     1'b1 ? clk : 1'd0;
    assign fsm26_in =
     fsm26_out == 3'd5 ? 3'd0 :
     fsm26_out != 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? incr26_out : 3'd0;
    assign fsm26_write_en =
     fsm26_out != 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm26_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm27_clk =
     1'b1 ? clk : 1'd0;
    assign fsm27_in =
     fsm27_out == 1'd1 ? 1'd0 :
     fsm27_out != 1'd1 & fsm44_out == 8'd80 & go ? incr27_out : 1'd0;
    assign fsm27_write_en =
     fsm27_out != 1'd1 & fsm44_out == 8'd80 & go | fsm27_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm28_clk =
     1'b1 ? clk : 1'd0;
    assign fsm28_in =
     fsm28_out == 3'd5 ? 3'd0 :
     fsm28_out != 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? incr28_out : 3'd0;
    assign fsm28_write_en =
     fsm28_out != 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm28_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm29_clk =
     1'b1 ? clk : 1'd0;
    assign fsm29_in =
     fsm29_out == 1'd1 ? 1'd0 :
     fsm29_out != 1'd1 & fsm44_out == 8'd86 & go ? incr29_out : 1'd0;
    assign fsm29_write_en =
     fsm29_out != 1'd1 & fsm44_out == 8'd86 & go | fsm29_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm3_clk =
     1'b1 ? clk : 1'd0;
    assign fsm3_in =
     fsm3_out == 1'd1 ? 1'd0 :
     fsm3_out != 1'd1 & fsm44_out == 8'd8 & go ? incr3_out : 1'd0;
    assign fsm3_write_en =
     fsm3_out != 1'd1 & fsm44_out == 8'd8 & go | fsm3_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm30_clk =
     1'b1 ? clk : 1'd0;
    assign fsm30_in =
     fsm30_out == 3'd5 ? 3'd0 :
     fsm30_out != 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? incr30_out : 3'd0;
    assign fsm30_write_en =
     fsm30_out != 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm30_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm31_clk =
     1'b1 ? clk : 1'd0;
    assign fsm31_in =
     fsm31_out == 1'd1 ? 1'd0 :
     fsm31_out != 1'd1 & fsm44_out == 8'd92 & go ? incr31_out : 1'd0;
    assign fsm31_write_en =
     fsm31_out != 1'd1 & fsm44_out == 8'd92 & go | fsm31_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm32_clk =
     1'b1 ? clk : 1'd0;
    assign fsm32_in =
     fsm32_out == 3'd5 ? 3'd0 :
     fsm32_out != 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? incr32_out : 3'd0;
    assign fsm32_write_en =
     fsm32_out != 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm32_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm33_clk =
     1'b1 ? clk : 1'd0;
    assign fsm33_in =
     fsm33_out == 1'd1 ? 1'd0 :
     fsm33_out != 1'd1 & fsm44_out == 8'd98 & go ? incr33_out : 1'd0;
    assign fsm33_write_en =
     fsm33_out != 1'd1 & fsm44_out == 8'd98 & go | fsm33_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm34_clk =
     1'b1 ? clk : 1'd0;
    assign fsm34_in =
     fsm34_out == 3'd5 ? 3'd0 :
     fsm34_out != 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? incr34_out : 3'd0;
    assign fsm34_write_en =
     fsm34_out != 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm34_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm35_clk =
     1'b1 ? clk : 1'd0;
    assign fsm35_in =
     fsm35_out == 1'd1 ? 1'd0 :
     fsm35_out != 1'd1 & fsm44_out == 8'd104 & go ? incr35_out : 1'd0;
    assign fsm35_write_en =
     fsm35_out != 1'd1 & fsm44_out == 8'd104 & go | fsm35_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm36_clk =
     1'b1 ? clk : 1'd0;
    assign fsm36_in =
     fsm36_out == 3'd5 ? 3'd0 :
     fsm36_out != 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? incr36_out : 3'd0;
    assign fsm36_write_en =
     fsm36_out != 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm36_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm37_clk =
     1'b1 ? clk : 1'd0;
    assign fsm37_in =
     fsm37_out == 1'd1 ? 1'd0 :
     fsm37_out != 1'd1 & fsm44_out == 8'd110 & go ? incr37_out : 1'd0;
    assign fsm37_write_en =
     fsm37_out != 1'd1 & fsm44_out == 8'd110 & go | fsm37_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm38_clk =
     1'b1 ? clk : 1'd0;
    assign fsm38_in =
     fsm38_out == 3'd5 ? 3'd0 :
     fsm38_out != 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go ? incr38_out : 3'd0;
    assign fsm38_write_en =
     fsm38_out != 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm38_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm39_clk =
     1'b1 ? clk : 1'd0;
    assign fsm39_in =
     fsm39_out == 1'd1 ? 1'd0 :
     fsm39_out != 1'd1 & fsm44_out == 8'd116 & go ? incr39_out : 1'd0;
    assign fsm39_write_en =
     fsm39_out != 1'd1 & fsm44_out == 8'd116 & go | fsm39_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm4_clk =
     1'b1 ? clk : 1'd0;
    assign fsm4_in =
     fsm4_out == 3'd5 ? 3'd0 :
     fsm4_out != 3'd5 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go ? incr4_out : 3'd0;
    assign fsm4_write_en =
     fsm4_out != 3'd5 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm4_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm40_clk =
     1'b1 ? clk : 1'd0;
    assign fsm40_in =
     fsm40_out == 3'd5 ? 3'd0 :
     fsm40_out != 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go ? incr40_out : 3'd0;
    assign fsm40_write_en =
     fsm40_out != 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go | fsm40_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm41_clk =
     1'b1 ? clk : 1'd0;
    assign fsm41_in =
     fsm41_out == 1'd1 ? 1'd0 :
     fsm41_out != 1'd1 & fsm44_out == 8'd122 & go ? incr41_out : 1'd0;
    assign fsm41_write_en =
     fsm41_out != 1'd1 & fsm44_out == 8'd122 & go | fsm41_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm42_clk =
     1'b1 ? clk : 1'd0;
    assign fsm42_in =
     fsm42_out == 3'd5 ? 3'd0 :
     fsm42_out != 3'd5 & fsm44_out >= 8'd123 & fsm44_out < 8'd128 & go ? incr42_out : 3'd0;
    assign fsm42_write_en =
     fsm42_out != 3'd5 & fsm44_out >= 8'd123 & fsm44_out < 8'd128 & go | fsm42_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm43_clk =
     1'b1 ? clk : 1'd0;
    assign fsm43_in =
     fsm43_out == 1'd1 ? 1'd0 :
     fsm43_out != 1'd1 & fsm44_out == 8'd128 & go ? incr43_out : 1'd0;
    assign fsm43_write_en =
     fsm43_out != 1'd1 & fsm44_out == 8'd128 & go | fsm43_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm44_clk =
     1'b1 ? clk : 1'd0;
    assign fsm44_in =
     fsm44_out == 8'd134 ? 8'd0 :
     fsm44_out != 8'd134 & go ? incr44_out : 8'd0;
    assign fsm44_write_en =
     fsm44_out != 8'd134 & go | fsm44_out == 8'd134 ? 1'd1 : 1'd0;
    assign fsm5_clk =
     1'b1 ? clk : 1'd0;
    assign fsm5_in =
     fsm5_out == 1'd1 ? 1'd0 :
     fsm5_out != 1'd1 & fsm44_out == 8'd14 & go ? incr5_out : 1'd0;
    assign fsm5_write_en =
     fsm5_out != 1'd1 & fsm44_out == 8'd14 & go | fsm5_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm6_clk =
     1'b1 ? clk : 1'd0;
    assign fsm6_in =
     fsm6_out == 3'd5 ? 3'd0 :
     fsm6_out != 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go ? incr6_out : 3'd0;
    assign fsm6_write_en =
     fsm6_out != 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm6_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm7_clk =
     1'b1 ? clk : 1'd0;
    assign fsm7_in =
     fsm7_out == 1'd1 ? 1'd0 :
     fsm7_out != 1'd1 & fsm44_out == 8'd20 & go ? incr7_out : 1'd0;
    assign fsm7_write_en =
     fsm7_out != 1'd1 & fsm44_out == 8'd20 & go | fsm7_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm8_clk =
     1'b1 ? clk : 1'd0;
    assign fsm8_in =
     fsm8_out == 3'd5 ? 3'd0 :
     fsm8_out != 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go ? incr8_out : 3'd0;
    assign fsm8_write_en =
     fsm8_out != 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm8_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm9_clk =
     1'b1 ? clk : 1'd0;
    assign fsm9_in =
     fsm9_out == 1'd1 ? 1'd0 :
     fsm9_out != 1'd1 & fsm44_out == 8'd26 & go ? incr9_out : 1'd0;
    assign fsm9_write_en =
     fsm9_out != 1'd1 & fsm44_out == 8'd26 & go | fsm9_out == 1'd1 ? 1'd1 : 1'd0;
    assign incr_left =
     fsm44_out == 8'd0 & go ? 1'd1 : 1'd0;
    assign incr_right =
     fsm44_out == 8'd0 & go ? fsm_out : 1'd0;
    assign incr0_left =
     fsm44_out == 8'd1 & go ? 1'd1 : 1'd0;
    assign incr0_right =
     fsm44_out == 8'd1 & go ? fsm0_out : 1'd0;
    assign incr1_left =
     fsm44_out == 8'd2 & go ? 1'd1 : 1'd0;
    assign incr1_right =
     fsm44_out == 8'd2 & go ? fsm1_out : 1'd0;
    assign incr10_left =
     fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go ? 3'd1 : 3'd0;
    assign incr10_right =
     fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go ? fsm10_out : 3'd0;
    assign incr11_left =
     fsm44_out == 8'd32 & go ? 1'd1 : 1'd0;
    assign incr11_right =
     fsm44_out == 8'd32 & go ? fsm11_out : 1'd0;
    assign incr12_left =
     fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go ? 3'd1 : 3'd0;
    assign incr12_right =
     fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go ? fsm12_out : 3'd0;
    assign incr13_left =
     fsm44_out == 8'd38 & go ? 1'd1 : 1'd0;
    assign incr13_right =
     fsm44_out == 8'd38 & go ? fsm13_out : 1'd0;
    assign incr14_left =
     fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go ? 3'd1 : 3'd0;
    assign incr14_right =
     fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go ? fsm14_out : 3'd0;
    assign incr15_left =
     fsm44_out == 8'd44 & go ? 1'd1 : 1'd0;
    assign incr15_right =
     fsm44_out == 8'd44 & go ? fsm15_out : 1'd0;
    assign incr16_left =
     fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go ? 3'd1 : 3'd0;
    assign incr16_right =
     fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go ? fsm16_out : 3'd0;
    assign incr17_left =
     fsm44_out == 8'd50 & go ? 1'd1 : 1'd0;
    assign incr17_right =
     fsm44_out == 8'd50 & go ? fsm17_out : 1'd0;
    assign incr18_left =
     fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? 3'd1 : 3'd0;
    assign incr18_right =
     fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? fsm18_out : 3'd0;
    assign incr19_left =
     fsm44_out == 8'd56 & go ? 1'd1 : 1'd0;
    assign incr19_right =
     fsm44_out == 8'd56 & go ? fsm19_out : 1'd0;
    assign incr2_left =
     fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go ? 3'd1 : 3'd0;
    assign incr2_right =
     fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go ? fsm2_out : 3'd0;
    assign incr20_left =
     fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? 3'd1 : 3'd0;
    assign incr20_right =
     fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? fsm20_out : 3'd0;
    assign incr21_left =
     fsm44_out == 8'd62 & go ? 1'd1 : 1'd0;
    assign incr21_right =
     fsm44_out == 8'd62 & go ? fsm21_out : 1'd0;
    assign incr22_left =
     fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? 3'd1 : 3'd0;
    assign incr22_right =
     fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? fsm22_out : 3'd0;
    assign incr23_left =
     fsm44_out == 8'd68 & go ? 1'd1 : 1'd0;
    assign incr23_right =
     fsm44_out == 8'd68 & go ? fsm23_out : 1'd0;
    assign incr24_left =
     fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? 3'd1 : 3'd0;
    assign incr24_right =
     fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? fsm24_out : 3'd0;
    assign incr25_left =
     fsm44_out == 8'd74 & go ? 1'd1 : 1'd0;
    assign incr25_right =
     fsm44_out == 8'd74 & go ? fsm25_out : 1'd0;
    assign incr26_left =
     fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? 3'd1 : 3'd0;
    assign incr26_right =
     fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? fsm26_out : 3'd0;
    assign incr27_left =
     fsm44_out == 8'd80 & go ? 1'd1 : 1'd0;
    assign incr27_right =
     fsm44_out == 8'd80 & go ? fsm27_out : 1'd0;
    assign incr28_left =
     fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? 3'd1 : 3'd0;
    assign incr28_right =
     fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? fsm28_out : 3'd0;
    assign incr29_left =
     fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign incr29_right =
     fsm44_out == 8'd86 & go ? fsm29_out : 1'd0;
    assign incr3_left =
     fsm44_out == 8'd8 & go ? 1'd1 : 1'd0;
    assign incr3_right =
     fsm44_out == 8'd8 & go ? fsm3_out : 1'd0;
    assign incr30_left =
     fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? 3'd1 : 3'd0;
    assign incr30_right =
     fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? fsm30_out : 3'd0;
    assign incr31_left =
     fsm44_out == 8'd92 & go ? 1'd1 : 1'd0;
    assign incr31_right =
     fsm44_out == 8'd92 & go ? fsm31_out : 1'd0;
    assign incr32_left =
     fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? 3'd1 : 3'd0;
    assign incr32_right =
     fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? fsm32_out : 3'd0;
    assign incr33_left =
     fsm44_out == 8'd98 & go ? 1'd1 : 1'd0;
    assign incr33_right =
     fsm44_out == 8'd98 & go ? fsm33_out : 1'd0;
    assign incr34_left =
     fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? 3'd1 : 3'd0;
    assign incr34_right =
     fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? fsm34_out : 3'd0;
    assign incr35_left =
     fsm44_out == 8'd104 & go ? 1'd1 : 1'd0;
    assign incr35_right =
     fsm44_out == 8'd104 & go ? fsm35_out : 1'd0;
    assign incr36_left =
     fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? 3'd1 : 3'd0;
    assign incr36_right =
     fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? fsm36_out : 3'd0;
    assign incr37_left =
     fsm44_out == 8'd110 & go ? 1'd1 : 1'd0;
    assign incr37_right =
     fsm44_out == 8'd110 & go ? fsm37_out : 1'd0;
    assign incr38_left =
     fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go ? 3'd1 : 3'd0;
    assign incr38_right =
     fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go ? fsm38_out : 3'd0;
    assign incr39_left =
     fsm44_out == 8'd116 & go ? 1'd1 : 1'd0;
    assign incr39_right =
     fsm44_out == 8'd116 & go ? fsm39_out : 1'd0;
    assign incr4_left =
     fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go ? 3'd1 : 3'd0;
    assign incr4_right =
     fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go ? fsm4_out : 3'd0;
    assign incr40_left =
     fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go ? 3'd1 : 3'd0;
    assign incr40_right =
     fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go ? fsm40_out : 3'd0;
    assign incr41_left =
     fsm44_out == 8'd122 & go ? 1'd1 : 1'd0;
    assign incr41_right =
     fsm44_out == 8'd122 & go ? fsm41_out : 1'd0;
    assign incr42_left =
     fsm44_out >= 8'd123 & fsm44_out < 8'd128 & go ? 3'd1 : 3'd0;
    assign incr42_right =
     fsm44_out >= 8'd123 & fsm44_out < 8'd128 & go ? fsm42_out : 3'd0;
    assign incr43_left =
     fsm44_out == 8'd128 & go ? 1'd1 : 1'd0;
    assign incr43_right =
     fsm44_out == 8'd128 & go ? fsm43_out : 1'd0;
    assign incr44_left =
     go ? 8'd1 : 8'd0;
    assign incr44_right =
     go ? fsm44_out : 8'd0;
    assign incr5_left =
     fsm44_out == 8'd14 & go ? 1'd1 : 1'd0;
    assign incr5_right =
     fsm44_out == 8'd14 & go ? fsm5_out : 1'd0;
    assign incr6_left =
     fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go ? 3'd1 : 3'd0;
    assign incr6_right =
     fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go ? fsm6_out : 3'd0;
    assign incr7_left =
     fsm44_out == 8'd20 & go ? 1'd1 : 1'd0;
    assign incr7_right =
     fsm44_out == 8'd20 & go ? fsm7_out : 1'd0;
    assign incr8_left =
     fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go ? 3'd1 : 3'd0;
    assign incr8_right =
     fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go ? fsm8_out : 3'd0;
    assign incr9_left =
     fsm44_out == 8'd26 & go ? 1'd1 : 1'd0;
    assign incr9_right =
     fsm44_out == 8'd26 & go ? fsm9_out : 1'd0;
    assign l0_add_left =
     fsm0_out < 1'd1 & fsm44_out == 8'd1 & go | fsm2_out < 3'd1 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go ? 4'd1 : 4'd0;
    assign l0_add_right =
     fsm0_out < 1'd1 & fsm44_out == 8'd1 & go | fsm2_out < 3'd1 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go ? l0_idx_out : 4'd0;
    assign l0_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l0_idx_in =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go ? 4'd15 :
     fsm0_out < 1'd1 & fsm44_out == 8'd1 & go | fsm2_out < 3'd1 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go ? l0_add_out : 4'd0;
    assign l0_idx_write_en =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go | fsm0_out < 1'd1 & fsm44_out == 8'd1 & go | fsm2_out < 3'd1 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go ? 1'd1 : 1'd0;
    assign l1_add_left =
     fsm2_out < 3'd1 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go ? 4'd1 : 4'd0;
    assign l1_add_right =
     fsm2_out < 3'd1 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go ? l1_idx_out : 4'd0;
    assign l1_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l1_idx_in =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go ? 4'd15 :
     fsm2_out < 3'd1 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go ? l1_add_out : 4'd0;
    assign l1_idx_write_en =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go | fsm2_out < 3'd1 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go ? 1'd1 : 1'd0;
    assign l2_add_left =
     fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? 4'd1 : 4'd0;
    assign l2_add_right =
     fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? l2_idx_out : 4'd0;
    assign l2_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l2_idx_in =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go ? 4'd15 :
     fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? l2_add_out : 4'd0;
    assign l2_idx_write_en =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? 1'd1 : 1'd0;
    assign l3_add_left =
     fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? 4'd1 : 4'd0;
    assign l3_add_right =
     fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? l3_idx_out : 4'd0;
    assign l3_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l3_idx_in =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go ? 4'd15 :
     fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? l3_add_out : 4'd0;
    assign l3_idx_write_en =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? 1'd1 : 1'd0;
    assign l4_add_left =
     fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? 4'd1 : 4'd0;
    assign l4_add_right =
     fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? l4_idx_out : 4'd0;
    assign l4_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l4_idx_in =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go ? 4'd15 :
     fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? l4_add_out : 4'd0;
    assign l4_idx_write_en =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? 1'd1 : 1'd0;
    assign l5_add_left =
     fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? 4'd1 : 4'd0;
    assign l5_add_right =
     fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? l5_idx_out : 4'd0;
    assign l5_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l5_idx_in =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go ? 4'd15 :
     fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? l5_add_out : 4'd0;
    assign l5_idx_write_en =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? 1'd1 : 1'd0;
    assign l6_add_left =
     fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd1 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? 4'd1 : 4'd0;
    assign l6_add_right =
     fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd1 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? l6_idx_out : 4'd0;
    assign l6_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l6_idx_in =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go ? 4'd15 :
     fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd1 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? l6_add_out : 4'd0;
    assign l6_idx_write_en =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd1 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? 1'd1 : 1'd0;
    assign l7_add_left =
     fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd1 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd1 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? 4'd1 : 4'd0;
    assign l7_add_right =
     fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd1 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd1 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? l7_idx_out : 4'd0;
    assign l7_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l7_idx_in =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go ? 4'd15 :
     fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd1 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd1 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? l7_add_out : 4'd0;
    assign l7_idx_write_en =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd1 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd1 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? 1'd1 : 1'd0;
    assign left_0_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_0_in =
     fsm1_out < 1'd1 & fsm44_out == 8'd2 & go | fsm3_out < 1'd1 & fsm44_out == 8'd8 & go | fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go ? l0_read_data : 32'd0;
    assign left_0_0_write_en =
     fsm1_out < 1'd1 & fsm44_out == 8'd2 & go | fsm3_out < 1'd1 & fsm44_out == 8'd8 & go | fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go ? 1'd1 : 1'd0;
    assign left_0_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_1_in =
     fsm3_out < 1'd1 & fsm44_out == 8'd8 & go | fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go ? left_0_0_out : 32'd0;
    assign left_0_1_write_en =
     fsm3_out < 1'd1 & fsm44_out == 8'd8 & go | fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go ? 1'd1 : 1'd0;
    assign left_0_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_2_in =
     fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go ? left_0_1_out : 32'd0;
    assign left_0_2_write_en =
     fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go ? 1'd1 : 1'd0;
    assign left_0_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_3_in =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? left_0_2_out : 32'd0;
    assign left_0_3_write_en =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? 1'd1 : 1'd0;
    assign left_0_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_4_in =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? left_0_3_out : 32'd0;
    assign left_0_4_write_en =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? 1'd1 : 1'd0;
    assign left_0_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_5_in =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? left_0_4_out : 32'd0;
    assign left_0_5_write_en =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? 1'd1 : 1'd0;
    assign left_0_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_6_in =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? left_0_5_out : 32'd0;
    assign left_0_6_write_en =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? 1'd1 : 1'd0;
    assign left_0_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_7_in =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? left_0_6_out : 32'd0;
    assign left_0_7_write_en =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign left_1_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_0_in =
     fsm3_out < 1'd1 & fsm44_out == 8'd8 & go | fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go ? l1_read_data : 32'd0;
    assign left_1_0_write_en =
     fsm3_out < 1'd1 & fsm44_out == 8'd8 & go | fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go ? 1'd1 : 1'd0;
    assign left_1_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_1_in =
     fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go ? left_1_0_out : 32'd0;
    assign left_1_1_write_en =
     fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go ? 1'd1 : 1'd0;
    assign left_1_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_2_in =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? left_1_1_out : 32'd0;
    assign left_1_2_write_en =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? 1'd1 : 1'd0;
    assign left_1_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_3_in =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? left_1_2_out : 32'd0;
    assign left_1_3_write_en =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? 1'd1 : 1'd0;
    assign left_1_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_4_in =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? left_1_3_out : 32'd0;
    assign left_1_4_write_en =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? 1'd1 : 1'd0;
    assign left_1_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_5_in =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? left_1_4_out : 32'd0;
    assign left_1_5_write_en =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? 1'd1 : 1'd0;
    assign left_1_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_6_in =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? left_1_5_out : 32'd0;
    assign left_1_6_write_en =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign left_1_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_7_in =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? left_1_6_out : 32'd0;
    assign left_1_7_write_en =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? 1'd1 : 1'd0;
    assign left_2_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_0_in =
     fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go ? l2_read_data : 32'd0;
    assign left_2_0_write_en =
     fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go ? 1'd1 : 1'd0;
    assign left_2_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_1_in =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? left_2_0_out : 32'd0;
    assign left_2_1_write_en =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? 1'd1 : 1'd0;
    assign left_2_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_2_in =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? left_2_1_out : 32'd0;
    assign left_2_2_write_en =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? 1'd1 : 1'd0;
    assign left_2_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_3_in =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? left_2_2_out : 32'd0;
    assign left_2_3_write_en =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? 1'd1 : 1'd0;
    assign left_2_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_4_in =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? left_2_3_out : 32'd0;
    assign left_2_4_write_en =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? 1'd1 : 1'd0;
    assign left_2_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_5_in =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? left_2_4_out : 32'd0;
    assign left_2_5_write_en =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign left_2_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_6_in =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? left_2_5_out : 32'd0;
    assign left_2_6_write_en =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? 1'd1 : 1'd0;
    assign left_2_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_7_in =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? left_2_6_out : 32'd0;
    assign left_2_7_write_en =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? 1'd1 : 1'd0;
    assign left_3_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_0_in =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? l3_read_data : 32'd0;
    assign left_3_0_write_en =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? 1'd1 : 1'd0;
    assign left_3_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_1_in =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? left_3_0_out : 32'd0;
    assign left_3_1_write_en =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? 1'd1 : 1'd0;
    assign left_3_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_2_in =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? left_3_1_out : 32'd0;
    assign left_3_2_write_en =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? 1'd1 : 1'd0;
    assign left_3_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_3_in =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? left_3_2_out : 32'd0;
    assign left_3_3_write_en =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? 1'd1 : 1'd0;
    assign left_3_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_4_in =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? left_3_3_out : 32'd0;
    assign left_3_4_write_en =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign left_3_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_5_in =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? left_3_4_out : 32'd0;
    assign left_3_5_write_en =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? 1'd1 : 1'd0;
    assign left_3_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_6_in =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? left_3_5_out : 32'd0;
    assign left_3_6_write_en =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? 1'd1 : 1'd0;
    assign left_3_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_7_in =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? left_3_6_out : 32'd0;
    assign left_3_7_write_en =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? 1'd1 : 1'd0;
    assign left_4_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_0_in =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? l4_read_data : 32'd0;
    assign left_4_0_write_en =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? 1'd1 : 1'd0;
    assign left_4_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_1_in =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? left_4_0_out : 32'd0;
    assign left_4_1_write_en =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? 1'd1 : 1'd0;
    assign left_4_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_2_in =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? left_4_1_out : 32'd0;
    assign left_4_2_write_en =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? 1'd1 : 1'd0;
    assign left_4_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_3_in =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? left_4_2_out : 32'd0;
    assign left_4_3_write_en =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign left_4_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_4_in =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? left_4_3_out : 32'd0;
    assign left_4_4_write_en =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? 1'd1 : 1'd0;
    assign left_4_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_5_in =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? left_4_4_out : 32'd0;
    assign left_4_5_write_en =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? 1'd1 : 1'd0;
    assign left_4_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_6_in =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? left_4_5_out : 32'd0;
    assign left_4_6_write_en =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? 1'd1 : 1'd0;
    assign left_4_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_7_in =
     fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go ? left_4_6_out : 32'd0;
    assign left_4_7_write_en =
     fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go ? 1'd1 : 1'd0;
    assign left_5_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_0_in =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? l5_read_data : 32'd0;
    assign left_5_0_write_en =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? 1'd1 : 1'd0;
    assign left_5_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_1_in =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? left_5_0_out : 32'd0;
    assign left_5_1_write_en =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? 1'd1 : 1'd0;
    assign left_5_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_2_in =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? left_5_1_out : 32'd0;
    assign left_5_2_write_en =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign left_5_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_3_in =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? left_5_2_out : 32'd0;
    assign left_5_3_write_en =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? 1'd1 : 1'd0;
    assign left_5_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_4_in =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? left_5_3_out : 32'd0;
    assign left_5_4_write_en =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? 1'd1 : 1'd0;
    assign left_5_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_5_in =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? left_5_4_out : 32'd0;
    assign left_5_5_write_en =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? 1'd1 : 1'd0;
    assign left_5_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_6_in =
     fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go ? left_5_5_out : 32'd0;
    assign left_5_6_write_en =
     fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go ? 1'd1 : 1'd0;
    assign left_5_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_7_in =
     fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go ? left_5_6_out : 32'd0;
    assign left_5_7_write_en =
     fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go ? 1'd1 : 1'd0;
    assign left_6_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_0_in =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? l6_read_data : 32'd0;
    assign left_6_0_write_en =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? 1'd1 : 1'd0;
    assign left_6_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_1_in =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? left_6_0_out : 32'd0;
    assign left_6_1_write_en =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign left_6_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_2_in =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? left_6_1_out : 32'd0;
    assign left_6_2_write_en =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? 1'd1 : 1'd0;
    assign left_6_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_3_in =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? left_6_2_out : 32'd0;
    assign left_6_3_write_en =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? 1'd1 : 1'd0;
    assign left_6_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_4_in =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? left_6_3_out : 32'd0;
    assign left_6_4_write_en =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? 1'd1 : 1'd0;
    assign left_6_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_5_in =
     fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go ? left_6_4_out : 32'd0;
    assign left_6_5_write_en =
     fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go ? 1'd1 : 1'd0;
    assign left_6_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_6_in =
     fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go ? left_6_5_out : 32'd0;
    assign left_6_6_write_en =
     fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go ? 1'd1 : 1'd0;
    assign left_6_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_7_in =
     fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go | fsm41_out < 1'd1 & fsm44_out == 8'd122 & go ? left_6_6_out : 32'd0;
    assign left_6_7_write_en =
     fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go | fsm41_out < 1'd1 & fsm44_out == 8'd122 & go ? 1'd1 : 1'd0;
    assign left_7_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_0_in =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? l7_read_data : 32'd0;
    assign left_7_0_write_en =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign left_7_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_1_in =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? left_7_0_out : 32'd0;
    assign left_7_1_write_en =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? 1'd1 : 1'd0;
    assign left_7_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_2_in =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? left_7_1_out : 32'd0;
    assign left_7_2_write_en =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? 1'd1 : 1'd0;
    assign left_7_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_3_in =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? left_7_2_out : 32'd0;
    assign left_7_3_write_en =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? 1'd1 : 1'd0;
    assign left_7_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_4_in =
     fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go ? left_7_3_out : 32'd0;
    assign left_7_4_write_en =
     fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go ? 1'd1 : 1'd0;
    assign left_7_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_5_in =
     fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go ? left_7_4_out : 32'd0;
    assign left_7_5_write_en =
     fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go ? 1'd1 : 1'd0;
    assign left_7_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_6_in =
     fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go | fsm41_out < 1'd1 & fsm44_out == 8'd122 & go ? left_7_5_out : 32'd0;
    assign left_7_6_write_en =
     fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go | fsm41_out < 1'd1 & fsm44_out == 8'd122 & go ? 1'd1 : 1'd0;
    assign left_7_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_7_in =
     fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go | fsm41_out < 1'd1 & fsm44_out == 8'd122 & go | fsm43_out < 1'd1 & fsm44_out == 8'd128 & go ? left_7_6_out : 32'd0;
    assign left_7_7_write_en =
     fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go | fsm41_out < 1'd1 & fsm44_out == 8'd122 & go | fsm43_out < 1'd1 & fsm44_out == 8'd128 & go ? 1'd1 : 1'd0;
    assign pe_0_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_0_go =
     fsm2_out < 3'd5 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd5 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go ? 1'd1 : 1'd0;
    assign pe_0_0_left =
     fsm2_out < 3'd5 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd5 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go ? left_0_0_out : 32'd0;
    assign pe_0_0_top =
     fsm2_out < 3'd5 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd5 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go ? top_0_0_out : 32'd0;
    assign pe_0_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_1_go =
     fsm4_out < 3'd5 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? 1'd1 : 1'd0;
    assign pe_0_1_left =
     fsm4_out < 3'd5 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? left_0_1_out : 32'd0;
    assign pe_0_1_top =
     fsm4_out < 3'd5 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? top_0_1_out : 32'd0;
    assign pe_0_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_2_go =
     fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? 1'd1 : 1'd0;
    assign pe_0_2_left =
     fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? left_0_2_out : 32'd0;
    assign pe_0_2_top =
     fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? top_0_2_out : 32'd0;
    assign pe_0_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_3_go =
     fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? 1'd1 : 1'd0;
    assign pe_0_3_left =
     fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? left_0_3_out : 32'd0;
    assign pe_0_3_top =
     fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? top_0_3_out : 32'd0;
    assign pe_0_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_4_go =
     fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? 1'd1 : 1'd0;
    assign pe_0_4_left =
     fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? left_0_4_out : 32'd0;
    assign pe_0_4_top =
     fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? top_0_4_out : 32'd0;
    assign pe_0_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_5_go =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? 1'd1 : 1'd0;
    assign pe_0_5_left =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? left_0_5_out : 32'd0;
    assign pe_0_5_top =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? top_0_5_out : 32'd0;
    assign pe_0_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_6_go =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? 1'd1 : 1'd0;
    assign pe_0_6_left =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? left_0_6_out : 32'd0;
    assign pe_0_6_top =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? top_0_6_out : 32'd0;
    assign pe_0_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_7_go =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? 1'd1 : 1'd0;
    assign pe_0_7_left =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? left_0_7_out : 32'd0;
    assign pe_0_7_top =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? top_0_7_out : 32'd0;
    assign pe_1_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_0_go =
     fsm4_out < 3'd5 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? 1'd1 : 1'd0;
    assign pe_1_0_left =
     fsm4_out < 3'd5 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? left_1_0_out : 32'd0;
    assign pe_1_0_top =
     fsm4_out < 3'd5 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? top_1_0_out : 32'd0;
    assign pe_1_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_1_go =
     fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? 1'd1 : 1'd0;
    assign pe_1_1_left =
     fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? left_1_1_out : 32'd0;
    assign pe_1_1_top =
     fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? top_1_1_out : 32'd0;
    assign pe_1_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_2_go =
     fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? 1'd1 : 1'd0;
    assign pe_1_2_left =
     fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? left_1_2_out : 32'd0;
    assign pe_1_2_top =
     fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? top_1_2_out : 32'd0;
    assign pe_1_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_3_go =
     fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? 1'd1 : 1'd0;
    assign pe_1_3_left =
     fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? left_1_3_out : 32'd0;
    assign pe_1_3_top =
     fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? top_1_3_out : 32'd0;
    assign pe_1_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_4_go =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? 1'd1 : 1'd0;
    assign pe_1_4_left =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? left_1_4_out : 32'd0;
    assign pe_1_4_top =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? top_1_4_out : 32'd0;
    assign pe_1_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_5_go =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? 1'd1 : 1'd0;
    assign pe_1_5_left =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? left_1_5_out : 32'd0;
    assign pe_1_5_top =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? top_1_5_out : 32'd0;
    assign pe_1_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_6_go =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? 1'd1 : 1'd0;
    assign pe_1_6_left =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? left_1_6_out : 32'd0;
    assign pe_1_6_top =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? top_1_6_out : 32'd0;
    assign pe_1_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_7_go =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? 1'd1 : 1'd0;
    assign pe_1_7_left =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? left_1_7_out : 32'd0;
    assign pe_1_7_top =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? top_1_7_out : 32'd0;
    assign pe_2_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_0_go =
     fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? 1'd1 : 1'd0;
    assign pe_2_0_left =
     fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? left_2_0_out : 32'd0;
    assign pe_2_0_top =
     fsm6_out < 3'd5 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? top_2_0_out : 32'd0;
    assign pe_2_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_1_go =
     fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? 1'd1 : 1'd0;
    assign pe_2_1_left =
     fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? left_2_1_out : 32'd0;
    assign pe_2_1_top =
     fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? top_2_1_out : 32'd0;
    assign pe_2_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_2_go =
     fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? 1'd1 : 1'd0;
    assign pe_2_2_left =
     fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? left_2_2_out : 32'd0;
    assign pe_2_2_top =
     fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? top_2_2_out : 32'd0;
    assign pe_2_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_3_go =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? 1'd1 : 1'd0;
    assign pe_2_3_left =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? left_2_3_out : 32'd0;
    assign pe_2_3_top =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? top_2_3_out : 32'd0;
    assign pe_2_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_4_go =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? 1'd1 : 1'd0;
    assign pe_2_4_left =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? left_2_4_out : 32'd0;
    assign pe_2_4_top =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? top_2_4_out : 32'd0;
    assign pe_2_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_5_go =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? 1'd1 : 1'd0;
    assign pe_2_5_left =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? left_2_5_out : 32'd0;
    assign pe_2_5_top =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? top_2_5_out : 32'd0;
    assign pe_2_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_6_go =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? 1'd1 : 1'd0;
    assign pe_2_6_left =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? left_2_6_out : 32'd0;
    assign pe_2_6_top =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? top_2_6_out : 32'd0;
    assign pe_2_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_7_go =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? 1'd1 : 1'd0;
    assign pe_2_7_left =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? left_2_7_out : 32'd0;
    assign pe_2_7_top =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? top_2_7_out : 32'd0;
    assign pe_3_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_0_go =
     fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? 1'd1 : 1'd0;
    assign pe_3_0_left =
     fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? left_3_0_out : 32'd0;
    assign pe_3_0_top =
     fsm8_out < 3'd5 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? top_3_0_out : 32'd0;
    assign pe_3_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_1_go =
     fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? 1'd1 : 1'd0;
    assign pe_3_1_left =
     fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? left_3_1_out : 32'd0;
    assign pe_3_1_top =
     fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? top_3_1_out : 32'd0;
    assign pe_3_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_2_go =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? 1'd1 : 1'd0;
    assign pe_3_2_left =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? left_3_2_out : 32'd0;
    assign pe_3_2_top =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? top_3_2_out : 32'd0;
    assign pe_3_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_3_go =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? 1'd1 : 1'd0;
    assign pe_3_3_left =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? left_3_3_out : 32'd0;
    assign pe_3_3_top =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? top_3_3_out : 32'd0;
    assign pe_3_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_4_go =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? 1'd1 : 1'd0;
    assign pe_3_4_left =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? left_3_4_out : 32'd0;
    assign pe_3_4_top =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? top_3_4_out : 32'd0;
    assign pe_3_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_5_go =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? 1'd1 : 1'd0;
    assign pe_3_5_left =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? left_3_5_out : 32'd0;
    assign pe_3_5_top =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? top_3_5_out : 32'd0;
    assign pe_3_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_6_go =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? 1'd1 : 1'd0;
    assign pe_3_6_left =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? left_3_6_out : 32'd0;
    assign pe_3_6_top =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? top_3_6_out : 32'd0;
    assign pe_3_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_7_go =
     fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? 1'd1 : 1'd0;
    assign pe_3_7_left =
     fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? left_3_7_out : 32'd0;
    assign pe_3_7_top =
     fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? top_3_7_out : 32'd0;
    assign pe_4_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_0_go =
     fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? 1'd1 : 1'd0;
    assign pe_4_0_left =
     fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? left_4_0_out : 32'd0;
    assign pe_4_0_top =
     fsm10_out < 3'd5 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? top_4_0_out : 32'd0;
    assign pe_4_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_1_go =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? 1'd1 : 1'd0;
    assign pe_4_1_left =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? left_4_1_out : 32'd0;
    assign pe_4_1_top =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? top_4_1_out : 32'd0;
    assign pe_4_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_2_go =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? 1'd1 : 1'd0;
    assign pe_4_2_left =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? left_4_2_out : 32'd0;
    assign pe_4_2_top =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? top_4_2_out : 32'd0;
    assign pe_4_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_3_go =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? 1'd1 : 1'd0;
    assign pe_4_3_left =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? left_4_3_out : 32'd0;
    assign pe_4_3_top =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? top_4_3_out : 32'd0;
    assign pe_4_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_4_go =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? 1'd1 : 1'd0;
    assign pe_4_4_left =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? left_4_4_out : 32'd0;
    assign pe_4_4_top =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? top_4_4_out : 32'd0;
    assign pe_4_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_5_go =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? 1'd1 : 1'd0;
    assign pe_4_5_left =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? left_4_5_out : 32'd0;
    assign pe_4_5_top =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? top_4_5_out : 32'd0;
    assign pe_4_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_6_go =
     fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? 1'd1 : 1'd0;
    assign pe_4_6_left =
     fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? left_4_6_out : 32'd0;
    assign pe_4_6_top =
     fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? top_4_6_out : 32'd0;
    assign pe_4_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_7_go =
     fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go ? 1'd1 : 1'd0;
    assign pe_4_7_left =
     fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go ? left_4_7_out : 32'd0;
    assign pe_4_7_top =
     fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go ? top_4_7_out : 32'd0;
    assign pe_5_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_0_go =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? 1'd1 : 1'd0;
    assign pe_5_0_left =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? left_5_0_out : 32'd0;
    assign pe_5_0_top =
     fsm12_out < 3'd5 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? top_5_0_out : 32'd0;
    assign pe_5_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_1_go =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? 1'd1 : 1'd0;
    assign pe_5_1_left =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? left_5_1_out : 32'd0;
    assign pe_5_1_top =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? top_5_1_out : 32'd0;
    assign pe_5_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_2_go =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? 1'd1 : 1'd0;
    assign pe_5_2_left =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? left_5_2_out : 32'd0;
    assign pe_5_2_top =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? top_5_2_out : 32'd0;
    assign pe_5_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_3_go =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? 1'd1 : 1'd0;
    assign pe_5_3_left =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? left_5_3_out : 32'd0;
    assign pe_5_3_top =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? top_5_3_out : 32'd0;
    assign pe_5_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_4_go =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? 1'd1 : 1'd0;
    assign pe_5_4_left =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? left_5_4_out : 32'd0;
    assign pe_5_4_top =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? top_5_4_out : 32'd0;
    assign pe_5_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_5_go =
     fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? 1'd1 : 1'd0;
    assign pe_5_5_left =
     fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? left_5_5_out : 32'd0;
    assign pe_5_5_top =
     fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? top_5_5_out : 32'd0;
    assign pe_5_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_6_go =
     fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go ? 1'd1 : 1'd0;
    assign pe_5_6_left =
     fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go ? left_5_6_out : 32'd0;
    assign pe_5_6_top =
     fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go ? top_5_6_out : 32'd0;
    assign pe_5_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_7_go =
     fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go ? 1'd1 : 1'd0;
    assign pe_5_7_left =
     fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go ? left_5_7_out : 32'd0;
    assign pe_5_7_top =
     fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go ? top_5_7_out : 32'd0;
    assign pe_6_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_0_go =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? 1'd1 : 1'd0;
    assign pe_6_0_left =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? left_6_0_out : 32'd0;
    assign pe_6_0_top =
     fsm14_out < 3'd5 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? top_6_0_out : 32'd0;
    assign pe_6_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_1_go =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? 1'd1 : 1'd0;
    assign pe_6_1_left =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? left_6_1_out : 32'd0;
    assign pe_6_1_top =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? top_6_1_out : 32'd0;
    assign pe_6_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_2_go =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? 1'd1 : 1'd0;
    assign pe_6_2_left =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? left_6_2_out : 32'd0;
    assign pe_6_2_top =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? top_6_2_out : 32'd0;
    assign pe_6_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_3_go =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? 1'd1 : 1'd0;
    assign pe_6_3_left =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? left_6_3_out : 32'd0;
    assign pe_6_3_top =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? top_6_3_out : 32'd0;
    assign pe_6_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_4_go =
     fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? 1'd1 : 1'd0;
    assign pe_6_4_left =
     fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? left_6_4_out : 32'd0;
    assign pe_6_4_top =
     fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? top_6_4_out : 32'd0;
    assign pe_6_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_5_go =
     fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go ? 1'd1 : 1'd0;
    assign pe_6_5_left =
     fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go ? left_6_5_out : 32'd0;
    assign pe_6_5_top =
     fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go ? top_6_5_out : 32'd0;
    assign pe_6_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_6_go =
     fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go ? 1'd1 : 1'd0;
    assign pe_6_6_left =
     fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go ? left_6_6_out : 32'd0;
    assign pe_6_6_top =
     fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go ? top_6_6_out : 32'd0;
    assign pe_6_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_7_go =
     fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go | fsm42_out < 3'd5 & fsm44_out >= 8'd123 & fsm44_out < 8'd128 & go ? 1'd1 : 1'd0;
    assign pe_6_7_left =
     fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go | fsm42_out < 3'd5 & fsm44_out >= 8'd123 & fsm44_out < 8'd128 & go ? left_6_7_out : 32'd0;
    assign pe_6_7_top =
     fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go | fsm42_out < 3'd5 & fsm44_out >= 8'd123 & fsm44_out < 8'd128 & go ? top_6_7_out : 32'd0;
    assign pe_7_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_0_go =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? 1'd1 : 1'd0;
    assign pe_7_0_left =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? left_7_0_out : 32'd0;
    assign pe_7_0_top =
     fsm16_out < 3'd5 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go ? top_7_0_out : 32'd0;
    assign pe_7_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_1_go =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? 1'd1 : 1'd0;
    assign pe_7_1_left =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? left_7_1_out : 32'd0;
    assign pe_7_1_top =
     fsm18_out < 3'd5 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go ? top_7_1_out : 32'd0;
    assign pe_7_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_2_go =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? 1'd1 : 1'd0;
    assign pe_7_2_left =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? left_7_2_out : 32'd0;
    assign pe_7_2_top =
     fsm20_out < 3'd5 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go ? top_7_2_out : 32'd0;
    assign pe_7_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_3_go =
     fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? 1'd1 : 1'd0;
    assign pe_7_3_left =
     fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? left_7_3_out : 32'd0;
    assign pe_7_3_top =
     fsm22_out < 3'd5 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go ? top_7_3_out : 32'd0;
    assign pe_7_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_4_go =
     fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go ? 1'd1 : 1'd0;
    assign pe_7_4_left =
     fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go ? left_7_4_out : 32'd0;
    assign pe_7_4_top =
     fsm24_out < 3'd5 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go ? top_7_4_out : 32'd0;
    assign pe_7_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_5_go =
     fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go ? 1'd1 : 1'd0;
    assign pe_7_5_left =
     fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go ? left_7_5_out : 32'd0;
    assign pe_7_5_top =
     fsm26_out < 3'd5 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go ? top_7_5_out : 32'd0;
    assign pe_7_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_6_go =
     fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go | fsm42_out < 3'd5 & fsm44_out >= 8'd123 & fsm44_out < 8'd128 & go ? 1'd1 : 1'd0;
    assign pe_7_6_left =
     fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go | fsm42_out < 3'd5 & fsm44_out >= 8'd123 & fsm44_out < 8'd128 & go ? left_7_6_out : 32'd0;
    assign pe_7_6_top =
     fsm28_out < 3'd5 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go | fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go | fsm42_out < 3'd5 & fsm44_out >= 8'd123 & fsm44_out < 8'd128 & go ? top_7_6_out : 32'd0;
    assign pe_7_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_7_go =
     fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go | fsm42_out < 3'd5 & fsm44_out >= 8'd123 & fsm44_out < 8'd128 & go | fsm44_out >= 8'd129 & fsm44_out < 8'd134 & go ? 1'd1 : 1'd0;
    assign pe_7_7_left =
     fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go | fsm42_out < 3'd5 & fsm44_out >= 8'd123 & fsm44_out < 8'd128 & go | fsm44_out >= 8'd129 & fsm44_out < 8'd134 & go ? left_7_7_out : 32'd0;
    assign pe_7_7_top =
     fsm30_out < 3'd5 & fsm44_out >= 8'd87 & fsm44_out < 8'd92 & go | fsm32_out < 3'd5 & fsm44_out >= 8'd93 & fsm44_out < 8'd98 & go | fsm34_out < 3'd5 & fsm44_out >= 8'd99 & fsm44_out < 8'd104 & go | fsm36_out < 3'd5 & fsm44_out >= 8'd105 & fsm44_out < 8'd110 & go | fsm38_out < 3'd5 & fsm44_out >= 8'd111 & fsm44_out < 8'd116 & go | fsm40_out < 3'd5 & fsm44_out >= 8'd117 & fsm44_out < 8'd122 & go | fsm42_out < 3'd5 & fsm44_out >= 8'd123 & fsm44_out < 8'd128 & go | fsm44_out >= 8'd129 & fsm44_out < 8'd134 & go ? top_7_7_out : 32'd0;
    assign t0_add_left =
     fsm0_out < 1'd1 & fsm44_out == 8'd1 & go | fsm2_out < 3'd1 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go ? 4'd1 : 4'd0;
    assign t0_add_right =
     fsm0_out < 1'd1 & fsm44_out == 8'd1 & go | fsm2_out < 3'd1 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go ? t0_idx_out : 4'd0;
    assign t0_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t0_idx_in =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go ? 4'd15 :
     fsm0_out < 1'd1 & fsm44_out == 8'd1 & go | fsm2_out < 3'd1 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go ? t0_add_out : 4'd0;
    assign t0_idx_write_en =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go | fsm0_out < 1'd1 & fsm44_out == 8'd1 & go | fsm2_out < 3'd1 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go ? 1'd1 : 1'd0;
    assign t1_add_left =
     fsm2_out < 3'd1 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go ? 4'd1 : 4'd0;
    assign t1_add_right =
     fsm2_out < 3'd1 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go ? t1_idx_out : 4'd0;
    assign t1_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t1_idx_in =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go ? 4'd15 :
     fsm2_out < 3'd1 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go ? t1_add_out : 4'd0;
    assign t1_idx_write_en =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go | fsm2_out < 3'd1 & fsm44_out >= 8'd3 & fsm44_out < 8'd8 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go ? 1'd1 : 1'd0;
    assign t2_add_left =
     fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? 4'd1 : 4'd0;
    assign t2_add_right =
     fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? t2_idx_out : 4'd0;
    assign t2_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t2_idx_in =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go ? 4'd15 :
     fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? t2_add_out : 4'd0;
    assign t2_idx_write_en =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go | fsm4_out < 3'd1 & fsm44_out >= 8'd9 & fsm44_out < 8'd14 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go ? 1'd1 : 1'd0;
    assign t3_add_left =
     fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? 4'd1 : 4'd0;
    assign t3_add_right =
     fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? t3_idx_out : 4'd0;
    assign t3_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t3_idx_in =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go ? 4'd15 :
     fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? t3_add_out : 4'd0;
    assign t3_idx_write_en =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go | fsm6_out < 3'd1 & fsm44_out >= 8'd15 & fsm44_out < 8'd20 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go ? 1'd1 : 1'd0;
    assign t4_add_left =
     fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? 4'd1 : 4'd0;
    assign t4_add_right =
     fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? t4_idx_out : 4'd0;
    assign t4_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t4_idx_in =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go ? 4'd15 :
     fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? t4_add_out : 4'd0;
    assign t4_idx_write_en =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go | fsm8_out < 3'd1 & fsm44_out >= 8'd21 & fsm44_out < 8'd26 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go ? 1'd1 : 1'd0;
    assign t5_add_left =
     fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? 4'd1 : 4'd0;
    assign t5_add_right =
     fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? t5_idx_out : 4'd0;
    assign t5_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t5_idx_in =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go ? 4'd15 :
     fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? t5_add_out : 4'd0;
    assign t5_idx_write_en =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go | fsm10_out < 3'd1 & fsm44_out >= 8'd27 & fsm44_out < 8'd32 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go ? 1'd1 : 1'd0;
    assign t6_add_left =
     fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd1 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? 4'd1 : 4'd0;
    assign t6_add_right =
     fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd1 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? t6_idx_out : 4'd0;
    assign t6_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t6_idx_in =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go ? 4'd15 :
     fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd1 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? t6_add_out : 4'd0;
    assign t6_idx_write_en =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go | fsm12_out < 3'd1 & fsm44_out >= 8'd33 & fsm44_out < 8'd38 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd1 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go ? 1'd1 : 1'd0;
    assign t7_add_left =
     fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd1 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd1 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? 4'd1 : 4'd0;
    assign t7_add_right =
     fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd1 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd1 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? t7_idx_out : 4'd0;
    assign t7_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t7_idx_in =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go ? 4'd15 :
     fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd1 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd1 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? t7_add_out : 4'd0;
    assign t7_idx_write_en =
     fsm_out < 1'd1 & fsm44_out == 8'd0 & go | fsm14_out < 3'd1 & fsm44_out >= 8'd39 & fsm44_out < 8'd44 & go | fsm16_out < 3'd1 & fsm44_out >= 8'd45 & fsm44_out < 8'd50 & go | fsm18_out < 3'd1 & fsm44_out >= 8'd51 & fsm44_out < 8'd56 & go | fsm20_out < 3'd1 & fsm44_out >= 8'd57 & fsm44_out < 8'd62 & go | fsm22_out < 3'd1 & fsm44_out >= 8'd63 & fsm44_out < 8'd68 & go | fsm24_out < 3'd1 & fsm44_out >= 8'd69 & fsm44_out < 8'd74 & go | fsm26_out < 3'd1 & fsm44_out >= 8'd75 & fsm44_out < 8'd80 & go | fsm28_out < 3'd1 & fsm44_out >= 8'd81 & fsm44_out < 8'd86 & go ? 1'd1 : 1'd0;
    assign top_0_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_0_in =
     fsm1_out < 1'd1 & fsm44_out == 8'd2 & go | fsm3_out < 1'd1 & fsm44_out == 8'd8 & go | fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go ? t0_read_data : 32'd0;
    assign top_0_0_write_en =
     fsm1_out < 1'd1 & fsm44_out == 8'd2 & go | fsm3_out < 1'd1 & fsm44_out == 8'd8 & go | fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go ? 1'd1 : 1'd0;
    assign top_0_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_1_in =
     fsm3_out < 1'd1 & fsm44_out == 8'd8 & go | fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go ? t1_read_data : 32'd0;
    assign top_0_1_write_en =
     fsm3_out < 1'd1 & fsm44_out == 8'd8 & go | fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go ? 1'd1 : 1'd0;
    assign top_0_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_2_in =
     fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go ? t2_read_data : 32'd0;
    assign top_0_2_write_en =
     fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go ? 1'd1 : 1'd0;
    assign top_0_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_3_in =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? t3_read_data : 32'd0;
    assign top_0_3_write_en =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? 1'd1 : 1'd0;
    assign top_0_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_4_in =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? t4_read_data : 32'd0;
    assign top_0_4_write_en =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? 1'd1 : 1'd0;
    assign top_0_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_5_in =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? t5_read_data : 32'd0;
    assign top_0_5_write_en =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? 1'd1 : 1'd0;
    assign top_0_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_6_in =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? t6_read_data : 32'd0;
    assign top_0_6_write_en =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? 1'd1 : 1'd0;
    assign top_0_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_7_in =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? t7_read_data : 32'd0;
    assign top_0_7_write_en =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign top_1_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_0_in =
     fsm3_out < 1'd1 & fsm44_out == 8'd8 & go | fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go ? top_0_0_out : 32'd0;
    assign top_1_0_write_en =
     fsm3_out < 1'd1 & fsm44_out == 8'd8 & go | fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go ? 1'd1 : 1'd0;
    assign top_1_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_1_in =
     fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go ? top_0_1_out : 32'd0;
    assign top_1_1_write_en =
     fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go ? 1'd1 : 1'd0;
    assign top_1_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_2_in =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? top_0_2_out : 32'd0;
    assign top_1_2_write_en =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? 1'd1 : 1'd0;
    assign top_1_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_3_in =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? top_0_3_out : 32'd0;
    assign top_1_3_write_en =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? 1'd1 : 1'd0;
    assign top_1_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_4_in =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? top_0_4_out : 32'd0;
    assign top_1_4_write_en =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? 1'd1 : 1'd0;
    assign top_1_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_5_in =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? top_0_5_out : 32'd0;
    assign top_1_5_write_en =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? 1'd1 : 1'd0;
    assign top_1_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_6_in =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? top_0_6_out : 32'd0;
    assign top_1_6_write_en =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign top_1_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_7_in =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? top_0_7_out : 32'd0;
    assign top_1_7_write_en =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? 1'd1 : 1'd0;
    assign top_2_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_0_in =
     fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go ? top_1_0_out : 32'd0;
    assign top_2_0_write_en =
     fsm5_out < 1'd1 & fsm44_out == 8'd14 & go | fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go ? 1'd1 : 1'd0;
    assign top_2_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_1_in =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? top_1_1_out : 32'd0;
    assign top_2_1_write_en =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? 1'd1 : 1'd0;
    assign top_2_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_2_in =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? top_1_2_out : 32'd0;
    assign top_2_2_write_en =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? 1'd1 : 1'd0;
    assign top_2_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_3_in =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? top_1_3_out : 32'd0;
    assign top_2_3_write_en =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? 1'd1 : 1'd0;
    assign top_2_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_4_in =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? top_1_4_out : 32'd0;
    assign top_2_4_write_en =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? 1'd1 : 1'd0;
    assign top_2_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_5_in =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? top_1_5_out : 32'd0;
    assign top_2_5_write_en =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign top_2_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_6_in =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? top_1_6_out : 32'd0;
    assign top_2_6_write_en =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? 1'd1 : 1'd0;
    assign top_2_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_7_in =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? top_1_7_out : 32'd0;
    assign top_2_7_write_en =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? 1'd1 : 1'd0;
    assign top_3_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_0_in =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? top_2_0_out : 32'd0;
    assign top_3_0_write_en =
     fsm7_out < 1'd1 & fsm44_out == 8'd20 & go | fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go ? 1'd1 : 1'd0;
    assign top_3_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_1_in =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? top_2_1_out : 32'd0;
    assign top_3_1_write_en =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? 1'd1 : 1'd0;
    assign top_3_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_2_in =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? top_2_2_out : 32'd0;
    assign top_3_2_write_en =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? 1'd1 : 1'd0;
    assign top_3_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_3_in =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? top_2_3_out : 32'd0;
    assign top_3_3_write_en =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? 1'd1 : 1'd0;
    assign top_3_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_4_in =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? top_2_4_out : 32'd0;
    assign top_3_4_write_en =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign top_3_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_5_in =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? top_2_5_out : 32'd0;
    assign top_3_5_write_en =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? 1'd1 : 1'd0;
    assign top_3_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_6_in =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? top_2_6_out : 32'd0;
    assign top_3_6_write_en =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? 1'd1 : 1'd0;
    assign top_3_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_7_in =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? top_2_7_out : 32'd0;
    assign top_3_7_write_en =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? 1'd1 : 1'd0;
    assign top_4_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_0_in =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? top_3_0_out : 32'd0;
    assign top_4_0_write_en =
     fsm9_out < 1'd1 & fsm44_out == 8'd26 & go | fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go ? 1'd1 : 1'd0;
    assign top_4_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_1_in =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? top_3_1_out : 32'd0;
    assign top_4_1_write_en =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? 1'd1 : 1'd0;
    assign top_4_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_2_in =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? top_3_2_out : 32'd0;
    assign top_4_2_write_en =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? 1'd1 : 1'd0;
    assign top_4_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_3_in =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? top_3_3_out : 32'd0;
    assign top_4_3_write_en =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign top_4_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_4_in =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? top_3_4_out : 32'd0;
    assign top_4_4_write_en =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? 1'd1 : 1'd0;
    assign top_4_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_5_in =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? top_3_5_out : 32'd0;
    assign top_4_5_write_en =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? 1'd1 : 1'd0;
    assign top_4_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_6_in =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? top_3_6_out : 32'd0;
    assign top_4_6_write_en =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? 1'd1 : 1'd0;
    assign top_4_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_7_in =
     fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go ? top_3_7_out : 32'd0;
    assign top_4_7_write_en =
     fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go ? 1'd1 : 1'd0;
    assign top_5_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_0_in =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? top_4_0_out : 32'd0;
    assign top_5_0_write_en =
     fsm11_out < 1'd1 & fsm44_out == 8'd32 & go | fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go ? 1'd1 : 1'd0;
    assign top_5_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_1_in =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? top_4_1_out : 32'd0;
    assign top_5_1_write_en =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? 1'd1 : 1'd0;
    assign top_5_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_2_in =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? top_4_2_out : 32'd0;
    assign top_5_2_write_en =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign top_5_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_3_in =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? top_4_3_out : 32'd0;
    assign top_5_3_write_en =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? 1'd1 : 1'd0;
    assign top_5_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_4_in =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? top_4_4_out : 32'd0;
    assign top_5_4_write_en =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? 1'd1 : 1'd0;
    assign top_5_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_5_in =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? top_4_5_out : 32'd0;
    assign top_5_5_write_en =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? 1'd1 : 1'd0;
    assign top_5_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_6_in =
     fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go ? top_4_6_out : 32'd0;
    assign top_5_6_write_en =
     fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go ? 1'd1 : 1'd0;
    assign top_5_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_7_in =
     fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go ? top_4_7_out : 32'd0;
    assign top_5_7_write_en =
     fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go ? 1'd1 : 1'd0;
    assign top_6_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_0_in =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? top_5_0_out : 32'd0;
    assign top_6_0_write_en =
     fsm13_out < 1'd1 & fsm44_out == 8'd38 & go | fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go ? 1'd1 : 1'd0;
    assign top_6_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_1_in =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? top_5_1_out : 32'd0;
    assign top_6_1_write_en =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign top_6_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_2_in =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? top_5_2_out : 32'd0;
    assign top_6_2_write_en =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? 1'd1 : 1'd0;
    assign top_6_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_3_in =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? top_5_3_out : 32'd0;
    assign top_6_3_write_en =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? 1'd1 : 1'd0;
    assign top_6_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_4_in =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? top_5_4_out : 32'd0;
    assign top_6_4_write_en =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? 1'd1 : 1'd0;
    assign top_6_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_5_in =
     fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go ? top_5_5_out : 32'd0;
    assign top_6_5_write_en =
     fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go ? 1'd1 : 1'd0;
    assign top_6_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_6_in =
     fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go ? top_5_6_out : 32'd0;
    assign top_6_6_write_en =
     fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go ? 1'd1 : 1'd0;
    assign top_6_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_7_in =
     fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go | fsm41_out < 1'd1 & fsm44_out == 8'd122 & go ? top_5_7_out : 32'd0;
    assign top_6_7_write_en =
     fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go | fsm41_out < 1'd1 & fsm44_out == 8'd122 & go ? 1'd1 : 1'd0;
    assign top_7_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_0_in =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? top_6_0_out : 32'd0;
    assign top_7_0_write_en =
     fsm15_out < 1'd1 & fsm44_out == 8'd44 & go | fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go ? 1'd1 : 1'd0;
    assign top_7_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_1_in =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? top_6_1_out : 32'd0;
    assign top_7_1_write_en =
     fsm17_out < 1'd1 & fsm44_out == 8'd50 & go | fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go ? 1'd1 : 1'd0;
    assign top_7_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_2_in =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? top_6_2_out : 32'd0;
    assign top_7_2_write_en =
     fsm19_out < 1'd1 & fsm44_out == 8'd56 & go | fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go ? 1'd1 : 1'd0;
    assign top_7_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_3_in =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? top_6_3_out : 32'd0;
    assign top_7_3_write_en =
     fsm21_out < 1'd1 & fsm44_out == 8'd62 & go | fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go ? 1'd1 : 1'd0;
    assign top_7_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_4_in =
     fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go ? top_6_4_out : 32'd0;
    assign top_7_4_write_en =
     fsm23_out < 1'd1 & fsm44_out == 8'd68 & go | fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go ? 1'd1 : 1'd0;
    assign top_7_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_5_in =
     fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go ? top_6_5_out : 32'd0;
    assign top_7_5_write_en =
     fsm25_out < 1'd1 & fsm44_out == 8'd74 & go | fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go ? 1'd1 : 1'd0;
    assign top_7_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_6_in =
     fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go | fsm41_out < 1'd1 & fsm44_out == 8'd122 & go ? top_6_6_out : 32'd0;
    assign top_7_6_write_en =
     fsm27_out < 1'd1 & fsm44_out == 8'd80 & go | fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go | fsm41_out < 1'd1 & fsm44_out == 8'd122 & go ? 1'd1 : 1'd0;
    assign top_7_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_7_in =
     fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go | fsm41_out < 1'd1 & fsm44_out == 8'd122 & go | fsm43_out < 1'd1 & fsm44_out == 8'd128 & go ? top_6_7_out : 32'd0;
    assign top_7_7_write_en =
     fsm29_out < 1'd1 & fsm44_out == 8'd86 & go | fsm31_out < 1'd1 & fsm44_out == 8'd92 & go | fsm33_out < 1'd1 & fsm44_out == 8'd98 & go | fsm35_out < 1'd1 & fsm44_out == 8'd104 & go | fsm37_out < 1'd1 & fsm44_out == 8'd110 & go | fsm39_out < 1'd1 & fsm44_out == 8'd116 & go | fsm41_out < 1'd1 & fsm44_out == 8'd122 & go | fsm43_out < 1'd1 & fsm44_out == 8'd128 & go ? 1'd1 : 1'd0;
endmodule

module mac_pe (
    input logic [31:0] top,
    input logic [31:0] left,
    output logic [31:0] out,
    input logic go,
    input logic clk,
    output logic done
);
    logic [31:0] acc_in;
    logic acc_write_en;
    logic acc_clk;
    logic [31:0] acc_out;
    logic acc_done;
    logic [31:0] mul_reg_in;
    logic mul_reg_write_en;
    logic mul_reg_clk;
    logic [31:0] mul_reg_out;
    logic mul_reg_done;
    logic [31:0] add_left;
    logic [31:0] add_right;
    logic [31:0] add_out;
    logic mul_clk;
    logic mul_go;
    logic [31:0] mul_left;
    logic [31:0] mul_right;
    logic [31:0] mul_out;
    logic mul_done;
    logic [2:0] fsm_in;
    logic fsm_write_en;
    logic fsm_clk;
    logic [2:0] fsm_out;
    logic fsm_done;
    logic [2:0] incr_left;
    logic [2:0] incr_right;
    logic [2:0] incr_out;
    initial begin
        acc_in = 32'd0;
        acc_write_en = 1'd0;
        acc_clk = 1'd0;
        mul_reg_in = 32'd0;
        mul_reg_write_en = 1'd0;
        mul_reg_clk = 1'd0;
        add_left = 32'd0;
        add_right = 32'd0;
        mul_clk = 1'd0;
        mul_go = 1'd0;
        mul_left = 32'd0;
        mul_right = 32'd0;
        fsm_in = 3'd0;
        fsm_write_en = 1'd0;
        fsm_clk = 1'd0;
        incr_left = 3'd0;
        incr_right = 3'd0;
    end
    std_reg # (
        .width(32)
    ) acc (
        .clk(acc_clk),
        .done(acc_done),
        .in(acc_in),
        .out(acc_out),
        .write_en(acc_write_en)
    );
    std_reg # (
        .width(32)
    ) mul_reg (
        .clk(mul_reg_clk),
        .done(mul_reg_done),
        .in(mul_reg_in),
        .out(mul_reg_out),
        .write_en(mul_reg_write_en)
    );
    std_add # (
        .width(32)
    ) add (
        .left(add_left),
        .out(add_out),
        .right(add_right)
    );
    std_mult_pipe # (
        .width(32)
    ) mul (
        .clk(mul_clk),
        .done(mul_done),
        .go(mul_go),
        .left(mul_left),
        .out(mul_out),
        .right(mul_right)
    );
    std_reg # (
        .width(3)
    ) fsm (
        .clk(fsm_clk),
        .done(fsm_done),
        .in(fsm_in),
        .out(fsm_out),
        .write_en(fsm_write_en)
    );
    std_add # (
        .width(3)
    ) incr (
        .left(incr_left),
        .out(incr_out),
        .right(incr_right)
    );
    assign done =
     fsm_out == 3'd5 ? 1'd1 : 1'd0;
    assign out =
     1'b1 ? acc_out : 32'd0;
    assign acc_clk =
     1'b1 ? clk : 1'd0;
    assign acc_in =
     fsm_out == 3'd4 & go ? add_out : 32'd0;
    assign acc_write_en =
     fsm_out == 3'd4 & go ? 1'd1 : 1'd0;
    assign add_left =
     fsm_out == 3'd4 & go ? acc_out : 32'd0;
    assign add_right =
     fsm_out == 3'd4 & go ? mul_reg_out : 32'd0;
    assign fsm_clk =
     1'b1 ? clk : 1'd0;
    assign fsm_in =
     fsm_out == 3'd5 ? 3'd0 :
     fsm_out != 3'd5 & go ? incr_out : 3'd0;
    assign fsm_write_en =
     fsm_out != 3'd5 & go | fsm_out == 3'd5 ? 1'd1 : 1'd0;
    assign incr_left =
     go ? 3'd1 : 3'd0;
    assign incr_right =
     go ? fsm_out : 3'd0;
    assign mul_clk =
     1'b1 ? clk : 1'd0;
    assign mul_go =
     ~mul_done & fsm_out < 3'd4 & go ? 1'd1 : 1'd0;
    assign mul_left =
     fsm_out < 3'd4 & go ? top : 32'd0;
    assign mul_right =
     fsm_out < 3'd4 & go ? left : 32'd0;
    assign mul_reg_clk =
     1'b1 ? clk : 1'd0;
    assign mul_reg_in =
     mul_done & fsm_out < 3'd4 & go ? mul_out : 32'd0;
    assign mul_reg_write_en =
     mul_done & fsm_out < 3'd4 & go ? 1'd1 : 1'd0;
endmodule
