
/// This is mostly used for testing the static guarantees currently.
/// A realistic implementation would probably take four cycles.
module pipelined_mult (
    input wire clk,
    input wire reset,
    // inputs
    input wire [31:0] left,
    input wire [31:0] right,
    // The input has been committed
    output wire [31:0] out
);

logic [31:0] lt, rt, buff0, buff1, buff2, tmp_prod;

assign out = buff2;
assign tmp_prod = lt * rt;

always_ff @(posedge clk) begin
    if (reset) begin
        lt <= 0;
        rt <= 0;
        buff0 <= 0;
        buff1 <= 0;
        buff2 <= 0;
    end else begin
        lt <= left;
        rt <= right;
        buff0 <= tmp_prod;
        buff1 <= buff0;
        buff2 <= buff1;
    end
end

endmodule

module bb_pipelined_mult(
	               input wire [31:0] left,
	               input wire [31:0] right,
	               output wire [31:0] out,
	               input wire clk
	               );
`ifdef __ICARUS__
   reg [31:0] reg0;
   reg [31:0] reg1;
   reg [31:0] reg2;
   reg [31:0] reg3;
   always @( posedge clk ) begin
      reg0 <= left * right;
      reg1 <= reg0;
      reg2 <= reg1;
      reg3 <= reg2;
   end
   assign out = reg3;
`elsif VERILATOR
   reg [31:0] reg0;
   reg [31:0] reg1;
   reg [31:0] reg2;
   reg [31:0] reg3;
   always @( posedge clk ) begin
      reg0 <= left * right;
      reg1 <= reg0;
      reg2 <= reg1;
      reg3 <= reg2;
   end
   assign out = reg3;
`else
   // mul_uint32 is a black box module generated by Xilinx's IP Core generator.
   // Generation commands are in the synth.tcl file.
   mul_uint32 mul_uint32 (
                   .A(left),
                   .B(right),
                   .P(out),
                   .CLK(clk)
                   );
`endif
endmodule
/* verilator lint_off MULTITOP */
/// =================== Unsigned, Fixed Point =========================
module std_fp_add #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  assign out = left + right;
endmodule

module std_fp_sub #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module std_fp_mult_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16,
    parameter SIGNED = 0
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    input  logic             go,
    input  logic             clk,
    input  logic             reset,
    output logic [WIDTH-1:0] out,
    output logic             done
);
  logic [WIDTH-1:0]          rtmp;
  logic [WIDTH-1:0]          ltmp;
  logic [(WIDTH << 1) - 1:0] out_tmp;
  // Buffer used to walk through the 3 cycles of the pipeline.
  logic done_buf[1:0];

  assign done = done_buf[1];

  assign out = out_tmp[(WIDTH << 1) - INT_WIDTH - 1 : WIDTH - INT_WIDTH];

  // If the done buffer is completely empty and go is high then execution
  // just started.
  logic start;
  assign start = go;

  // Start sending the done signal.
  always_ff @(posedge clk) begin
    if (start)
      done_buf[0] <= 1;
    else
      done_buf[0] <= 0;
  end

  // Push the done signal through the pipeline.
  always_ff @(posedge clk) begin
    if (go) begin
      done_buf[1] <= done_buf[0];
    end else begin
      done_buf[1] <= 0;
    end
  end

  // Register the inputs
  always_ff @(posedge clk) begin
    if (reset) begin
      rtmp <= 0;
      ltmp <= 0;
    end else if (go) begin
      if (SIGNED) begin
        rtmp <= $signed(right);
        ltmp <= $signed(left);
      end else begin
        rtmp <= right;
        ltmp <= left;
      end
    end else begin
      rtmp <= 0;
      ltmp <= 0;
    end

  end

  // Compute the output and save it into out_tmp
  always_ff @(posedge clk) begin
    if (reset) begin
      out_tmp <= 0;
    end else if (go) begin
      if (SIGNED) begin
        // In the first cycle, this performs an invalid computation because
        // ltmp and rtmp only get their actual values in cycle 1
        out_tmp <= $signed(
          { {WIDTH{ltmp[WIDTH-1]}}, ltmp} *
          { {WIDTH{rtmp[WIDTH-1]}}, rtmp}
        );
      end else begin
        out_tmp <= ltmp * rtmp;
      end
    end else begin
      out_tmp <= out_tmp;
    end
  end
endmodule

/* verilator lint_off WIDTH */
module std_fp_div_pipe #(
  parameter WIDTH = 32,
  parameter INT_WIDTH = 16,
  parameter FRAC_WIDTH = 16
) (
    input  logic             go,
    input  logic             clk,
    input  logic             reset,
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out_remainder,
    output logic [WIDTH-1:0] out_quotient,
    output logic             done
);
    localparam ITERATIONS = WIDTH + FRAC_WIDTH;

    logic [WIDTH-1:0] quotient, quotient_next;
    logic [WIDTH:0] acc, acc_next;
    logic [$clog2(ITERATIONS)-1:0] idx;
    logic start, running, finished, dividend_is_zero;

    assign start = go && !running;
    assign dividend_is_zero = start && left == 0;
    assign finished = idx == ITERATIONS - 1 && running;

    always_ff @(posedge clk) begin
      if (reset || finished || dividend_is_zero)
        running <= 0;
      else if (start)
        running <= 1;
      else
        running <= running;
    end

    always_comb begin
      if (acc >= {1'b0, right}) begin
        acc_next = acc - right;
        {acc_next, quotient_next} = {acc_next[WIDTH-1:0], quotient, 1'b1};
      end else begin
        {acc_next, quotient_next} = {acc, quotient} << 1;
      end
    end

    // `done` signaling
    always_ff @(posedge clk) begin
      if (dividend_is_zero || finished)
        done <= 1;
      else
        done <= 0;
    end

    always_ff @(posedge clk) begin
      if (running)
        idx <= idx + 1;
      else
        idx <= 0;
    end

    always_ff @(posedge clk) begin
      if (reset) begin
        out_quotient <= 0;
        out_remainder <= 0;
      end else if (start) begin
        out_quotient <= 0;
        out_remainder <= left;
      end else if (go == 0) begin
        out_quotient <= out_quotient;
        out_remainder <= out_remainder;
      end else if (dividend_is_zero) begin
        out_quotient <= 0;
        out_remainder <= 0;
      end else if (finished) begin
        out_quotient <= quotient_next;
        out_remainder <= out_remainder;
      end else begin
        out_quotient <= out_quotient;
        if (right <= out_remainder)
          out_remainder <= out_remainder - right;
        else
          out_remainder <= out_remainder;
      end
    end

    always_ff @(posedge clk) begin
      if (reset) begin
        acc <= 0;
        quotient <= 0;
      end else if (start) begin
        {acc, quotient} <= {{WIDTH{1'b0}}, left, 1'b0};
      end else begin
        acc <= acc_next;
        quotient <= quotient_next;
      end
    end
endmodule

module std_fp_gt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic             out
);
  assign out = left > right;
endmodule

/// =================== Signed, Fixed Point =========================
module std_fp_sadd #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left + right);
endmodule

module std_fp_ssub #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);

  assign out = $signed(left - right);
endmodule

module std_fp_smult_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  [WIDTH-1:0]              left,
    input  [WIDTH-1:0]              right,
    input  logic                    reset,
    input  logic                    go,
    input  logic                    clk,
    output logic [WIDTH-1:0]        out,
    output logic                    done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(INT_WIDTH),
    .FRAC_WIDTH(FRAC_WIDTH),
    .SIGNED(1)
  ) comp (
    .clk(clk),
    .done(done),
    .reset(reset),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

module std_fp_sdiv_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input                     clk,
    input                     go,
    input                     reset,
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out_quotient,
    output signed [WIDTH-1:0] out_remainder,
    output logic              done
);

  logic signed [WIDTH-1:0] left_abs, right_abs, comp_out_q, comp_out_r, right_save, out_rem_intermediate;

  // Registers to figure out how to transform outputs.
  logic different_signs, left_sign, right_sign;

  // Latch the value of control registers so that their available after
  // go signal becomes low.
  always_ff @(posedge clk) begin
    if (go) begin
      right_save <= right_abs;
      left_sign <= left[WIDTH-1];
      right_sign <= right[WIDTH-1];
    end else begin
      left_sign <= left_sign;
      right_save <= right_save;
      right_sign <= right_sign;
    end
  end

  assign right_abs = right[WIDTH-1] ? -right : right;
  assign left_abs = left[WIDTH-1] ? -left : left;

  assign different_signs = left_sign ^ right_sign;
  assign out_quotient = different_signs ? -comp_out_q : comp_out_q;

  // Remainder is computed as:
  //  t0 = |left| % |right|
  //  t1 = if left * right < 0 and t0 != 0 then |right| - t0 else t0
  //  rem = if right < 0 then -t1 else t1
  assign out_rem_intermediate = different_signs & |comp_out_r ? $signed(right_save - comp_out_r) : comp_out_r;
  assign out_remainder = right_sign ? -out_rem_intermediate : out_rem_intermediate;

  std_fp_div_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(INT_WIDTH),
    .FRAC_WIDTH(FRAC_WIDTH)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left_abs),
    .right(right_abs),
    .out_quotient(comp_out_q),
    .out_remainder(comp_out_r)
  );
endmodule

module std_fp_sgt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic signed [WIDTH-1:0] left,
    input  logic signed [WIDTH-1:0] right,
    output logic signed             out
);
  assign out = $signed(left > right);
endmodule

module std_fp_slt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
   input logic signed [WIDTH-1:0] left,
   input logic signed [WIDTH-1:0] right,
   output logic signed            out
);
  assign out = $signed(left < right);
endmodule

/// =================== Unsigned, Bitnum =========================
module std_mult_pipe #(
    parameter WIDTH = 32
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    input  logic             reset,
    input  logic             go,
    input  logic             clk,
    output logic [WIDTH-1:0] out,
    output logic             done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(WIDTH),
    .FRAC_WIDTH(0),
    .SIGNED(0)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

module std_div_pipe #(
    parameter WIDTH = 32
) (
    input                    reset,
    input                    clk,
    input                    go,
    input        [WIDTH-1:0] left,
    input        [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out_remainder,
    output logic [WIDTH-1:0] out_quotient,
    output logic             done
);

  logic [WIDTH-1:0] dividend;
  logic [(WIDTH-1)*2:0] divisor;
  logic [WIDTH-1:0] quotient;
  logic [WIDTH-1:0] quotient_msk;
  logic start, running, finished, dividend_is_zero;

  assign start = go && !running;
  assign finished = quotient_msk == 0 && running;
  assign dividend_is_zero = start && left == 0;

  always_ff @(posedge clk) begin
    // Early return if the divisor is zero.
    if (finished || dividend_is_zero)
      done <= 1;
    else
      done <= 0;
  end

  always_ff @(posedge clk) begin
    if (reset || finished || dividend_is_zero)
      running <= 0;
    else if (start)
      running <= 1;
    else
      running <= running;
  end

  // Outputs
  always_ff @(posedge clk) begin
    if (dividend_is_zero || start) begin
      out_quotient <= 0;
      out_remainder <= 0;
    end else if (finished) begin
      out_quotient <= quotient;
      out_remainder <= dividend;
    end else begin
      // Otherwise, explicitly latch the values.
      out_quotient <= out_quotient;
      out_remainder <= out_remainder;
    end
  end

  // Calculate the quotient mask.
  always_ff @(posedge clk) begin
    if (start)
      quotient_msk <= 1 << WIDTH - 1;
    else if (running)
      quotient_msk <= quotient_msk >> 1;
    else
      quotient_msk <= quotient_msk;
  end

  // Calculate the quotient.
  always_ff @(posedge clk) begin
    if (start)
      quotient <= 0;
    else if (divisor <= dividend)
      quotient <= quotient | quotient_msk;
    else
      quotient <= quotient;
  end

  // Calculate the dividend.
  always_ff @(posedge clk) begin
    if (start)
      dividend <= left;
    else if (divisor <= dividend)
      dividend <= dividend - divisor;
    else
      dividend <= dividend;
  end

  always_ff @(posedge clk) begin
    if (start) begin
      divisor <= right << WIDTH - 1;
    end else if (finished) begin
      divisor <= 0;
    end else begin
      divisor <= divisor >> 1;
    end
  end

  // Simulation self test against unsynthesizable implementation.
  `ifdef VERILATOR
    logic [WIDTH-1:0] l, r;
    always_ff @(posedge clk) begin
      if (go) begin
        l <= left;
        r <= right;
      end else begin
        l <= l;
        r <= r;
      end
    end

    always @(posedge clk) begin
      if (done && $unsigned(out_remainder) != $unsigned(l % r))
        $error(
          "\nstd_div_pipe (Remainder): Computed and golden outputs do not match!\n",
          "left: %0d", $unsigned(l),
          "  right: %0d\n", $unsigned(r),
          "expected: %0d", $unsigned(l % r),
          "  computed: %0d", $unsigned(out_remainder)
        );

      if (done && $unsigned(out_quotient) != $unsigned(l / r))
        $error(
          "\nstd_div_pipe (Quotient): Computed and golden outputs do not match!\n",
          "left: %0d", $unsigned(l),
          "  right: %0d\n", $unsigned(r),
          "expected: %0d", $unsigned(l / r),
          "  computed: %0d", $unsigned(out_quotient)
        );
    end
  `endif
endmodule

/// =================== Signed, Bitnum =========================
module std_sadd #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left + right);
endmodule

module std_ssub #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left - right);
endmodule

module std_smult_pipe #(
    parameter WIDTH = 32
) (
    input  logic                    reset,
    input  logic                    go,
    input  logic                    clk,
    input  signed       [WIDTH-1:0] left,
    input  signed       [WIDTH-1:0] right,
    output logic signed [WIDTH-1:0] out,
    output logic                    done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(WIDTH),
    .FRAC_WIDTH(0),
    .SIGNED(1)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

/* verilator lint_off WIDTH */
module std_sdiv_pipe #(
    parameter WIDTH = 32
) (
    input                           reset,
    input                           clk,
    input                           go,
    input  logic signed [WIDTH-1:0] left,
    input  logic signed [WIDTH-1:0] right,
    output logic signed [WIDTH-1:0] out_quotient,
    output logic signed [WIDTH-1:0] out_remainder,
    output logic                    done
);

  logic signed [WIDTH-1:0] left_abs, right_abs, comp_out_q, comp_out_r, right_save, out_rem_intermediate;

  // Registers to figure out how to transform outputs.
  logic different_signs, left_sign, right_sign;

  // Latch the value of control registers so that their available after
  // go signal becomes low.
  always_ff @(posedge clk) begin
    if (go) begin
      right_save <= right_abs;
      left_sign <= left[WIDTH-1];
      right_sign <= right[WIDTH-1];
    end else begin
      left_sign <= left_sign;
      right_save <= right_save;
      right_sign <= right_sign;
    end
  end

  assign right_abs = right[WIDTH-1] ? -right : right;
  assign left_abs = left[WIDTH-1] ? -left : left;

  assign different_signs = left_sign ^ right_sign;
  assign out_quotient = different_signs ? -comp_out_q : comp_out_q;

  // Remainder is computed as:
  //  t0 = |left| % |right|
  //  t1 = if left * right < 0 and t0 != 0 then |right| - t0 else t0
  //  rem = if right < 0 then -t1 else t1
  assign out_rem_intermediate = different_signs & |comp_out_r ? $signed(right_save - comp_out_r) : comp_out_r;
  assign out_remainder = right_sign ? -out_rem_intermediate : out_rem_intermediate;

  std_div_pipe #(
    .WIDTH(WIDTH)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left_abs),
    .right(right_abs),
    .out_quotient(comp_out_q),
    .out_remainder(comp_out_r)
  );

  // Simulation self test against unsynthesizable implementation.
  `ifdef VERILATOR
    logic signed [WIDTH-1:0] l, r;
    always_ff @(posedge clk) begin
      if (go) begin
        l <= left;
        r <= right;
      end else begin
        l <= l;
        r <= r;
      end
    end

    always @(posedge clk) begin
      if (done && out_quotient != $signed(l / r))
        $error(
          "\nstd_sdiv_pipe (Quotient): Computed and golden outputs do not match!\n",
          "left: %0d", l,
          "  right: %0d\n", r,
          "expected: %0d", $signed(l / r),
          "  computed: %0d", $signed(out_quotient),
        );
      if (done && out_remainder != $signed(((l % r) + r) % r))
        $error(
          "\nstd_sdiv_pipe (Remainder): Computed and golden outputs do not match!\n",
          "left: %0d", l,
          "  right: %0d\n", r,
          "expected: %0d", $signed(((l % r) + r) % r),
          "  computed: %0d", $signed(out_remainder),
        );
    end
  `endif
endmodule

module std_sgt #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left > right);
endmodule

module std_slt #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left < right);
endmodule

module std_seq #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left == right);
endmodule

module std_sneq #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left != right);
endmodule

module std_sge #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left >= right);
endmodule

module std_sle #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left <= right);
endmodule

module std_slsh #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = left <<< right;
endmodule

module std_srsh #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = left >>> right;
endmodule

/**
 * Core primitives for Calyx.
 * Implements core primitives used by the compiler.
 *
 * Conventions:
 * - All parameter names must be SNAKE_CASE and all caps.
 * - Port names must be snake_case, no caps.
 */
`default_nettype none

module std_slice #(
    parameter IN_WIDTH  = 32,
    parameter OUT_WIDTH = 32
) (
   input wire                   logic [ IN_WIDTH-1:0] in,
   output logic [OUT_WIDTH-1:0] out
);
  assign out = in[OUT_WIDTH-1:0];

  `ifdef VERILATOR
    always_comb begin
      if (IN_WIDTH < OUT_WIDTH)
        $error(
          "std_slice: Input width less than output width\n",
          "IN_WIDTH: %0d", IN_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_pad #(
    parameter IN_WIDTH  = 32,
    parameter OUT_WIDTH = 32
) (
   input wire logic [IN_WIDTH-1:0]  in,
   output logic     [OUT_WIDTH-1:0] out
);
  localparam EXTEND = OUT_WIDTH - IN_WIDTH;
  assign out = { {EXTEND {1'b0}}, in};

  `ifdef VERILATOR
    always_comb begin
      if (IN_WIDTH > OUT_WIDTH)
        $error(
          "std_pad: Output width less than input width\n",
          "IN_WIDTH: %0d", IN_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_cat #(
  parameter LEFT_WIDTH  = 32,
  parameter RIGHT_WIDTH = 32,
  parameter OUT_WIDTH = 64
) (
  input wire logic [LEFT_WIDTH-1:0] left,
  input wire logic [RIGHT_WIDTH-1:0] right,
  output logic [OUT_WIDTH-1:0] out
);
  assign out = {left, right};

  `ifdef VERILATOR
    always_comb begin
      if (LEFT_WIDTH + RIGHT_WIDTH != OUT_WIDTH)
        $error(
          "std_cat: Output width must equal sum of input widths\n",
          "LEFT_WIDTH: %0d", LEFT_WIDTH,
          "RIGHT_WIDTH: %0d", RIGHT_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_not #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] in,
   output logic [WIDTH-1:0] out
);
  assign out = ~in;
endmodule

module std_and #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left & right;
endmodule

module std_or #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left | right;
endmodule

module std_xor #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left ^ right;
endmodule

module std_sub #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module std_gt #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left > right;
endmodule

module std_lt #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left < right;
endmodule

module std_eq #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left == right;
endmodule

module std_neq #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left != right;
endmodule

module std_ge #(
    parameter WIDTH = 32
) (
    input wire   logic [WIDTH-1:0] left,
    input wire   logic [WIDTH-1:0] right,
    output logic out
);
  assign out = left >= right;
endmodule

module std_le #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left <= right;
endmodule

module std_lsh #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left << right;
endmodule

module std_rsh #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left >> right;
endmodule

/// this primitive is intended to be used
/// for lowering purposes (not in source programs)
module std_mux #(
    parameter WIDTH = 32
) (
   input wire               logic cond,
   input wire               logic [WIDTH-1:0] tru,
   input wire               logic [WIDTH-1:0] fal,
   output logic [WIDTH-1:0] out
);
  assign out = cond ? tru : fal;
endmodule

module std_mem_d1 #(
    parameter WIDTH = 32,
    parameter SIZE = 16,
    parameter IDX_SIZE = 4
) (
   input wire                logic [IDX_SIZE-1:0] addr0,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  logic [WIDTH-1:0] mem[SIZE-1:0];

  /* verilator lint_off WIDTH */
  assign read_data = mem[addr0];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= SIZE)
        $error(
          "std_mem_d1: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "SIZE: %0d", SIZE
        );
    end
  `endif
endmodule

module std_mem_d2 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0];

  assign read_data = mem[addr0][addr1];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d2: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d2: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
    end
  `endif
endmodule

module std_mem_d3 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D2_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4,
    parameter D2_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [D2_IDX_SIZE-1:0] addr2,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0][D2_SIZE-1:0];

  assign read_data = mem[addr0][addr1][addr2];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1][addr2] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
      if (addr2 >= D2_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr2: %0d\n", addr2,
          "D2_SIZE: %0d", D2_SIZE
        );
    end
  `endif
endmodule

module std_mem_d4 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D2_SIZE = 16,
    parameter D3_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4,
    parameter D2_IDX_SIZE = 4,
    parameter D3_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [D2_IDX_SIZE-1:0] addr2,
   input wire                logic [D3_IDX_SIZE-1:0] addr3,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0][D2_SIZE-1:0][D3_SIZE-1:0];

  assign read_data = mem[addr0][addr1][addr2][addr3];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1][addr2][addr3] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
      if (addr2 >= D2_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr2: %0d\n", addr2,
          "D2_SIZE: %0d", D2_SIZE
        );
      if (addr3 >= D3_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr3: %0d\n", addr3,
          "D3_SIZE: %0d", D3_SIZE
        );
    end
  `endif
endmodule

`default_nettype wire

module undef #(
    parameter WIDTH = 32
) (
   output logic [WIDTH-1:0] out
);
assign out = 'x;
endmodule

module std_const #(
    parameter WIDTH = 32,
    parameter VALUE = 32
) (
   output logic [WIDTH-1:0] out
);
assign out = VALUE;
endmodule

module std_wire #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] in,
   output logic [WIDTH-1:0] out
);
assign out = in;
endmodule

module std_add #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] left,
   input logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
assign out = left + right;
endmodule

module std_reg #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] in,
   input logic write_en,
   input logic clk,
   input logic reset,
   output logic [WIDTH-1:0] out,
   output logic done
);
always_ff @(posedge clk) begin
    if (reset) begin
       out <= 0;
       done <= 0;
    end else if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module mac_pe(
  input logic [31:0] top,
  input logic [31:0] left,
  input logic mul_ready,
  output logic [31:0] out,
  input logic go,
  input logic clk,
  input logic reset,
  output logic done
);
// COMPONENT START: mac_pe
logic [31:0] acc_in;
logic acc_write_en;
logic acc_clk;
logic acc_reset;
logic [31:0] acc_out;
logic acc_done;
logic [31:0] add_left;
logic [31:0] add_right;
logic [31:0] add_out;
logic mul_clk;
logic [31:0] mul_left;
logic [31:0] mul_right;
logic [31:0] mul_out;
logic fsm_in;
logic fsm_write_en;
logic fsm_clk;
logic fsm_reset;
logic fsm_out;
logic fsm_done;
logic ud_out;
logic adder_left;
logic adder_right;
logic adder_out;
logic signal_reg_in;
logic signal_reg_write_en;
logic signal_reg_clk;
logic signal_reg_reset;
logic signal_reg_out;
logic signal_reg_done;
logic early_reset_static_par_go_in;
logic early_reset_static_par_go_out;
logic early_reset_static_par_done_in;
logic early_reset_static_par_done_out;
logic wrapper_early_reset_static_par_go_in;
logic wrapper_early_reset_static_par_go_out;
logic wrapper_early_reset_static_par_done_in;
logic wrapper_early_reset_static_par_done_out;
std_reg # (
    .WIDTH(32)
) acc (
    .clk(acc_clk),
    .done(acc_done),
    .in(acc_in),
    .out(acc_out),
    .reset(acc_reset),
    .write_en(acc_write_en)
);
std_add # (
    .WIDTH(32)
) add (
    .left(add_left),
    .out(add_out),
    .right(add_right)
);
bb_pipelined_mult mul (
    .clk(mul_clk),
    .left(mul_left),
    .out(mul_out),
    .right(mul_right)
);
std_reg # (
    .WIDTH(1)
) fsm (
    .clk(fsm_clk),
    .done(fsm_done),
    .in(fsm_in),
    .out(fsm_out),
    .reset(fsm_reset),
    .write_en(fsm_write_en)
);
undef # (
    .WIDTH(1)
) ud (
    .out(ud_out)
);
std_add # (
    .WIDTH(1)
) adder (
    .left(adder_left),
    .out(adder_out),
    .right(adder_right)
);
std_reg # (
    .WIDTH(1)
) signal_reg (
    .clk(signal_reg_clk),
    .done(signal_reg_done),
    .in(signal_reg_in),
    .out(signal_reg_out),
    .reset(signal_reg_reset),
    .write_en(signal_reg_write_en)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_go (
    .in(early_reset_static_par_go_in),
    .out(early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_done (
    .in(early_reset_static_par_done_in),
    .out(early_reset_static_par_done_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_go (
    .in(wrapper_early_reset_static_par_go_in),
    .out(wrapper_early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_done (
    .in(wrapper_early_reset_static_par_done_in),
    .out(wrapper_early_reset_static_par_done_out)
);
wire _guard0 = 1;
wire _guard1 = early_reset_static_par_go_out;
wire _guard2 = early_reset_static_par_go_out;
wire _guard3 = wrapper_early_reset_static_par_done_out;
wire _guard4 = early_reset_static_par_go_out;
wire _guard5 = fsm_out != 1'd0;
wire _guard6 = early_reset_static_par_go_out;
wire _guard7 = _guard5 & _guard6;
wire _guard8 = fsm_out == 1'd0;
wire _guard9 = early_reset_static_par_go_out;
wire _guard10 = _guard8 & _guard9;
wire _guard11 = early_reset_static_par_go_out;
wire _guard12 = early_reset_static_par_go_out;
wire _guard13 = fsm_out == 1'd0;
wire _guard14 = signal_reg_out;
wire _guard15 = _guard13 & _guard14;
wire _guard16 = fsm_out == 1'd0;
wire _guard17 = signal_reg_out;
wire _guard18 = _guard16 & _guard17;
wire _guard19 = fsm_out == 1'd0;
wire _guard20 = signal_reg_out;
wire _guard21 = ~_guard20;
wire _guard22 = _guard19 & _guard21;
wire _guard23 = wrapper_early_reset_static_par_go_out;
wire _guard24 = _guard22 & _guard23;
wire _guard25 = _guard18 | _guard24;
wire _guard26 = fsm_out == 1'd0;
wire _guard27 = signal_reg_out;
wire _guard28 = ~_guard27;
wire _guard29 = _guard26 & _guard28;
wire _guard30 = wrapper_early_reset_static_par_go_out;
wire _guard31 = _guard29 & _guard30;
wire _guard32 = fsm_out == 1'd0;
wire _guard33 = signal_reg_out;
wire _guard34 = _guard32 & _guard33;
wire _guard35 = early_reset_static_par_go_out;
wire _guard36 = early_reset_static_par_go_out;
wire _guard37 = early_reset_static_par_go_out;
wire _guard38 = early_reset_static_par_go_out;
wire _guard39 = wrapper_early_reset_static_par_go_out;
assign acc_write_en =
  _guard1 ? mul_ready :
  1'd0;
assign acc_clk = clk;
assign acc_reset = reset;
assign acc_in = add_out;
assign done = _guard3;
assign out = acc_out;
assign fsm_write_en = _guard4;
assign fsm_clk = clk;
assign fsm_reset = reset;
assign fsm_in =
  _guard7 ? adder_out :
  _guard10 ? 1'd0 :
  1'd0;
assign adder_left =
  _guard11 ? fsm_out :
  1'd0;
assign adder_right = _guard12;
assign wrapper_early_reset_static_par_go_in = go;
assign wrapper_early_reset_static_par_done_in = _guard15;
assign early_reset_static_par_done_in = ud_out;
assign signal_reg_write_en = _guard25;
assign signal_reg_clk = clk;
assign signal_reg_reset = reset;
assign signal_reg_in =
  _guard31 ? 1'd1 :
  _guard34 ? 1'd0 :
  1'd0;
assign add_left = acc_out;
assign add_right = mul_out;
assign mul_clk = clk;
assign mul_left =
  _guard37 ? top :
  32'd0;
assign mul_right =
  _guard38 ? left :
  32'd0;
assign early_reset_static_par_go_in = _guard39;
// COMPONENT END: mac_pe
endmodule
module main(
  input logic go,
  input logic clk,
  input logic reset,
  output logic done,
  output logic [3:0] t0_addr0,
  output logic [31:0] t0_write_data,
  output logic t0_write_en,
  output logic t0_clk,
  output logic t0_reset,
  input logic [31:0] t0_read_data,
  input logic t0_done,
  output logic [3:0] t1_addr0,
  output logic [31:0] t1_write_data,
  output logic t1_write_en,
  output logic t1_clk,
  output logic t1_reset,
  input logic [31:0] t1_read_data,
  input logic t1_done,
  output logic [3:0] t2_addr0,
  output logic [31:0] t2_write_data,
  output logic t2_write_en,
  output logic t2_clk,
  output logic t2_reset,
  input logic [31:0] t2_read_data,
  input logic t2_done,
  output logic [3:0] t3_addr0,
  output logic [31:0] t3_write_data,
  output logic t3_write_en,
  output logic t3_clk,
  output logic t3_reset,
  input logic [31:0] t3_read_data,
  input logic t3_done,
  output logic [3:0] t4_addr0,
  output logic [31:0] t4_write_data,
  output logic t4_write_en,
  output logic t4_clk,
  output logic t4_reset,
  input logic [31:0] t4_read_data,
  input logic t4_done,
  output logic [3:0] t5_addr0,
  output logic [31:0] t5_write_data,
  output logic t5_write_en,
  output logic t5_clk,
  output logic t5_reset,
  input logic [31:0] t5_read_data,
  input logic t5_done,
  output logic [3:0] t6_addr0,
  output logic [31:0] t6_write_data,
  output logic t6_write_en,
  output logic t6_clk,
  output logic t6_reset,
  input logic [31:0] t6_read_data,
  input logic t6_done,
  output logic [3:0] t7_addr0,
  output logic [31:0] t7_write_data,
  output logic t7_write_en,
  output logic t7_clk,
  output logic t7_reset,
  input logic [31:0] t7_read_data,
  input logic t7_done,
  output logic [3:0] l0_addr0,
  output logic [31:0] l0_write_data,
  output logic l0_write_en,
  output logic l0_clk,
  output logic l0_reset,
  input logic [31:0] l0_read_data,
  input logic l0_done,
  output logic [3:0] l1_addr0,
  output logic [31:0] l1_write_data,
  output logic l1_write_en,
  output logic l1_clk,
  output logic l1_reset,
  input logic [31:0] l1_read_data,
  input logic l1_done,
  output logic [3:0] l2_addr0,
  output logic [31:0] l2_write_data,
  output logic l2_write_en,
  output logic l2_clk,
  output logic l2_reset,
  input logic [31:0] l2_read_data,
  input logic l2_done,
  output logic [3:0] l3_addr0,
  output logic [31:0] l3_write_data,
  output logic l3_write_en,
  output logic l3_clk,
  output logic l3_reset,
  input logic [31:0] l3_read_data,
  input logic l3_done,
  output logic [3:0] l4_addr0,
  output logic [31:0] l4_write_data,
  output logic l4_write_en,
  output logic l4_clk,
  output logic l4_reset,
  input logic [31:0] l4_read_data,
  input logic l4_done,
  output logic [3:0] l5_addr0,
  output logic [31:0] l5_write_data,
  output logic l5_write_en,
  output logic l5_clk,
  output logic l5_reset,
  input logic [31:0] l5_read_data,
  input logic l5_done,
  output logic [3:0] l6_addr0,
  output logic [31:0] l6_write_data,
  output logic l6_write_en,
  output logic l6_clk,
  output logic l6_reset,
  input logic [31:0] l6_read_data,
  input logic l6_done,
  output logic [3:0] l7_addr0,
  output logic [31:0] l7_write_data,
  output logic l7_write_en,
  output logic l7_clk,
  output logic l7_reset,
  input logic [31:0] l7_read_data,
  input logic l7_done,
  output logic [3:0] out_mem_0_addr0,
  output logic [31:0] out_mem_0_write_data,
  output logic out_mem_0_write_en,
  output logic out_mem_0_clk,
  output logic out_mem_0_reset,
  input logic [31:0] out_mem_0_read_data,
  input logic out_mem_0_done,
  output logic [3:0] out_mem_1_addr0,
  output logic [31:0] out_mem_1_write_data,
  output logic out_mem_1_write_en,
  output logic out_mem_1_clk,
  output logic out_mem_1_reset,
  input logic [31:0] out_mem_1_read_data,
  input logic out_mem_1_done,
  output logic [3:0] out_mem_2_addr0,
  output logic [31:0] out_mem_2_write_data,
  output logic out_mem_2_write_en,
  output logic out_mem_2_clk,
  output logic out_mem_2_reset,
  input logic [31:0] out_mem_2_read_data,
  input logic out_mem_2_done,
  output logic [3:0] out_mem_3_addr0,
  output logic [31:0] out_mem_3_write_data,
  output logic out_mem_3_write_en,
  output logic out_mem_3_clk,
  output logic out_mem_3_reset,
  input logic [31:0] out_mem_3_read_data,
  input logic out_mem_3_done,
  output logic [3:0] out_mem_4_addr0,
  output logic [31:0] out_mem_4_write_data,
  output logic out_mem_4_write_en,
  output logic out_mem_4_clk,
  output logic out_mem_4_reset,
  input logic [31:0] out_mem_4_read_data,
  input logic out_mem_4_done,
  output logic [3:0] out_mem_5_addr0,
  output logic [31:0] out_mem_5_write_data,
  output logic out_mem_5_write_en,
  output logic out_mem_5_clk,
  output logic out_mem_5_reset,
  input logic [31:0] out_mem_5_read_data,
  input logic out_mem_5_done,
  output logic [3:0] out_mem_6_addr0,
  output logic [31:0] out_mem_6_write_data,
  output logic out_mem_6_write_en,
  output logic out_mem_6_clk,
  output logic out_mem_6_reset,
  input logic [31:0] out_mem_6_read_data,
  input logic out_mem_6_done,
  output logic [3:0] out_mem_7_addr0,
  output logic [31:0] out_mem_7_write_data,
  output logic out_mem_7_write_en,
  output logic out_mem_7_clk,
  output logic out_mem_7_reset,
  input logic [31:0] out_mem_7_read_data,
  input logic out_mem_7_done
);
// COMPONENT START: main
logic [31:0] pe_0_0_top;
logic [31:0] pe_0_0_left;
logic pe_0_0_mul_ready;
logic [31:0] pe_0_0_out;
logic pe_0_0_go;
logic pe_0_0_clk;
logic pe_0_0_reset;
logic pe_0_0_done;
logic [31:0] top_0_0_in;
logic top_0_0_write_en;
logic top_0_0_clk;
logic top_0_0_reset;
logic [31:0] top_0_0_out;
logic top_0_0_done;
logic [31:0] left_0_0_in;
logic left_0_0_write_en;
logic left_0_0_clk;
logic left_0_0_reset;
logic [31:0] left_0_0_out;
logic left_0_0_done;
logic [31:0] pe_0_1_top;
logic [31:0] pe_0_1_left;
logic pe_0_1_mul_ready;
logic [31:0] pe_0_1_out;
logic pe_0_1_go;
logic pe_0_1_clk;
logic pe_0_1_reset;
logic pe_0_1_done;
logic [31:0] top_0_1_in;
logic top_0_1_write_en;
logic top_0_1_clk;
logic top_0_1_reset;
logic [31:0] top_0_1_out;
logic top_0_1_done;
logic [31:0] left_0_1_in;
logic left_0_1_write_en;
logic left_0_1_clk;
logic left_0_1_reset;
logic [31:0] left_0_1_out;
logic left_0_1_done;
logic [31:0] pe_0_2_top;
logic [31:0] pe_0_2_left;
logic pe_0_2_mul_ready;
logic [31:0] pe_0_2_out;
logic pe_0_2_go;
logic pe_0_2_clk;
logic pe_0_2_reset;
logic pe_0_2_done;
logic [31:0] top_0_2_in;
logic top_0_2_write_en;
logic top_0_2_clk;
logic top_0_2_reset;
logic [31:0] top_0_2_out;
logic top_0_2_done;
logic [31:0] left_0_2_in;
logic left_0_2_write_en;
logic left_0_2_clk;
logic left_0_2_reset;
logic [31:0] left_0_2_out;
logic left_0_2_done;
logic [31:0] pe_0_3_top;
logic [31:0] pe_0_3_left;
logic pe_0_3_mul_ready;
logic [31:0] pe_0_3_out;
logic pe_0_3_go;
logic pe_0_3_clk;
logic pe_0_3_reset;
logic pe_0_3_done;
logic [31:0] top_0_3_in;
logic top_0_3_write_en;
logic top_0_3_clk;
logic top_0_3_reset;
logic [31:0] top_0_3_out;
logic top_0_3_done;
logic [31:0] left_0_3_in;
logic left_0_3_write_en;
logic left_0_3_clk;
logic left_0_3_reset;
logic [31:0] left_0_3_out;
logic left_0_3_done;
logic [31:0] pe_0_4_top;
logic [31:0] pe_0_4_left;
logic pe_0_4_mul_ready;
logic [31:0] pe_0_4_out;
logic pe_0_4_go;
logic pe_0_4_clk;
logic pe_0_4_reset;
logic pe_0_4_done;
logic [31:0] top_0_4_in;
logic top_0_4_write_en;
logic top_0_4_clk;
logic top_0_4_reset;
logic [31:0] top_0_4_out;
logic top_0_4_done;
logic [31:0] left_0_4_in;
logic left_0_4_write_en;
logic left_0_4_clk;
logic left_0_4_reset;
logic [31:0] left_0_4_out;
logic left_0_4_done;
logic [31:0] pe_0_5_top;
logic [31:0] pe_0_5_left;
logic pe_0_5_mul_ready;
logic [31:0] pe_0_5_out;
logic pe_0_5_go;
logic pe_0_5_clk;
logic pe_0_5_reset;
logic pe_0_5_done;
logic [31:0] top_0_5_in;
logic top_0_5_write_en;
logic top_0_5_clk;
logic top_0_5_reset;
logic [31:0] top_0_5_out;
logic top_0_5_done;
logic [31:0] left_0_5_in;
logic left_0_5_write_en;
logic left_0_5_clk;
logic left_0_5_reset;
logic [31:0] left_0_5_out;
logic left_0_5_done;
logic [31:0] pe_0_6_top;
logic [31:0] pe_0_6_left;
logic pe_0_6_mul_ready;
logic [31:0] pe_0_6_out;
logic pe_0_6_go;
logic pe_0_6_clk;
logic pe_0_6_reset;
logic pe_0_6_done;
logic [31:0] top_0_6_in;
logic top_0_6_write_en;
logic top_0_6_clk;
logic top_0_6_reset;
logic [31:0] top_0_6_out;
logic top_0_6_done;
logic [31:0] left_0_6_in;
logic left_0_6_write_en;
logic left_0_6_clk;
logic left_0_6_reset;
logic [31:0] left_0_6_out;
logic left_0_6_done;
logic [31:0] pe_0_7_top;
logic [31:0] pe_0_7_left;
logic pe_0_7_mul_ready;
logic [31:0] pe_0_7_out;
logic pe_0_7_go;
logic pe_0_7_clk;
logic pe_0_7_reset;
logic pe_0_7_done;
logic [31:0] top_0_7_in;
logic top_0_7_write_en;
logic top_0_7_clk;
logic top_0_7_reset;
logic [31:0] top_0_7_out;
logic top_0_7_done;
logic [31:0] left_0_7_in;
logic left_0_7_write_en;
logic left_0_7_clk;
logic left_0_7_reset;
logic [31:0] left_0_7_out;
logic left_0_7_done;
logic [31:0] pe_1_0_top;
logic [31:0] pe_1_0_left;
logic pe_1_0_mul_ready;
logic [31:0] pe_1_0_out;
logic pe_1_0_go;
logic pe_1_0_clk;
logic pe_1_0_reset;
logic pe_1_0_done;
logic [31:0] top_1_0_in;
logic top_1_0_write_en;
logic top_1_0_clk;
logic top_1_0_reset;
logic [31:0] top_1_0_out;
logic top_1_0_done;
logic [31:0] left_1_0_in;
logic left_1_0_write_en;
logic left_1_0_clk;
logic left_1_0_reset;
logic [31:0] left_1_0_out;
logic left_1_0_done;
logic [31:0] pe_1_1_top;
logic [31:0] pe_1_1_left;
logic pe_1_1_mul_ready;
logic [31:0] pe_1_1_out;
logic pe_1_1_go;
logic pe_1_1_clk;
logic pe_1_1_reset;
logic pe_1_1_done;
logic [31:0] top_1_1_in;
logic top_1_1_write_en;
logic top_1_1_clk;
logic top_1_1_reset;
logic [31:0] top_1_1_out;
logic top_1_1_done;
logic [31:0] left_1_1_in;
logic left_1_1_write_en;
logic left_1_1_clk;
logic left_1_1_reset;
logic [31:0] left_1_1_out;
logic left_1_1_done;
logic [31:0] pe_1_2_top;
logic [31:0] pe_1_2_left;
logic pe_1_2_mul_ready;
logic [31:0] pe_1_2_out;
logic pe_1_2_go;
logic pe_1_2_clk;
logic pe_1_2_reset;
logic pe_1_2_done;
logic [31:0] top_1_2_in;
logic top_1_2_write_en;
logic top_1_2_clk;
logic top_1_2_reset;
logic [31:0] top_1_2_out;
logic top_1_2_done;
logic [31:0] left_1_2_in;
logic left_1_2_write_en;
logic left_1_2_clk;
logic left_1_2_reset;
logic [31:0] left_1_2_out;
logic left_1_2_done;
logic [31:0] pe_1_3_top;
logic [31:0] pe_1_3_left;
logic pe_1_3_mul_ready;
logic [31:0] pe_1_3_out;
logic pe_1_3_go;
logic pe_1_3_clk;
logic pe_1_3_reset;
logic pe_1_3_done;
logic [31:0] top_1_3_in;
logic top_1_3_write_en;
logic top_1_3_clk;
logic top_1_3_reset;
logic [31:0] top_1_3_out;
logic top_1_3_done;
logic [31:0] left_1_3_in;
logic left_1_3_write_en;
logic left_1_3_clk;
logic left_1_3_reset;
logic [31:0] left_1_3_out;
logic left_1_3_done;
logic [31:0] pe_1_4_top;
logic [31:0] pe_1_4_left;
logic pe_1_4_mul_ready;
logic [31:0] pe_1_4_out;
logic pe_1_4_go;
logic pe_1_4_clk;
logic pe_1_4_reset;
logic pe_1_4_done;
logic [31:0] top_1_4_in;
logic top_1_4_write_en;
logic top_1_4_clk;
logic top_1_4_reset;
logic [31:0] top_1_4_out;
logic top_1_4_done;
logic [31:0] left_1_4_in;
logic left_1_4_write_en;
logic left_1_4_clk;
logic left_1_4_reset;
logic [31:0] left_1_4_out;
logic left_1_4_done;
logic [31:0] pe_1_5_top;
logic [31:0] pe_1_5_left;
logic pe_1_5_mul_ready;
logic [31:0] pe_1_5_out;
logic pe_1_5_go;
logic pe_1_5_clk;
logic pe_1_5_reset;
logic pe_1_5_done;
logic [31:0] top_1_5_in;
logic top_1_5_write_en;
logic top_1_5_clk;
logic top_1_5_reset;
logic [31:0] top_1_5_out;
logic top_1_5_done;
logic [31:0] left_1_5_in;
logic left_1_5_write_en;
logic left_1_5_clk;
logic left_1_5_reset;
logic [31:0] left_1_5_out;
logic left_1_5_done;
logic [31:0] pe_1_6_top;
logic [31:0] pe_1_6_left;
logic pe_1_6_mul_ready;
logic [31:0] pe_1_6_out;
logic pe_1_6_go;
logic pe_1_6_clk;
logic pe_1_6_reset;
logic pe_1_6_done;
logic [31:0] top_1_6_in;
logic top_1_6_write_en;
logic top_1_6_clk;
logic top_1_6_reset;
logic [31:0] top_1_6_out;
logic top_1_6_done;
logic [31:0] left_1_6_in;
logic left_1_6_write_en;
logic left_1_6_clk;
logic left_1_6_reset;
logic [31:0] left_1_6_out;
logic left_1_6_done;
logic [31:0] pe_1_7_top;
logic [31:0] pe_1_7_left;
logic pe_1_7_mul_ready;
logic [31:0] pe_1_7_out;
logic pe_1_7_go;
logic pe_1_7_clk;
logic pe_1_7_reset;
logic pe_1_7_done;
logic [31:0] top_1_7_in;
logic top_1_7_write_en;
logic top_1_7_clk;
logic top_1_7_reset;
logic [31:0] top_1_7_out;
logic top_1_7_done;
logic [31:0] left_1_7_in;
logic left_1_7_write_en;
logic left_1_7_clk;
logic left_1_7_reset;
logic [31:0] left_1_7_out;
logic left_1_7_done;
logic [31:0] pe_2_0_top;
logic [31:0] pe_2_0_left;
logic pe_2_0_mul_ready;
logic [31:0] pe_2_0_out;
logic pe_2_0_go;
logic pe_2_0_clk;
logic pe_2_0_reset;
logic pe_2_0_done;
logic [31:0] top_2_0_in;
logic top_2_0_write_en;
logic top_2_0_clk;
logic top_2_0_reset;
logic [31:0] top_2_0_out;
logic top_2_0_done;
logic [31:0] left_2_0_in;
logic left_2_0_write_en;
logic left_2_0_clk;
logic left_2_0_reset;
logic [31:0] left_2_0_out;
logic left_2_0_done;
logic [31:0] pe_2_1_top;
logic [31:0] pe_2_1_left;
logic pe_2_1_mul_ready;
logic [31:0] pe_2_1_out;
logic pe_2_1_go;
logic pe_2_1_clk;
logic pe_2_1_reset;
logic pe_2_1_done;
logic [31:0] top_2_1_in;
logic top_2_1_write_en;
logic top_2_1_clk;
logic top_2_1_reset;
logic [31:0] top_2_1_out;
logic top_2_1_done;
logic [31:0] left_2_1_in;
logic left_2_1_write_en;
logic left_2_1_clk;
logic left_2_1_reset;
logic [31:0] left_2_1_out;
logic left_2_1_done;
logic [31:0] pe_2_2_top;
logic [31:0] pe_2_2_left;
logic pe_2_2_mul_ready;
logic [31:0] pe_2_2_out;
logic pe_2_2_go;
logic pe_2_2_clk;
logic pe_2_2_reset;
logic pe_2_2_done;
logic [31:0] top_2_2_in;
logic top_2_2_write_en;
logic top_2_2_clk;
logic top_2_2_reset;
logic [31:0] top_2_2_out;
logic top_2_2_done;
logic [31:0] left_2_2_in;
logic left_2_2_write_en;
logic left_2_2_clk;
logic left_2_2_reset;
logic [31:0] left_2_2_out;
logic left_2_2_done;
logic [31:0] pe_2_3_top;
logic [31:0] pe_2_3_left;
logic pe_2_3_mul_ready;
logic [31:0] pe_2_3_out;
logic pe_2_3_go;
logic pe_2_3_clk;
logic pe_2_3_reset;
logic pe_2_3_done;
logic [31:0] top_2_3_in;
logic top_2_3_write_en;
logic top_2_3_clk;
logic top_2_3_reset;
logic [31:0] top_2_3_out;
logic top_2_3_done;
logic [31:0] left_2_3_in;
logic left_2_3_write_en;
logic left_2_3_clk;
logic left_2_3_reset;
logic [31:0] left_2_3_out;
logic left_2_3_done;
logic [31:0] pe_2_4_top;
logic [31:0] pe_2_4_left;
logic pe_2_4_mul_ready;
logic [31:0] pe_2_4_out;
logic pe_2_4_go;
logic pe_2_4_clk;
logic pe_2_4_reset;
logic pe_2_4_done;
logic [31:0] top_2_4_in;
logic top_2_4_write_en;
logic top_2_4_clk;
logic top_2_4_reset;
logic [31:0] top_2_4_out;
logic top_2_4_done;
logic [31:0] left_2_4_in;
logic left_2_4_write_en;
logic left_2_4_clk;
logic left_2_4_reset;
logic [31:0] left_2_4_out;
logic left_2_4_done;
logic [31:0] pe_2_5_top;
logic [31:0] pe_2_5_left;
logic pe_2_5_mul_ready;
logic [31:0] pe_2_5_out;
logic pe_2_5_go;
logic pe_2_5_clk;
logic pe_2_5_reset;
logic pe_2_5_done;
logic [31:0] top_2_5_in;
logic top_2_5_write_en;
logic top_2_5_clk;
logic top_2_5_reset;
logic [31:0] top_2_5_out;
logic top_2_5_done;
logic [31:0] left_2_5_in;
logic left_2_5_write_en;
logic left_2_5_clk;
logic left_2_5_reset;
logic [31:0] left_2_5_out;
logic left_2_5_done;
logic [31:0] pe_2_6_top;
logic [31:0] pe_2_6_left;
logic pe_2_6_mul_ready;
logic [31:0] pe_2_6_out;
logic pe_2_6_go;
logic pe_2_6_clk;
logic pe_2_6_reset;
logic pe_2_6_done;
logic [31:0] top_2_6_in;
logic top_2_6_write_en;
logic top_2_6_clk;
logic top_2_6_reset;
logic [31:0] top_2_6_out;
logic top_2_6_done;
logic [31:0] left_2_6_in;
logic left_2_6_write_en;
logic left_2_6_clk;
logic left_2_6_reset;
logic [31:0] left_2_6_out;
logic left_2_6_done;
logic [31:0] pe_2_7_top;
logic [31:0] pe_2_7_left;
logic pe_2_7_mul_ready;
logic [31:0] pe_2_7_out;
logic pe_2_7_go;
logic pe_2_7_clk;
logic pe_2_7_reset;
logic pe_2_7_done;
logic [31:0] top_2_7_in;
logic top_2_7_write_en;
logic top_2_7_clk;
logic top_2_7_reset;
logic [31:0] top_2_7_out;
logic top_2_7_done;
logic [31:0] left_2_7_in;
logic left_2_7_write_en;
logic left_2_7_clk;
logic left_2_7_reset;
logic [31:0] left_2_7_out;
logic left_2_7_done;
logic [31:0] pe_3_0_top;
logic [31:0] pe_3_0_left;
logic pe_3_0_mul_ready;
logic [31:0] pe_3_0_out;
logic pe_3_0_go;
logic pe_3_0_clk;
logic pe_3_0_reset;
logic pe_3_0_done;
logic [31:0] top_3_0_in;
logic top_3_0_write_en;
logic top_3_0_clk;
logic top_3_0_reset;
logic [31:0] top_3_0_out;
logic top_3_0_done;
logic [31:0] left_3_0_in;
logic left_3_0_write_en;
logic left_3_0_clk;
logic left_3_0_reset;
logic [31:0] left_3_0_out;
logic left_3_0_done;
logic [31:0] pe_3_1_top;
logic [31:0] pe_3_1_left;
logic pe_3_1_mul_ready;
logic [31:0] pe_3_1_out;
logic pe_3_1_go;
logic pe_3_1_clk;
logic pe_3_1_reset;
logic pe_3_1_done;
logic [31:0] top_3_1_in;
logic top_3_1_write_en;
logic top_3_1_clk;
logic top_3_1_reset;
logic [31:0] top_3_1_out;
logic top_3_1_done;
logic [31:0] left_3_1_in;
logic left_3_1_write_en;
logic left_3_1_clk;
logic left_3_1_reset;
logic [31:0] left_3_1_out;
logic left_3_1_done;
logic [31:0] pe_3_2_top;
logic [31:0] pe_3_2_left;
logic pe_3_2_mul_ready;
logic [31:0] pe_3_2_out;
logic pe_3_2_go;
logic pe_3_2_clk;
logic pe_3_2_reset;
logic pe_3_2_done;
logic [31:0] top_3_2_in;
logic top_3_2_write_en;
logic top_3_2_clk;
logic top_3_2_reset;
logic [31:0] top_3_2_out;
logic top_3_2_done;
logic [31:0] left_3_2_in;
logic left_3_2_write_en;
logic left_3_2_clk;
logic left_3_2_reset;
logic [31:0] left_3_2_out;
logic left_3_2_done;
logic [31:0] pe_3_3_top;
logic [31:0] pe_3_3_left;
logic pe_3_3_mul_ready;
logic [31:0] pe_3_3_out;
logic pe_3_3_go;
logic pe_3_3_clk;
logic pe_3_3_reset;
logic pe_3_3_done;
logic [31:0] top_3_3_in;
logic top_3_3_write_en;
logic top_3_3_clk;
logic top_3_3_reset;
logic [31:0] top_3_3_out;
logic top_3_3_done;
logic [31:0] left_3_3_in;
logic left_3_3_write_en;
logic left_3_3_clk;
logic left_3_3_reset;
logic [31:0] left_3_3_out;
logic left_3_3_done;
logic [31:0] pe_3_4_top;
logic [31:0] pe_3_4_left;
logic pe_3_4_mul_ready;
logic [31:0] pe_3_4_out;
logic pe_3_4_go;
logic pe_3_4_clk;
logic pe_3_4_reset;
logic pe_3_4_done;
logic [31:0] top_3_4_in;
logic top_3_4_write_en;
logic top_3_4_clk;
logic top_3_4_reset;
logic [31:0] top_3_4_out;
logic top_3_4_done;
logic [31:0] left_3_4_in;
logic left_3_4_write_en;
logic left_3_4_clk;
logic left_3_4_reset;
logic [31:0] left_3_4_out;
logic left_3_4_done;
logic [31:0] pe_3_5_top;
logic [31:0] pe_3_5_left;
logic pe_3_5_mul_ready;
logic [31:0] pe_3_5_out;
logic pe_3_5_go;
logic pe_3_5_clk;
logic pe_3_5_reset;
logic pe_3_5_done;
logic [31:0] top_3_5_in;
logic top_3_5_write_en;
logic top_3_5_clk;
logic top_3_5_reset;
logic [31:0] top_3_5_out;
logic top_3_5_done;
logic [31:0] left_3_5_in;
logic left_3_5_write_en;
logic left_3_5_clk;
logic left_3_5_reset;
logic [31:0] left_3_5_out;
logic left_3_5_done;
logic [31:0] pe_3_6_top;
logic [31:0] pe_3_6_left;
logic pe_3_6_mul_ready;
logic [31:0] pe_3_6_out;
logic pe_3_6_go;
logic pe_3_6_clk;
logic pe_3_6_reset;
logic pe_3_6_done;
logic [31:0] top_3_6_in;
logic top_3_6_write_en;
logic top_3_6_clk;
logic top_3_6_reset;
logic [31:0] top_3_6_out;
logic top_3_6_done;
logic [31:0] left_3_6_in;
logic left_3_6_write_en;
logic left_3_6_clk;
logic left_3_6_reset;
logic [31:0] left_3_6_out;
logic left_3_6_done;
logic [31:0] pe_3_7_top;
logic [31:0] pe_3_7_left;
logic pe_3_7_mul_ready;
logic [31:0] pe_3_7_out;
logic pe_3_7_go;
logic pe_3_7_clk;
logic pe_3_7_reset;
logic pe_3_7_done;
logic [31:0] top_3_7_in;
logic top_3_7_write_en;
logic top_3_7_clk;
logic top_3_7_reset;
logic [31:0] top_3_7_out;
logic top_3_7_done;
logic [31:0] left_3_7_in;
logic left_3_7_write_en;
logic left_3_7_clk;
logic left_3_7_reset;
logic [31:0] left_3_7_out;
logic left_3_7_done;
logic [31:0] pe_4_0_top;
logic [31:0] pe_4_0_left;
logic pe_4_0_mul_ready;
logic [31:0] pe_4_0_out;
logic pe_4_0_go;
logic pe_4_0_clk;
logic pe_4_0_reset;
logic pe_4_0_done;
logic [31:0] top_4_0_in;
logic top_4_0_write_en;
logic top_4_0_clk;
logic top_4_0_reset;
logic [31:0] top_4_0_out;
logic top_4_0_done;
logic [31:0] left_4_0_in;
logic left_4_0_write_en;
logic left_4_0_clk;
logic left_4_0_reset;
logic [31:0] left_4_0_out;
logic left_4_0_done;
logic [31:0] pe_4_1_top;
logic [31:0] pe_4_1_left;
logic pe_4_1_mul_ready;
logic [31:0] pe_4_1_out;
logic pe_4_1_go;
logic pe_4_1_clk;
logic pe_4_1_reset;
logic pe_4_1_done;
logic [31:0] top_4_1_in;
logic top_4_1_write_en;
logic top_4_1_clk;
logic top_4_1_reset;
logic [31:0] top_4_1_out;
logic top_4_1_done;
logic [31:0] left_4_1_in;
logic left_4_1_write_en;
logic left_4_1_clk;
logic left_4_1_reset;
logic [31:0] left_4_1_out;
logic left_4_1_done;
logic [31:0] pe_4_2_top;
logic [31:0] pe_4_2_left;
logic pe_4_2_mul_ready;
logic [31:0] pe_4_2_out;
logic pe_4_2_go;
logic pe_4_2_clk;
logic pe_4_2_reset;
logic pe_4_2_done;
logic [31:0] top_4_2_in;
logic top_4_2_write_en;
logic top_4_2_clk;
logic top_4_2_reset;
logic [31:0] top_4_2_out;
logic top_4_2_done;
logic [31:0] left_4_2_in;
logic left_4_2_write_en;
logic left_4_2_clk;
logic left_4_2_reset;
logic [31:0] left_4_2_out;
logic left_4_2_done;
logic [31:0] pe_4_3_top;
logic [31:0] pe_4_3_left;
logic pe_4_3_mul_ready;
logic [31:0] pe_4_3_out;
logic pe_4_3_go;
logic pe_4_3_clk;
logic pe_4_3_reset;
logic pe_4_3_done;
logic [31:0] top_4_3_in;
logic top_4_3_write_en;
logic top_4_3_clk;
logic top_4_3_reset;
logic [31:0] top_4_3_out;
logic top_4_3_done;
logic [31:0] left_4_3_in;
logic left_4_3_write_en;
logic left_4_3_clk;
logic left_4_3_reset;
logic [31:0] left_4_3_out;
logic left_4_3_done;
logic [31:0] pe_4_4_top;
logic [31:0] pe_4_4_left;
logic pe_4_4_mul_ready;
logic [31:0] pe_4_4_out;
logic pe_4_4_go;
logic pe_4_4_clk;
logic pe_4_4_reset;
logic pe_4_4_done;
logic [31:0] top_4_4_in;
logic top_4_4_write_en;
logic top_4_4_clk;
logic top_4_4_reset;
logic [31:0] top_4_4_out;
logic top_4_4_done;
logic [31:0] left_4_4_in;
logic left_4_4_write_en;
logic left_4_4_clk;
logic left_4_4_reset;
logic [31:0] left_4_4_out;
logic left_4_4_done;
logic [31:0] pe_4_5_top;
logic [31:0] pe_4_5_left;
logic pe_4_5_mul_ready;
logic [31:0] pe_4_5_out;
logic pe_4_5_go;
logic pe_4_5_clk;
logic pe_4_5_reset;
logic pe_4_5_done;
logic [31:0] top_4_5_in;
logic top_4_5_write_en;
logic top_4_5_clk;
logic top_4_5_reset;
logic [31:0] top_4_5_out;
logic top_4_5_done;
logic [31:0] left_4_5_in;
logic left_4_5_write_en;
logic left_4_5_clk;
logic left_4_5_reset;
logic [31:0] left_4_5_out;
logic left_4_5_done;
logic [31:0] pe_4_6_top;
logic [31:0] pe_4_6_left;
logic pe_4_6_mul_ready;
logic [31:0] pe_4_6_out;
logic pe_4_6_go;
logic pe_4_6_clk;
logic pe_4_6_reset;
logic pe_4_6_done;
logic [31:0] top_4_6_in;
logic top_4_6_write_en;
logic top_4_6_clk;
logic top_4_6_reset;
logic [31:0] top_4_6_out;
logic top_4_6_done;
logic [31:0] left_4_6_in;
logic left_4_6_write_en;
logic left_4_6_clk;
logic left_4_6_reset;
logic [31:0] left_4_6_out;
logic left_4_6_done;
logic [31:0] pe_4_7_top;
logic [31:0] pe_4_7_left;
logic pe_4_7_mul_ready;
logic [31:0] pe_4_7_out;
logic pe_4_7_go;
logic pe_4_7_clk;
logic pe_4_7_reset;
logic pe_4_7_done;
logic [31:0] top_4_7_in;
logic top_4_7_write_en;
logic top_4_7_clk;
logic top_4_7_reset;
logic [31:0] top_4_7_out;
logic top_4_7_done;
logic [31:0] left_4_7_in;
logic left_4_7_write_en;
logic left_4_7_clk;
logic left_4_7_reset;
logic [31:0] left_4_7_out;
logic left_4_7_done;
logic [31:0] pe_5_0_top;
logic [31:0] pe_5_0_left;
logic pe_5_0_mul_ready;
logic [31:0] pe_5_0_out;
logic pe_5_0_go;
logic pe_5_0_clk;
logic pe_5_0_reset;
logic pe_5_0_done;
logic [31:0] top_5_0_in;
logic top_5_0_write_en;
logic top_5_0_clk;
logic top_5_0_reset;
logic [31:0] top_5_0_out;
logic top_5_0_done;
logic [31:0] left_5_0_in;
logic left_5_0_write_en;
logic left_5_0_clk;
logic left_5_0_reset;
logic [31:0] left_5_0_out;
logic left_5_0_done;
logic [31:0] pe_5_1_top;
logic [31:0] pe_5_1_left;
logic pe_5_1_mul_ready;
logic [31:0] pe_5_1_out;
logic pe_5_1_go;
logic pe_5_1_clk;
logic pe_5_1_reset;
logic pe_5_1_done;
logic [31:0] top_5_1_in;
logic top_5_1_write_en;
logic top_5_1_clk;
logic top_5_1_reset;
logic [31:0] top_5_1_out;
logic top_5_1_done;
logic [31:0] left_5_1_in;
logic left_5_1_write_en;
logic left_5_1_clk;
logic left_5_1_reset;
logic [31:0] left_5_1_out;
logic left_5_1_done;
logic [31:0] pe_5_2_top;
logic [31:0] pe_5_2_left;
logic pe_5_2_mul_ready;
logic [31:0] pe_5_2_out;
logic pe_5_2_go;
logic pe_5_2_clk;
logic pe_5_2_reset;
logic pe_5_2_done;
logic [31:0] top_5_2_in;
logic top_5_2_write_en;
logic top_5_2_clk;
logic top_5_2_reset;
logic [31:0] top_5_2_out;
logic top_5_2_done;
logic [31:0] left_5_2_in;
logic left_5_2_write_en;
logic left_5_2_clk;
logic left_5_2_reset;
logic [31:0] left_5_2_out;
logic left_5_2_done;
logic [31:0] pe_5_3_top;
logic [31:0] pe_5_3_left;
logic pe_5_3_mul_ready;
logic [31:0] pe_5_3_out;
logic pe_5_3_go;
logic pe_5_3_clk;
logic pe_5_3_reset;
logic pe_5_3_done;
logic [31:0] top_5_3_in;
logic top_5_3_write_en;
logic top_5_3_clk;
logic top_5_3_reset;
logic [31:0] top_5_3_out;
logic top_5_3_done;
logic [31:0] left_5_3_in;
logic left_5_3_write_en;
logic left_5_3_clk;
logic left_5_3_reset;
logic [31:0] left_5_3_out;
logic left_5_3_done;
logic [31:0] pe_5_4_top;
logic [31:0] pe_5_4_left;
logic pe_5_4_mul_ready;
logic [31:0] pe_5_4_out;
logic pe_5_4_go;
logic pe_5_4_clk;
logic pe_5_4_reset;
logic pe_5_4_done;
logic [31:0] top_5_4_in;
logic top_5_4_write_en;
logic top_5_4_clk;
logic top_5_4_reset;
logic [31:0] top_5_4_out;
logic top_5_4_done;
logic [31:0] left_5_4_in;
logic left_5_4_write_en;
logic left_5_4_clk;
logic left_5_4_reset;
logic [31:0] left_5_4_out;
logic left_5_4_done;
logic [31:0] pe_5_5_top;
logic [31:0] pe_5_5_left;
logic pe_5_5_mul_ready;
logic [31:0] pe_5_5_out;
logic pe_5_5_go;
logic pe_5_5_clk;
logic pe_5_5_reset;
logic pe_5_5_done;
logic [31:0] top_5_5_in;
logic top_5_5_write_en;
logic top_5_5_clk;
logic top_5_5_reset;
logic [31:0] top_5_5_out;
logic top_5_5_done;
logic [31:0] left_5_5_in;
logic left_5_5_write_en;
logic left_5_5_clk;
logic left_5_5_reset;
logic [31:0] left_5_5_out;
logic left_5_5_done;
logic [31:0] pe_5_6_top;
logic [31:0] pe_5_6_left;
logic pe_5_6_mul_ready;
logic [31:0] pe_5_6_out;
logic pe_5_6_go;
logic pe_5_6_clk;
logic pe_5_6_reset;
logic pe_5_6_done;
logic [31:0] top_5_6_in;
logic top_5_6_write_en;
logic top_5_6_clk;
logic top_5_6_reset;
logic [31:0] top_5_6_out;
logic top_5_6_done;
logic [31:0] left_5_6_in;
logic left_5_6_write_en;
logic left_5_6_clk;
logic left_5_6_reset;
logic [31:0] left_5_6_out;
logic left_5_6_done;
logic [31:0] pe_5_7_top;
logic [31:0] pe_5_7_left;
logic pe_5_7_mul_ready;
logic [31:0] pe_5_7_out;
logic pe_5_7_go;
logic pe_5_7_clk;
logic pe_5_7_reset;
logic pe_5_7_done;
logic [31:0] top_5_7_in;
logic top_5_7_write_en;
logic top_5_7_clk;
logic top_5_7_reset;
logic [31:0] top_5_7_out;
logic top_5_7_done;
logic [31:0] left_5_7_in;
logic left_5_7_write_en;
logic left_5_7_clk;
logic left_5_7_reset;
logic [31:0] left_5_7_out;
logic left_5_7_done;
logic [31:0] pe_6_0_top;
logic [31:0] pe_6_0_left;
logic pe_6_0_mul_ready;
logic [31:0] pe_6_0_out;
logic pe_6_0_go;
logic pe_6_0_clk;
logic pe_6_0_reset;
logic pe_6_0_done;
logic [31:0] top_6_0_in;
logic top_6_0_write_en;
logic top_6_0_clk;
logic top_6_0_reset;
logic [31:0] top_6_0_out;
logic top_6_0_done;
logic [31:0] left_6_0_in;
logic left_6_0_write_en;
logic left_6_0_clk;
logic left_6_0_reset;
logic [31:0] left_6_0_out;
logic left_6_0_done;
logic [31:0] pe_6_1_top;
logic [31:0] pe_6_1_left;
logic pe_6_1_mul_ready;
logic [31:0] pe_6_1_out;
logic pe_6_1_go;
logic pe_6_1_clk;
logic pe_6_1_reset;
logic pe_6_1_done;
logic [31:0] top_6_1_in;
logic top_6_1_write_en;
logic top_6_1_clk;
logic top_6_1_reset;
logic [31:0] top_6_1_out;
logic top_6_1_done;
logic [31:0] left_6_1_in;
logic left_6_1_write_en;
logic left_6_1_clk;
logic left_6_1_reset;
logic [31:0] left_6_1_out;
logic left_6_1_done;
logic [31:0] pe_6_2_top;
logic [31:0] pe_6_2_left;
logic pe_6_2_mul_ready;
logic [31:0] pe_6_2_out;
logic pe_6_2_go;
logic pe_6_2_clk;
logic pe_6_2_reset;
logic pe_6_2_done;
logic [31:0] top_6_2_in;
logic top_6_2_write_en;
logic top_6_2_clk;
logic top_6_2_reset;
logic [31:0] top_6_2_out;
logic top_6_2_done;
logic [31:0] left_6_2_in;
logic left_6_2_write_en;
logic left_6_2_clk;
logic left_6_2_reset;
logic [31:0] left_6_2_out;
logic left_6_2_done;
logic [31:0] pe_6_3_top;
logic [31:0] pe_6_3_left;
logic pe_6_3_mul_ready;
logic [31:0] pe_6_3_out;
logic pe_6_3_go;
logic pe_6_3_clk;
logic pe_6_3_reset;
logic pe_6_3_done;
logic [31:0] top_6_3_in;
logic top_6_3_write_en;
logic top_6_3_clk;
logic top_6_3_reset;
logic [31:0] top_6_3_out;
logic top_6_3_done;
logic [31:0] left_6_3_in;
logic left_6_3_write_en;
logic left_6_3_clk;
logic left_6_3_reset;
logic [31:0] left_6_3_out;
logic left_6_3_done;
logic [31:0] pe_6_4_top;
logic [31:0] pe_6_4_left;
logic pe_6_4_mul_ready;
logic [31:0] pe_6_4_out;
logic pe_6_4_go;
logic pe_6_4_clk;
logic pe_6_4_reset;
logic pe_6_4_done;
logic [31:0] top_6_4_in;
logic top_6_4_write_en;
logic top_6_4_clk;
logic top_6_4_reset;
logic [31:0] top_6_4_out;
logic top_6_4_done;
logic [31:0] left_6_4_in;
logic left_6_4_write_en;
logic left_6_4_clk;
logic left_6_4_reset;
logic [31:0] left_6_4_out;
logic left_6_4_done;
logic [31:0] pe_6_5_top;
logic [31:0] pe_6_5_left;
logic pe_6_5_mul_ready;
logic [31:0] pe_6_5_out;
logic pe_6_5_go;
logic pe_6_5_clk;
logic pe_6_5_reset;
logic pe_6_5_done;
logic [31:0] top_6_5_in;
logic top_6_5_write_en;
logic top_6_5_clk;
logic top_6_5_reset;
logic [31:0] top_6_5_out;
logic top_6_5_done;
logic [31:0] left_6_5_in;
logic left_6_5_write_en;
logic left_6_5_clk;
logic left_6_5_reset;
logic [31:0] left_6_5_out;
logic left_6_5_done;
logic [31:0] pe_6_6_top;
logic [31:0] pe_6_6_left;
logic pe_6_6_mul_ready;
logic [31:0] pe_6_6_out;
logic pe_6_6_go;
logic pe_6_6_clk;
logic pe_6_6_reset;
logic pe_6_6_done;
logic [31:0] top_6_6_in;
logic top_6_6_write_en;
logic top_6_6_clk;
logic top_6_6_reset;
logic [31:0] top_6_6_out;
logic top_6_6_done;
logic [31:0] left_6_6_in;
logic left_6_6_write_en;
logic left_6_6_clk;
logic left_6_6_reset;
logic [31:0] left_6_6_out;
logic left_6_6_done;
logic [31:0] pe_6_7_top;
logic [31:0] pe_6_7_left;
logic pe_6_7_mul_ready;
logic [31:0] pe_6_7_out;
logic pe_6_7_go;
logic pe_6_7_clk;
logic pe_6_7_reset;
logic pe_6_7_done;
logic [31:0] top_6_7_in;
logic top_6_7_write_en;
logic top_6_7_clk;
logic top_6_7_reset;
logic [31:0] top_6_7_out;
logic top_6_7_done;
logic [31:0] left_6_7_in;
logic left_6_7_write_en;
logic left_6_7_clk;
logic left_6_7_reset;
logic [31:0] left_6_7_out;
logic left_6_7_done;
logic [31:0] pe_7_0_top;
logic [31:0] pe_7_0_left;
logic pe_7_0_mul_ready;
logic [31:0] pe_7_0_out;
logic pe_7_0_go;
logic pe_7_0_clk;
logic pe_7_0_reset;
logic pe_7_0_done;
logic [31:0] top_7_0_in;
logic top_7_0_write_en;
logic top_7_0_clk;
logic top_7_0_reset;
logic [31:0] top_7_0_out;
logic top_7_0_done;
logic [31:0] left_7_0_in;
logic left_7_0_write_en;
logic left_7_0_clk;
logic left_7_0_reset;
logic [31:0] left_7_0_out;
logic left_7_0_done;
logic [31:0] pe_7_1_top;
logic [31:0] pe_7_1_left;
logic pe_7_1_mul_ready;
logic [31:0] pe_7_1_out;
logic pe_7_1_go;
logic pe_7_1_clk;
logic pe_7_1_reset;
logic pe_7_1_done;
logic [31:0] top_7_1_in;
logic top_7_1_write_en;
logic top_7_1_clk;
logic top_7_1_reset;
logic [31:0] top_7_1_out;
logic top_7_1_done;
logic [31:0] left_7_1_in;
logic left_7_1_write_en;
logic left_7_1_clk;
logic left_7_1_reset;
logic [31:0] left_7_1_out;
logic left_7_1_done;
logic [31:0] pe_7_2_top;
logic [31:0] pe_7_2_left;
logic pe_7_2_mul_ready;
logic [31:0] pe_7_2_out;
logic pe_7_2_go;
logic pe_7_2_clk;
logic pe_7_2_reset;
logic pe_7_2_done;
logic [31:0] top_7_2_in;
logic top_7_2_write_en;
logic top_7_2_clk;
logic top_7_2_reset;
logic [31:0] top_7_2_out;
logic top_7_2_done;
logic [31:0] left_7_2_in;
logic left_7_2_write_en;
logic left_7_2_clk;
logic left_7_2_reset;
logic [31:0] left_7_2_out;
logic left_7_2_done;
logic [31:0] pe_7_3_top;
logic [31:0] pe_7_3_left;
logic pe_7_3_mul_ready;
logic [31:0] pe_7_3_out;
logic pe_7_3_go;
logic pe_7_3_clk;
logic pe_7_3_reset;
logic pe_7_3_done;
logic [31:0] top_7_3_in;
logic top_7_3_write_en;
logic top_7_3_clk;
logic top_7_3_reset;
logic [31:0] top_7_3_out;
logic top_7_3_done;
logic [31:0] left_7_3_in;
logic left_7_3_write_en;
logic left_7_3_clk;
logic left_7_3_reset;
logic [31:0] left_7_3_out;
logic left_7_3_done;
logic [31:0] pe_7_4_top;
logic [31:0] pe_7_4_left;
logic pe_7_4_mul_ready;
logic [31:0] pe_7_4_out;
logic pe_7_4_go;
logic pe_7_4_clk;
logic pe_7_4_reset;
logic pe_7_4_done;
logic [31:0] top_7_4_in;
logic top_7_4_write_en;
logic top_7_4_clk;
logic top_7_4_reset;
logic [31:0] top_7_4_out;
logic top_7_4_done;
logic [31:0] left_7_4_in;
logic left_7_4_write_en;
logic left_7_4_clk;
logic left_7_4_reset;
logic [31:0] left_7_4_out;
logic left_7_4_done;
logic [31:0] pe_7_5_top;
logic [31:0] pe_7_5_left;
logic pe_7_5_mul_ready;
logic [31:0] pe_7_5_out;
logic pe_7_5_go;
logic pe_7_5_clk;
logic pe_7_5_reset;
logic pe_7_5_done;
logic [31:0] top_7_5_in;
logic top_7_5_write_en;
logic top_7_5_clk;
logic top_7_5_reset;
logic [31:0] top_7_5_out;
logic top_7_5_done;
logic [31:0] left_7_5_in;
logic left_7_5_write_en;
logic left_7_5_clk;
logic left_7_5_reset;
logic [31:0] left_7_5_out;
logic left_7_5_done;
logic [31:0] pe_7_6_top;
logic [31:0] pe_7_6_left;
logic pe_7_6_mul_ready;
logic [31:0] pe_7_6_out;
logic pe_7_6_go;
logic pe_7_6_clk;
logic pe_7_6_reset;
logic pe_7_6_done;
logic [31:0] top_7_6_in;
logic top_7_6_write_en;
logic top_7_6_clk;
logic top_7_6_reset;
logic [31:0] top_7_6_out;
logic top_7_6_done;
logic [31:0] left_7_6_in;
logic left_7_6_write_en;
logic left_7_6_clk;
logic left_7_6_reset;
logic [31:0] left_7_6_out;
logic left_7_6_done;
logic [31:0] pe_7_7_top;
logic [31:0] pe_7_7_left;
logic pe_7_7_mul_ready;
logic [31:0] pe_7_7_out;
logic pe_7_7_go;
logic pe_7_7_clk;
logic pe_7_7_reset;
logic pe_7_7_done;
logic [31:0] top_7_7_in;
logic top_7_7_write_en;
logic top_7_7_clk;
logic top_7_7_reset;
logic [31:0] top_7_7_out;
logic top_7_7_done;
logic [31:0] left_7_7_in;
logic left_7_7_write_en;
logic left_7_7_clk;
logic left_7_7_reset;
logic [31:0] left_7_7_out;
logic left_7_7_done;
logic [3:0] t0_idx_in;
logic t0_idx_write_en;
logic t0_idx_clk;
logic t0_idx_reset;
logic [3:0] t0_idx_out;
logic t0_idx_done;
logic [3:0] t0_add_left;
logic [3:0] t0_add_right;
logic [3:0] t0_add_out;
logic [3:0] t1_idx_in;
logic t1_idx_write_en;
logic t1_idx_clk;
logic t1_idx_reset;
logic [3:0] t1_idx_out;
logic t1_idx_done;
logic [3:0] t1_add_left;
logic [3:0] t1_add_right;
logic [3:0] t1_add_out;
logic [3:0] t2_idx_in;
logic t2_idx_write_en;
logic t2_idx_clk;
logic t2_idx_reset;
logic [3:0] t2_idx_out;
logic t2_idx_done;
logic [3:0] t2_add_left;
logic [3:0] t2_add_right;
logic [3:0] t2_add_out;
logic [3:0] t3_idx_in;
logic t3_idx_write_en;
logic t3_idx_clk;
logic t3_idx_reset;
logic [3:0] t3_idx_out;
logic t3_idx_done;
logic [3:0] t3_add_left;
logic [3:0] t3_add_right;
logic [3:0] t3_add_out;
logic [3:0] t4_idx_in;
logic t4_idx_write_en;
logic t4_idx_clk;
logic t4_idx_reset;
logic [3:0] t4_idx_out;
logic t4_idx_done;
logic [3:0] t4_add_left;
logic [3:0] t4_add_right;
logic [3:0] t4_add_out;
logic [3:0] t5_idx_in;
logic t5_idx_write_en;
logic t5_idx_clk;
logic t5_idx_reset;
logic [3:0] t5_idx_out;
logic t5_idx_done;
logic [3:0] t5_add_left;
logic [3:0] t5_add_right;
logic [3:0] t5_add_out;
logic [3:0] t6_idx_in;
logic t6_idx_write_en;
logic t6_idx_clk;
logic t6_idx_reset;
logic [3:0] t6_idx_out;
logic t6_idx_done;
logic [3:0] t6_add_left;
logic [3:0] t6_add_right;
logic [3:0] t6_add_out;
logic [3:0] t7_idx_in;
logic t7_idx_write_en;
logic t7_idx_clk;
logic t7_idx_reset;
logic [3:0] t7_idx_out;
logic t7_idx_done;
logic [3:0] t7_add_left;
logic [3:0] t7_add_right;
logic [3:0] t7_add_out;
logic [3:0] l0_idx_in;
logic l0_idx_write_en;
logic l0_idx_clk;
logic l0_idx_reset;
logic [3:0] l0_idx_out;
logic l0_idx_done;
logic [3:0] l0_add_left;
logic [3:0] l0_add_right;
logic [3:0] l0_add_out;
logic [3:0] l1_idx_in;
logic l1_idx_write_en;
logic l1_idx_clk;
logic l1_idx_reset;
logic [3:0] l1_idx_out;
logic l1_idx_done;
logic [3:0] l1_add_left;
logic [3:0] l1_add_right;
logic [3:0] l1_add_out;
logic [3:0] l2_idx_in;
logic l2_idx_write_en;
logic l2_idx_clk;
logic l2_idx_reset;
logic [3:0] l2_idx_out;
logic l2_idx_done;
logic [3:0] l2_add_left;
logic [3:0] l2_add_right;
logic [3:0] l2_add_out;
logic [3:0] l3_idx_in;
logic l3_idx_write_en;
logic l3_idx_clk;
logic l3_idx_reset;
logic [3:0] l3_idx_out;
logic l3_idx_done;
logic [3:0] l3_add_left;
logic [3:0] l3_add_right;
logic [3:0] l3_add_out;
logic [3:0] l4_idx_in;
logic l4_idx_write_en;
logic l4_idx_clk;
logic l4_idx_reset;
logic [3:0] l4_idx_out;
logic l4_idx_done;
logic [3:0] l4_add_left;
logic [3:0] l4_add_right;
logic [3:0] l4_add_out;
logic [3:0] l5_idx_in;
logic l5_idx_write_en;
logic l5_idx_clk;
logic l5_idx_reset;
logic [3:0] l5_idx_out;
logic l5_idx_done;
logic [3:0] l5_add_left;
logic [3:0] l5_add_right;
logic [3:0] l5_add_out;
logic [3:0] l6_idx_in;
logic l6_idx_write_en;
logic l6_idx_clk;
logic l6_idx_reset;
logic [3:0] l6_idx_out;
logic l6_idx_done;
logic [3:0] l6_add_left;
logic [3:0] l6_add_right;
logic [3:0] l6_add_out;
logic [3:0] l7_idx_in;
logic l7_idx_write_en;
logic l7_idx_clk;
logic l7_idx_reset;
logic [3:0] l7_idx_out;
logic l7_idx_done;
logic [3:0] l7_add_left;
logic [3:0] l7_add_right;
logic [3:0] l7_add_out;
logic [4:0] idx_in;
logic idx_write_en;
logic idx_clk;
logic idx_reset;
logic [4:0] idx_out;
logic idx_done;
logic [4:0] idx_add_left;
logic [4:0] idx_add_right;
logic [4:0] idx_add_out;
logic idx_between_18_26_reg_in;
logic idx_between_18_26_reg_write_en;
logic idx_between_18_26_reg_clk;
logic idx_between_18_26_reg_reset;
logic idx_between_18_26_reg_out;
logic idx_between_18_26_reg_done;
logic [4:0] index_lt_26_left;
logic [4:0] index_lt_26_right;
logic index_lt_26_out;
logic [4:0] index_ge_18_left;
logic [4:0] index_ge_18_right;
logic index_ge_18_out;
logic idx_between_18_26_comb_left;
logic idx_between_18_26_comb_right;
logic idx_between_18_26_comb_out;
logic idx_between_3_7_reg_in;
logic idx_between_3_7_reg_write_en;
logic idx_between_3_7_reg_clk;
logic idx_between_3_7_reg_reset;
logic idx_between_3_7_reg_out;
logic idx_between_3_7_reg_done;
logic [4:0] index_lt_7_left;
logic [4:0] index_lt_7_right;
logic index_lt_7_out;
logic [4:0] index_ge_3_left;
logic [4:0] index_ge_3_right;
logic index_ge_3_out;
logic idx_between_3_7_comb_left;
logic idx_between_3_7_comb_right;
logic idx_between_3_7_comb_out;
logic idx_between_12_16_reg_in;
logic idx_between_12_16_reg_write_en;
logic idx_between_12_16_reg_clk;
logic idx_between_12_16_reg_reset;
logic idx_between_12_16_reg_out;
logic idx_between_12_16_reg_done;
logic [4:0] index_lt_16_left;
logic [4:0] index_lt_16_right;
logic index_lt_16_out;
logic [4:0] index_ge_12_left;
logic [4:0] index_ge_12_right;
logic index_ge_12_out;
logic idx_between_12_16_comb_left;
logic idx_between_12_16_comb_right;
logic idx_between_12_16_comb_out;
logic idx_between_26_27_reg_in;
logic idx_between_26_27_reg_write_en;
logic idx_between_26_27_reg_clk;
logic idx_between_26_27_reg_reset;
logic idx_between_26_27_reg_out;
logic idx_between_26_27_reg_done;
logic [4:0] index_lt_27_left;
logic [4:0] index_lt_27_right;
logic index_lt_27_out;
logic [4:0] index_ge_26_left;
logic [4:0] index_ge_26_right;
logic index_ge_26_out;
logic idx_between_26_27_comb_left;
logic idx_between_26_27_comb_right;
logic idx_between_26_27_comb_out;
logic idx_between_4_12_reg_in;
logic idx_between_4_12_reg_write_en;
logic idx_between_4_12_reg_clk;
logic idx_between_4_12_reg_reset;
logic idx_between_4_12_reg_out;
logic idx_between_4_12_reg_done;
logic [4:0] index_lt_12_left;
logic [4:0] index_lt_12_right;
logic index_lt_12_out;
logic [4:0] index_ge_4_left;
logic [4:0] index_ge_4_right;
logic index_ge_4_out;
logic idx_between_4_12_comb_left;
logic idx_between_4_12_comb_right;
logic idx_between_4_12_comb_out;
logic idx_between_21_22_reg_in;
logic idx_between_21_22_reg_write_en;
logic idx_between_21_22_reg_clk;
logic idx_between_21_22_reg_reset;
logic idx_between_21_22_reg_out;
logic idx_between_21_22_reg_done;
logic [4:0] index_lt_22_left;
logic [4:0] index_lt_22_right;
logic index_lt_22_out;
logic [4:0] index_ge_21_left;
logic [4:0] index_ge_21_right;
logic index_ge_21_out;
logic idx_between_21_22_comb_left;
logic idx_between_21_22_comb_right;
logic idx_between_21_22_comb_out;
logic idx_between_5_13_reg_in;
logic idx_between_5_13_reg_write_en;
logic idx_between_5_13_reg_clk;
logic idx_between_5_13_reg_reset;
logic idx_between_5_13_reg_out;
logic idx_between_5_13_reg_done;
logic [4:0] index_lt_13_left;
logic [4:0] index_lt_13_right;
logic index_lt_13_out;
logic [4:0] index_ge_5_left;
logic [4:0] index_ge_5_right;
logic index_ge_5_out;
logic idx_between_5_13_comb_left;
logic idx_between_5_13_comb_right;
logic idx_between_5_13_comb_out;
logic idx_between_22_23_reg_in;
logic idx_between_22_23_reg_write_en;
logic idx_between_22_23_reg_clk;
logic idx_between_22_23_reg_reset;
logic idx_between_22_23_reg_out;
logic idx_between_22_23_reg_done;
logic [4:0] index_lt_23_left;
logic [4:0] index_lt_23_right;
logic index_lt_23_out;
logic [4:0] index_ge_22_left;
logic [4:0] index_ge_22_right;
logic index_ge_22_out;
logic idx_between_22_23_comb_left;
logic idx_between_22_23_comb_right;
logic idx_between_22_23_comb_out;
logic idx_between_14_22_reg_in;
logic idx_between_14_22_reg_write_en;
logic idx_between_14_22_reg_clk;
logic idx_between_14_22_reg_reset;
logic idx_between_14_22_reg_out;
logic idx_between_14_22_reg_done;
logic [4:0] index_ge_14_left;
logic [4:0] index_ge_14_right;
logic index_ge_14_out;
logic idx_between_14_22_comb_left;
logic idx_between_14_22_comb_right;
logic idx_between_14_22_comb_out;
logic idx_between_8_12_reg_in;
logic idx_between_8_12_reg_write_en;
logic idx_between_8_12_reg_clk;
logic idx_between_8_12_reg_reset;
logic idx_between_8_12_reg_out;
logic idx_between_8_12_reg_done;
logic [4:0] index_ge_8_left;
logic [4:0] index_ge_8_right;
logic index_ge_8_out;
logic idx_between_8_12_comb_left;
logic idx_between_8_12_comb_right;
logic idx_between_8_12_comb_out;
logic idx_between_9_17_reg_in;
logic idx_between_9_17_reg_write_en;
logic idx_between_9_17_reg_clk;
logic idx_between_9_17_reg_reset;
logic idx_between_9_17_reg_out;
logic idx_between_9_17_reg_done;
logic [4:0] index_lt_17_left;
logic [4:0] index_lt_17_right;
logic index_lt_17_out;
logic [4:0] index_ge_9_left;
logic [4:0] index_ge_9_right;
logic index_ge_9_out;
logic idx_between_9_17_comb_left;
logic idx_between_9_17_comb_right;
logic idx_between_9_17_comb_out;
logic idx_between_0_8_reg_in;
logic idx_between_0_8_reg_write_en;
logic idx_between_0_8_reg_clk;
logic idx_between_0_8_reg_reset;
logic idx_between_0_8_reg_out;
logic idx_between_0_8_reg_done;
logic [4:0] index_lt_8_left;
logic [4:0] index_lt_8_right;
logic index_lt_8_out;
logic idx_between_17_18_reg_in;
logic idx_between_17_18_reg_write_en;
logic idx_between_17_18_reg_clk;
logic idx_between_17_18_reg_reset;
logic idx_between_17_18_reg_out;
logic idx_between_17_18_reg_done;
logic [4:0] index_lt_18_left;
logic [4:0] index_lt_18_right;
logic index_lt_18_out;
logic [4:0] index_ge_17_left;
logic [4:0] index_ge_17_right;
logic index_ge_17_out;
logic idx_between_17_18_comb_left;
logic idx_between_17_18_comb_right;
logic idx_between_17_18_comb_out;
logic idx_between_1_9_reg_in;
logic idx_between_1_9_reg_write_en;
logic idx_between_1_9_reg_clk;
logic idx_between_1_9_reg_reset;
logic idx_between_1_9_reg_out;
logic idx_between_1_9_reg_done;
logic [4:0] index_lt_9_left;
logic [4:0] index_lt_9_right;
logic index_lt_9_out;
logic [4:0] index_ge_1_left;
logic [4:0] index_ge_1_right;
logic index_ge_1_out;
logic idx_between_1_9_comb_left;
logic idx_between_1_9_comb_right;
logic idx_between_1_9_comb_out;
logic idx_between_10_18_reg_in;
logic idx_between_10_18_reg_write_en;
logic idx_between_10_18_reg_clk;
logic idx_between_10_18_reg_reset;
logic idx_between_10_18_reg_out;
logic idx_between_10_18_reg_done;
logic [4:0] index_ge_10_left;
logic [4:0] index_ge_10_right;
logic index_ge_10_out;
logic idx_between_10_18_comb_left;
logic idx_between_10_18_comb_right;
logic idx_between_10_18_comb_out;
logic idx_between_25_26_reg_in;
logic idx_between_25_26_reg_write_en;
logic idx_between_25_26_reg_clk;
logic idx_between_25_26_reg_reset;
logic idx_between_25_26_reg_out;
logic idx_between_25_26_reg_done;
logic [4:0] index_ge_25_left;
logic [4:0] index_ge_25_right;
logic index_ge_25_out;
logic idx_between_25_26_comb_left;
logic idx_between_25_26_comb_right;
logic idx_between_25_26_comb_out;
logic idx_between_27_28_reg_in;
logic idx_between_27_28_reg_write_en;
logic idx_between_27_28_reg_clk;
logic idx_between_27_28_reg_reset;
logic idx_between_27_28_reg_out;
logic idx_between_27_28_reg_done;
logic [4:0] index_lt_28_left;
logic [4:0] index_lt_28_right;
logic index_lt_28_out;
logic [4:0] index_ge_27_left;
logic [4:0] index_ge_27_right;
logic index_ge_27_out;
logic idx_between_27_28_comb_left;
logic idx_between_27_28_comb_right;
logic idx_between_27_28_comb_out;
logic idx_between_13_14_reg_in;
logic idx_between_13_14_reg_write_en;
logic idx_between_13_14_reg_clk;
logic idx_between_13_14_reg_reset;
logic idx_between_13_14_reg_out;
logic idx_between_13_14_reg_done;
logic [4:0] index_lt_14_left;
logic [4:0] index_lt_14_right;
logic index_lt_14_out;
logic [4:0] index_ge_13_left;
logic [4:0] index_ge_13_right;
logic index_ge_13_out;
logic idx_between_13_14_comb_left;
logic idx_between_13_14_comb_right;
logic idx_between_13_14_comb_out;
logic idx_between_19_27_reg_in;
logic idx_between_19_27_reg_write_en;
logic idx_between_19_27_reg_clk;
logic idx_between_19_27_reg_reset;
logic idx_between_19_27_reg_out;
logic idx_between_19_27_reg_done;
logic [4:0] index_ge_19_left;
logic [4:0] index_ge_19_right;
logic index_ge_19_out;
logic idx_between_19_27_comb_left;
logic idx_between_19_27_comb_right;
logic idx_between_19_27_comb_out;
logic idx_between_13_17_reg_in;
logic idx_between_13_17_reg_write_en;
logic idx_between_13_17_reg_clk;
logic idx_between_13_17_reg_reset;
logic idx_between_13_17_reg_out;
logic idx_between_13_17_reg_done;
logic idx_between_13_17_comb_left;
logic idx_between_13_17_comb_right;
logic idx_between_13_17_comb_out;
logic idx_between_6_14_reg_in;
logic idx_between_6_14_reg_write_en;
logic idx_between_6_14_reg_clk;
logic idx_between_6_14_reg_reset;
logic idx_between_6_14_reg_out;
logic idx_between_6_14_reg_done;
logic [4:0] index_ge_6_left;
logic [4:0] index_ge_6_right;
logic index_ge_6_out;
logic idx_between_6_14_comb_left;
logic idx_between_6_14_comb_right;
logic idx_between_6_14_comb_out;
logic idx_between_15_23_reg_in;
logic idx_between_15_23_reg_write_en;
logic idx_between_15_23_reg_clk;
logic idx_between_15_23_reg_reset;
logic idx_between_15_23_reg_out;
logic idx_between_15_23_reg_done;
logic [4:0] index_ge_15_left;
logic [4:0] index_ge_15_right;
logic index_ge_15_out;
logic idx_between_15_23_comb_left;
logic idx_between_15_23_comb_right;
logic idx_between_15_23_comb_out;
logic idx_between_18_19_reg_in;
logic idx_between_18_19_reg_write_en;
logic idx_between_18_19_reg_clk;
logic idx_between_18_19_reg_reset;
logic idx_between_18_19_reg_out;
logic idx_between_18_19_reg_done;
logic [4:0] index_lt_19_left;
logic [4:0] index_lt_19_right;
logic index_lt_19_out;
logic idx_between_18_19_comb_left;
logic idx_between_18_19_comb_right;
logic idx_between_18_19_comb_out;
logic idx_between_4_8_reg_in;
logic idx_between_4_8_reg_write_en;
logic idx_between_4_8_reg_clk;
logic idx_between_4_8_reg_reset;
logic idx_between_4_8_reg_out;
logic idx_between_4_8_reg_done;
logic idx_between_4_8_comb_left;
logic idx_between_4_8_comb_right;
logic idx_between_4_8_comb_out;
logic idx_between_5_9_reg_in;
logic idx_between_5_9_reg_write_en;
logic idx_between_5_9_reg_clk;
logic idx_between_5_9_reg_reset;
logic idx_between_5_9_reg_out;
logic idx_between_5_9_reg_done;
logic idx_between_5_9_comb_left;
logic idx_between_5_9_comb_right;
logic idx_between_5_9_comb_out;
logic idx_between_14_18_reg_in;
logic idx_between_14_18_reg_write_en;
logic idx_between_14_18_reg_clk;
logic idx_between_14_18_reg_reset;
logic idx_between_14_18_reg_out;
logic idx_between_14_18_reg_done;
logic idx_between_14_18_comb_left;
logic idx_between_14_18_comb_right;
logic idx_between_14_18_comb_out;
logic idx_between_14_15_reg_in;
logic idx_between_14_15_reg_write_en;
logic idx_between_14_15_reg_clk;
logic idx_between_14_15_reg_reset;
logic idx_between_14_15_reg_out;
logic idx_between_14_15_reg_done;
logic [4:0] index_lt_15_left;
logic [4:0] index_lt_15_right;
logic index_lt_15_out;
logic idx_between_14_15_comb_left;
logic idx_between_14_15_comb_right;
logic idx_between_14_15_comb_out;
logic idx_between_23_24_reg_in;
logic idx_between_23_24_reg_write_en;
logic idx_between_23_24_reg_clk;
logic idx_between_23_24_reg_reset;
logic idx_between_23_24_reg_out;
logic idx_between_23_24_reg_done;
logic [4:0] index_lt_24_left;
logic [4:0] index_lt_24_right;
logic index_lt_24_out;
logic [4:0] index_ge_23_left;
logic [4:0] index_ge_23_right;
logic index_ge_23_out;
logic idx_between_23_24_comb_left;
logic idx_between_23_24_comb_right;
logic idx_between_23_24_comb_out;
logic idx_between_9_13_reg_in;
logic idx_between_9_13_reg_write_en;
logic idx_between_9_13_reg_clk;
logic idx_between_9_13_reg_reset;
logic idx_between_9_13_reg_out;
logic idx_between_9_13_reg_done;
logic idx_between_9_13_comb_left;
logic idx_between_9_13_comb_right;
logic idx_between_9_13_comb_out;
logic idx_between_1_5_reg_in;
logic idx_between_1_5_reg_write_en;
logic idx_between_1_5_reg_clk;
logic idx_between_1_5_reg_reset;
logic idx_between_1_5_reg_out;
logic idx_between_1_5_reg_done;
logic [4:0] index_lt_5_left;
logic [4:0] index_lt_5_right;
logic index_lt_5_out;
logic idx_between_1_5_comb_left;
logic idx_between_1_5_comb_right;
logic idx_between_1_5_comb_out;
logic idx_between_10_14_reg_in;
logic idx_between_10_14_reg_write_en;
logic idx_between_10_14_reg_clk;
logic idx_between_10_14_reg_reset;
logic idx_between_10_14_reg_out;
logic idx_between_10_14_reg_done;
logic idx_between_10_14_comb_left;
logic idx_between_10_14_comb_right;
logic idx_between_10_14_comb_out;
logic idx_between_2_10_reg_in;
logic idx_between_2_10_reg_write_en;
logic idx_between_2_10_reg_clk;
logic idx_between_2_10_reg_reset;
logic idx_between_2_10_reg_out;
logic idx_between_2_10_reg_done;
logic [4:0] index_lt_10_left;
logic [4:0] index_lt_10_right;
logic index_lt_10_out;
logic [4:0] index_ge_2_left;
logic [4:0] index_ge_2_right;
logic index_ge_2_out;
logic idx_between_2_10_comb_left;
logic idx_between_2_10_comb_right;
logic idx_between_2_10_comb_out;
logic idx_between_11_19_reg_in;
logic idx_between_11_19_reg_write_en;
logic idx_between_11_19_reg_clk;
logic idx_between_11_19_reg_reset;
logic idx_between_11_19_reg_out;
logic idx_between_11_19_reg_done;
logic [4:0] index_ge_11_left;
logic [4:0] index_ge_11_right;
logic index_ge_11_out;
logic idx_between_11_19_comb_left;
logic idx_between_11_19_comb_right;
logic idx_between_11_19_comb_out;
logic idx_between_19_20_reg_in;
logic idx_between_19_20_reg_write_en;
logic idx_between_19_20_reg_clk;
logic idx_between_19_20_reg_reset;
logic idx_between_19_20_reg_out;
logic idx_between_19_20_reg_done;
logic [4:0] index_lt_20_left;
logic [4:0] index_lt_20_right;
logic index_lt_20_out;
logic idx_between_19_20_comb_left;
logic idx_between_19_20_comb_right;
logic idx_between_19_20_comb_out;
logic idx_between_15_16_reg_in;
logic idx_between_15_16_reg_write_en;
logic idx_between_15_16_reg_clk;
logic idx_between_15_16_reg_reset;
logic idx_between_15_16_reg_out;
logic idx_between_15_16_reg_done;
logic idx_between_15_16_comb_left;
logic idx_between_15_16_comb_right;
logic idx_between_15_16_comb_out;
logic idx_between_24_25_reg_in;
logic idx_between_24_25_reg_write_en;
logic idx_between_24_25_reg_clk;
logic idx_between_24_25_reg_reset;
logic idx_between_24_25_reg_out;
logic idx_between_24_25_reg_done;
logic [4:0] index_lt_25_left;
logic [4:0] index_lt_25_right;
logic index_lt_25_out;
logic [4:0] index_ge_24_left;
logic [4:0] index_ge_24_right;
logic index_ge_24_out;
logic idx_between_24_25_comb_left;
logic idx_between_24_25_comb_right;
logic idx_between_24_25_comb_out;
logic idx_between_6_10_reg_in;
logic idx_between_6_10_reg_write_en;
logic idx_between_6_10_reg_clk;
logic idx_between_6_10_reg_reset;
logic idx_between_6_10_reg_out;
logic idx_between_6_10_reg_done;
logic idx_between_6_10_comb_left;
logic idx_between_6_10_comb_right;
logic idx_between_6_10_comb_out;
logic idx_between_15_19_reg_in;
logic idx_between_15_19_reg_write_en;
logic idx_between_15_19_reg_clk;
logic idx_between_15_19_reg_reset;
logic idx_between_15_19_reg_out;
logic idx_between_15_19_reg_done;
logic idx_between_15_19_comb_left;
logic idx_between_15_19_comb_right;
logic idx_between_15_19_comb_out;
logic idx_between_7_15_reg_in;
logic idx_between_7_15_reg_write_en;
logic idx_between_7_15_reg_clk;
logic idx_between_7_15_reg_reset;
logic idx_between_7_15_reg_out;
logic idx_between_7_15_reg_done;
logic [4:0] index_ge_7_left;
logic [4:0] index_ge_7_right;
logic index_ge_7_out;
logic idx_between_7_15_comb_left;
logic idx_between_7_15_comb_right;
logic idx_between_7_15_comb_out;
logic idx_between_16_24_reg_in;
logic idx_between_16_24_reg_write_en;
logic idx_between_16_24_reg_clk;
logic idx_between_16_24_reg_reset;
logic idx_between_16_24_reg_out;
logic idx_between_16_24_reg_done;
logic [4:0] index_ge_16_left;
logic [4:0] index_ge_16_right;
logic index_ge_16_out;
logic idx_between_16_24_comb_left;
logic idx_between_16_24_comb_right;
logic idx_between_16_24_comb_out;
logic idx_between_3_11_reg_in;
logic idx_between_3_11_reg_write_en;
logic idx_between_3_11_reg_clk;
logic idx_between_3_11_reg_reset;
logic idx_between_3_11_reg_out;
logic idx_between_3_11_reg_done;
logic [4:0] index_lt_11_left;
logic [4:0] index_lt_11_right;
logic index_lt_11_out;
logic idx_between_3_11_comb_left;
logic idx_between_3_11_comb_right;
logic idx_between_3_11_comb_out;
logic idx_between_20_21_reg_in;
logic idx_between_20_21_reg_write_en;
logic idx_between_20_21_reg_clk;
logic idx_between_20_21_reg_reset;
logic idx_between_20_21_reg_out;
logic idx_between_20_21_reg_done;
logic [4:0] index_lt_21_left;
logic [4:0] index_lt_21_right;
logic index_lt_21_out;
logic [4:0] index_ge_20_left;
logic [4:0] index_ge_20_right;
logic index_ge_20_out;
logic idx_between_20_21_comb_left;
logic idx_between_20_21_comb_right;
logic idx_between_20_21_comb_out;
logic idx_between_12_20_reg_in;
logic idx_between_12_20_reg_write_en;
logic idx_between_12_20_reg_clk;
logic idx_between_12_20_reg_reset;
logic idx_between_12_20_reg_out;
logic idx_between_12_20_reg_done;
logic idx_between_12_20_comb_left;
logic idx_between_12_20_comb_right;
logic idx_between_12_20_comb_out;
logic idx_between_8_16_reg_in;
logic idx_between_8_16_reg_write_en;
logic idx_between_8_16_reg_clk;
logic idx_between_8_16_reg_reset;
logic idx_between_8_16_reg_out;
logic idx_between_8_16_reg_done;
logic idx_between_8_16_comb_left;
logic idx_between_8_16_comb_right;
logic idx_between_8_16_comb_out;
logic idx_between_7_11_reg_in;
logic idx_between_7_11_reg_write_en;
logic idx_between_7_11_reg_clk;
logic idx_between_7_11_reg_reset;
logic idx_between_7_11_reg_out;
logic idx_between_7_11_reg_done;
logic idx_between_7_11_comb_left;
logic idx_between_7_11_comb_right;
logic idx_between_7_11_comb_out;
logic idx_between_2_6_reg_in;
logic idx_between_2_6_reg_write_en;
logic idx_between_2_6_reg_clk;
logic idx_between_2_6_reg_reset;
logic idx_between_2_6_reg_out;
logic idx_between_2_6_reg_done;
logic [4:0] index_lt_6_left;
logic [4:0] index_lt_6_right;
logic index_lt_6_out;
logic idx_between_2_6_comb_left;
logic idx_between_2_6_comb_right;
logic idx_between_2_6_comb_out;
logic idx_between_11_15_reg_in;
logic idx_between_11_15_reg_write_en;
logic idx_between_11_15_reg_clk;
logic idx_between_11_15_reg_reset;
logic idx_between_11_15_reg_out;
logic idx_between_11_15_reg_done;
logic idx_between_11_15_comb_left;
logic idx_between_11_15_comb_right;
logic idx_between_11_15_comb_out;
logic idx_between_17_25_reg_in;
logic idx_between_17_25_reg_write_en;
logic idx_between_17_25_reg_clk;
logic idx_between_17_25_reg_reset;
logic idx_between_17_25_reg_out;
logic idx_between_17_25_reg_done;
logic idx_between_17_25_comb_left;
logic idx_between_17_25_comb_right;
logic idx_between_17_25_comb_out;
logic idx_between_13_21_reg_in;
logic idx_between_13_21_reg_write_en;
logic idx_between_13_21_reg_clk;
logic idx_between_13_21_reg_reset;
logic idx_between_13_21_reg_out;
logic idx_between_13_21_reg_done;
logic idx_between_13_21_comb_left;
logic idx_between_13_21_comb_right;
logic idx_between_13_21_comb_out;
logic idx_between_16_17_reg_in;
logic idx_between_16_17_reg_write_en;
logic idx_between_16_17_reg_clk;
logic idx_between_16_17_reg_reset;
logic idx_between_16_17_reg_out;
logic idx_between_16_17_reg_done;
logic idx_between_16_17_comb_left;
logic idx_between_16_17_comb_right;
logic idx_between_16_17_comb_out;
logic cond_in;
logic cond_write_en;
logic cond_clk;
logic cond_reset;
logic cond_out;
logic cond_done;
logic cond_wire_in;
logic cond_wire_out;
logic cond0_in;
logic cond0_write_en;
logic cond0_clk;
logic cond0_reset;
logic cond0_out;
logic cond0_done;
logic cond_wire0_in;
logic cond_wire0_out;
logic cond1_in;
logic cond1_write_en;
logic cond1_clk;
logic cond1_reset;
logic cond1_out;
logic cond1_done;
logic cond_wire1_in;
logic cond_wire1_out;
logic cond2_in;
logic cond2_write_en;
logic cond2_clk;
logic cond2_reset;
logic cond2_out;
logic cond2_done;
logic cond_wire2_in;
logic cond_wire2_out;
logic cond3_in;
logic cond3_write_en;
logic cond3_clk;
logic cond3_reset;
logic cond3_out;
logic cond3_done;
logic cond_wire3_in;
logic cond_wire3_out;
logic cond4_in;
logic cond4_write_en;
logic cond4_clk;
logic cond4_reset;
logic cond4_out;
logic cond4_done;
logic cond_wire4_in;
logic cond_wire4_out;
logic cond5_in;
logic cond5_write_en;
logic cond5_clk;
logic cond5_reset;
logic cond5_out;
logic cond5_done;
logic cond_wire5_in;
logic cond_wire5_out;
logic cond6_in;
logic cond6_write_en;
logic cond6_clk;
logic cond6_reset;
logic cond6_out;
logic cond6_done;
logic cond_wire6_in;
logic cond_wire6_out;
logic cond7_in;
logic cond7_write_en;
logic cond7_clk;
logic cond7_reset;
logic cond7_out;
logic cond7_done;
logic cond_wire7_in;
logic cond_wire7_out;
logic cond8_in;
logic cond8_write_en;
logic cond8_clk;
logic cond8_reset;
logic cond8_out;
logic cond8_done;
logic cond_wire8_in;
logic cond_wire8_out;
logic cond9_in;
logic cond9_write_en;
logic cond9_clk;
logic cond9_reset;
logic cond9_out;
logic cond9_done;
logic cond_wire9_in;
logic cond_wire9_out;
logic cond10_in;
logic cond10_write_en;
logic cond10_clk;
logic cond10_reset;
logic cond10_out;
logic cond10_done;
logic cond_wire10_in;
logic cond_wire10_out;
logic cond11_in;
logic cond11_write_en;
logic cond11_clk;
logic cond11_reset;
logic cond11_out;
logic cond11_done;
logic cond_wire11_in;
logic cond_wire11_out;
logic cond12_in;
logic cond12_write_en;
logic cond12_clk;
logic cond12_reset;
logic cond12_out;
logic cond12_done;
logic cond_wire12_in;
logic cond_wire12_out;
logic cond13_in;
logic cond13_write_en;
logic cond13_clk;
logic cond13_reset;
logic cond13_out;
logic cond13_done;
logic cond_wire13_in;
logic cond_wire13_out;
logic cond14_in;
logic cond14_write_en;
logic cond14_clk;
logic cond14_reset;
logic cond14_out;
logic cond14_done;
logic cond_wire14_in;
logic cond_wire14_out;
logic cond15_in;
logic cond15_write_en;
logic cond15_clk;
logic cond15_reset;
logic cond15_out;
logic cond15_done;
logic cond_wire15_in;
logic cond_wire15_out;
logic cond16_in;
logic cond16_write_en;
logic cond16_clk;
logic cond16_reset;
logic cond16_out;
logic cond16_done;
logic cond_wire16_in;
logic cond_wire16_out;
logic cond17_in;
logic cond17_write_en;
logic cond17_clk;
logic cond17_reset;
logic cond17_out;
logic cond17_done;
logic cond_wire17_in;
logic cond_wire17_out;
logic cond18_in;
logic cond18_write_en;
logic cond18_clk;
logic cond18_reset;
logic cond18_out;
logic cond18_done;
logic cond_wire18_in;
logic cond_wire18_out;
logic cond19_in;
logic cond19_write_en;
logic cond19_clk;
logic cond19_reset;
logic cond19_out;
logic cond19_done;
logic cond_wire19_in;
logic cond_wire19_out;
logic cond20_in;
logic cond20_write_en;
logic cond20_clk;
logic cond20_reset;
logic cond20_out;
logic cond20_done;
logic cond_wire20_in;
logic cond_wire20_out;
logic cond21_in;
logic cond21_write_en;
logic cond21_clk;
logic cond21_reset;
logic cond21_out;
logic cond21_done;
logic cond_wire21_in;
logic cond_wire21_out;
logic cond22_in;
logic cond22_write_en;
logic cond22_clk;
logic cond22_reset;
logic cond22_out;
logic cond22_done;
logic cond_wire22_in;
logic cond_wire22_out;
logic cond23_in;
logic cond23_write_en;
logic cond23_clk;
logic cond23_reset;
logic cond23_out;
logic cond23_done;
logic cond_wire23_in;
logic cond_wire23_out;
logic cond24_in;
logic cond24_write_en;
logic cond24_clk;
logic cond24_reset;
logic cond24_out;
logic cond24_done;
logic cond_wire24_in;
logic cond_wire24_out;
logic cond25_in;
logic cond25_write_en;
logic cond25_clk;
logic cond25_reset;
logic cond25_out;
logic cond25_done;
logic cond_wire25_in;
logic cond_wire25_out;
logic cond26_in;
logic cond26_write_en;
logic cond26_clk;
logic cond26_reset;
logic cond26_out;
logic cond26_done;
logic cond_wire26_in;
logic cond_wire26_out;
logic cond27_in;
logic cond27_write_en;
logic cond27_clk;
logic cond27_reset;
logic cond27_out;
logic cond27_done;
logic cond_wire27_in;
logic cond_wire27_out;
logic cond28_in;
logic cond28_write_en;
logic cond28_clk;
logic cond28_reset;
logic cond28_out;
logic cond28_done;
logic cond_wire28_in;
logic cond_wire28_out;
logic cond29_in;
logic cond29_write_en;
logic cond29_clk;
logic cond29_reset;
logic cond29_out;
logic cond29_done;
logic cond_wire29_in;
logic cond_wire29_out;
logic cond30_in;
logic cond30_write_en;
logic cond30_clk;
logic cond30_reset;
logic cond30_out;
logic cond30_done;
logic cond_wire30_in;
logic cond_wire30_out;
logic cond31_in;
logic cond31_write_en;
logic cond31_clk;
logic cond31_reset;
logic cond31_out;
logic cond31_done;
logic cond_wire31_in;
logic cond_wire31_out;
logic cond32_in;
logic cond32_write_en;
logic cond32_clk;
logic cond32_reset;
logic cond32_out;
logic cond32_done;
logic cond_wire32_in;
logic cond_wire32_out;
logic cond33_in;
logic cond33_write_en;
logic cond33_clk;
logic cond33_reset;
logic cond33_out;
logic cond33_done;
logic cond_wire33_in;
logic cond_wire33_out;
logic cond34_in;
logic cond34_write_en;
logic cond34_clk;
logic cond34_reset;
logic cond34_out;
logic cond34_done;
logic cond_wire34_in;
logic cond_wire34_out;
logic cond35_in;
logic cond35_write_en;
logic cond35_clk;
logic cond35_reset;
logic cond35_out;
logic cond35_done;
logic cond_wire35_in;
logic cond_wire35_out;
logic cond36_in;
logic cond36_write_en;
logic cond36_clk;
logic cond36_reset;
logic cond36_out;
logic cond36_done;
logic cond_wire36_in;
logic cond_wire36_out;
logic cond37_in;
logic cond37_write_en;
logic cond37_clk;
logic cond37_reset;
logic cond37_out;
logic cond37_done;
logic cond_wire37_in;
logic cond_wire37_out;
logic cond38_in;
logic cond38_write_en;
logic cond38_clk;
logic cond38_reset;
logic cond38_out;
logic cond38_done;
logic cond_wire38_in;
logic cond_wire38_out;
logic cond39_in;
logic cond39_write_en;
logic cond39_clk;
logic cond39_reset;
logic cond39_out;
logic cond39_done;
logic cond_wire39_in;
logic cond_wire39_out;
logic cond40_in;
logic cond40_write_en;
logic cond40_clk;
logic cond40_reset;
logic cond40_out;
logic cond40_done;
logic cond_wire40_in;
logic cond_wire40_out;
logic cond41_in;
logic cond41_write_en;
logic cond41_clk;
logic cond41_reset;
logic cond41_out;
logic cond41_done;
logic cond_wire41_in;
logic cond_wire41_out;
logic cond42_in;
logic cond42_write_en;
logic cond42_clk;
logic cond42_reset;
logic cond42_out;
logic cond42_done;
logic cond_wire42_in;
logic cond_wire42_out;
logic cond43_in;
logic cond43_write_en;
logic cond43_clk;
logic cond43_reset;
logic cond43_out;
logic cond43_done;
logic cond_wire43_in;
logic cond_wire43_out;
logic cond44_in;
logic cond44_write_en;
logic cond44_clk;
logic cond44_reset;
logic cond44_out;
logic cond44_done;
logic cond_wire44_in;
logic cond_wire44_out;
logic cond45_in;
logic cond45_write_en;
logic cond45_clk;
logic cond45_reset;
logic cond45_out;
logic cond45_done;
logic cond_wire45_in;
logic cond_wire45_out;
logic cond46_in;
logic cond46_write_en;
logic cond46_clk;
logic cond46_reset;
logic cond46_out;
logic cond46_done;
logic cond_wire46_in;
logic cond_wire46_out;
logic cond47_in;
logic cond47_write_en;
logic cond47_clk;
logic cond47_reset;
logic cond47_out;
logic cond47_done;
logic cond_wire47_in;
logic cond_wire47_out;
logic cond48_in;
logic cond48_write_en;
logic cond48_clk;
logic cond48_reset;
logic cond48_out;
logic cond48_done;
logic cond_wire48_in;
logic cond_wire48_out;
logic cond49_in;
logic cond49_write_en;
logic cond49_clk;
logic cond49_reset;
logic cond49_out;
logic cond49_done;
logic cond_wire49_in;
logic cond_wire49_out;
logic cond50_in;
logic cond50_write_en;
logic cond50_clk;
logic cond50_reset;
logic cond50_out;
logic cond50_done;
logic cond_wire50_in;
logic cond_wire50_out;
logic cond51_in;
logic cond51_write_en;
logic cond51_clk;
logic cond51_reset;
logic cond51_out;
logic cond51_done;
logic cond_wire51_in;
logic cond_wire51_out;
logic cond52_in;
logic cond52_write_en;
logic cond52_clk;
logic cond52_reset;
logic cond52_out;
logic cond52_done;
logic cond_wire52_in;
logic cond_wire52_out;
logic cond53_in;
logic cond53_write_en;
logic cond53_clk;
logic cond53_reset;
logic cond53_out;
logic cond53_done;
logic cond_wire53_in;
logic cond_wire53_out;
logic cond54_in;
logic cond54_write_en;
logic cond54_clk;
logic cond54_reset;
logic cond54_out;
logic cond54_done;
logic cond_wire54_in;
logic cond_wire54_out;
logic cond55_in;
logic cond55_write_en;
logic cond55_clk;
logic cond55_reset;
logic cond55_out;
logic cond55_done;
logic cond_wire55_in;
logic cond_wire55_out;
logic cond56_in;
logic cond56_write_en;
logic cond56_clk;
logic cond56_reset;
logic cond56_out;
logic cond56_done;
logic cond_wire56_in;
logic cond_wire56_out;
logic cond57_in;
logic cond57_write_en;
logic cond57_clk;
logic cond57_reset;
logic cond57_out;
logic cond57_done;
logic cond_wire57_in;
logic cond_wire57_out;
logic cond58_in;
logic cond58_write_en;
logic cond58_clk;
logic cond58_reset;
logic cond58_out;
logic cond58_done;
logic cond_wire58_in;
logic cond_wire58_out;
logic cond59_in;
logic cond59_write_en;
logic cond59_clk;
logic cond59_reset;
logic cond59_out;
logic cond59_done;
logic cond_wire59_in;
logic cond_wire59_out;
logic cond60_in;
logic cond60_write_en;
logic cond60_clk;
logic cond60_reset;
logic cond60_out;
logic cond60_done;
logic cond_wire60_in;
logic cond_wire60_out;
logic cond61_in;
logic cond61_write_en;
logic cond61_clk;
logic cond61_reset;
logic cond61_out;
logic cond61_done;
logic cond_wire61_in;
logic cond_wire61_out;
logic cond62_in;
logic cond62_write_en;
logic cond62_clk;
logic cond62_reset;
logic cond62_out;
logic cond62_done;
logic cond_wire62_in;
logic cond_wire62_out;
logic cond63_in;
logic cond63_write_en;
logic cond63_clk;
logic cond63_reset;
logic cond63_out;
logic cond63_done;
logic cond_wire63_in;
logic cond_wire63_out;
logic cond64_in;
logic cond64_write_en;
logic cond64_clk;
logic cond64_reset;
logic cond64_out;
logic cond64_done;
logic cond_wire64_in;
logic cond_wire64_out;
logic cond65_in;
logic cond65_write_en;
logic cond65_clk;
logic cond65_reset;
logic cond65_out;
logic cond65_done;
logic cond_wire65_in;
logic cond_wire65_out;
logic cond66_in;
logic cond66_write_en;
logic cond66_clk;
logic cond66_reset;
logic cond66_out;
logic cond66_done;
logic cond_wire66_in;
logic cond_wire66_out;
logic cond67_in;
logic cond67_write_en;
logic cond67_clk;
logic cond67_reset;
logic cond67_out;
logic cond67_done;
logic cond_wire67_in;
logic cond_wire67_out;
logic cond68_in;
logic cond68_write_en;
logic cond68_clk;
logic cond68_reset;
logic cond68_out;
logic cond68_done;
logic cond_wire68_in;
logic cond_wire68_out;
logic cond69_in;
logic cond69_write_en;
logic cond69_clk;
logic cond69_reset;
logic cond69_out;
logic cond69_done;
logic cond_wire69_in;
logic cond_wire69_out;
logic cond70_in;
logic cond70_write_en;
logic cond70_clk;
logic cond70_reset;
logic cond70_out;
logic cond70_done;
logic cond_wire70_in;
logic cond_wire70_out;
logic cond71_in;
logic cond71_write_en;
logic cond71_clk;
logic cond71_reset;
logic cond71_out;
logic cond71_done;
logic cond_wire71_in;
logic cond_wire71_out;
logic cond72_in;
logic cond72_write_en;
logic cond72_clk;
logic cond72_reset;
logic cond72_out;
logic cond72_done;
logic cond_wire72_in;
logic cond_wire72_out;
logic cond73_in;
logic cond73_write_en;
logic cond73_clk;
logic cond73_reset;
logic cond73_out;
logic cond73_done;
logic cond_wire73_in;
logic cond_wire73_out;
logic cond74_in;
logic cond74_write_en;
logic cond74_clk;
logic cond74_reset;
logic cond74_out;
logic cond74_done;
logic cond_wire74_in;
logic cond_wire74_out;
logic cond75_in;
logic cond75_write_en;
logic cond75_clk;
logic cond75_reset;
logic cond75_out;
logic cond75_done;
logic cond_wire75_in;
logic cond_wire75_out;
logic cond76_in;
logic cond76_write_en;
logic cond76_clk;
logic cond76_reset;
logic cond76_out;
logic cond76_done;
logic cond_wire76_in;
logic cond_wire76_out;
logic cond77_in;
logic cond77_write_en;
logic cond77_clk;
logic cond77_reset;
logic cond77_out;
logic cond77_done;
logic cond_wire77_in;
logic cond_wire77_out;
logic cond78_in;
logic cond78_write_en;
logic cond78_clk;
logic cond78_reset;
logic cond78_out;
logic cond78_done;
logic cond_wire78_in;
logic cond_wire78_out;
logic cond79_in;
logic cond79_write_en;
logic cond79_clk;
logic cond79_reset;
logic cond79_out;
logic cond79_done;
logic cond_wire79_in;
logic cond_wire79_out;
logic cond80_in;
logic cond80_write_en;
logic cond80_clk;
logic cond80_reset;
logic cond80_out;
logic cond80_done;
logic cond_wire80_in;
logic cond_wire80_out;
logic cond81_in;
logic cond81_write_en;
logic cond81_clk;
logic cond81_reset;
logic cond81_out;
logic cond81_done;
logic cond_wire81_in;
logic cond_wire81_out;
logic cond82_in;
logic cond82_write_en;
logic cond82_clk;
logic cond82_reset;
logic cond82_out;
logic cond82_done;
logic cond_wire82_in;
logic cond_wire82_out;
logic cond83_in;
logic cond83_write_en;
logic cond83_clk;
logic cond83_reset;
logic cond83_out;
logic cond83_done;
logic cond_wire83_in;
logic cond_wire83_out;
logic cond84_in;
logic cond84_write_en;
logic cond84_clk;
logic cond84_reset;
logic cond84_out;
logic cond84_done;
logic cond_wire84_in;
logic cond_wire84_out;
logic cond85_in;
logic cond85_write_en;
logic cond85_clk;
logic cond85_reset;
logic cond85_out;
logic cond85_done;
logic cond_wire85_in;
logic cond_wire85_out;
logic cond86_in;
logic cond86_write_en;
logic cond86_clk;
logic cond86_reset;
logic cond86_out;
logic cond86_done;
logic cond_wire86_in;
logic cond_wire86_out;
logic cond87_in;
logic cond87_write_en;
logic cond87_clk;
logic cond87_reset;
logic cond87_out;
logic cond87_done;
logic cond_wire87_in;
logic cond_wire87_out;
logic cond88_in;
logic cond88_write_en;
logic cond88_clk;
logic cond88_reset;
logic cond88_out;
logic cond88_done;
logic cond_wire88_in;
logic cond_wire88_out;
logic cond89_in;
logic cond89_write_en;
logic cond89_clk;
logic cond89_reset;
logic cond89_out;
logic cond89_done;
logic cond_wire89_in;
logic cond_wire89_out;
logic cond90_in;
logic cond90_write_en;
logic cond90_clk;
logic cond90_reset;
logic cond90_out;
logic cond90_done;
logic cond_wire90_in;
logic cond_wire90_out;
logic cond91_in;
logic cond91_write_en;
logic cond91_clk;
logic cond91_reset;
logic cond91_out;
logic cond91_done;
logic cond_wire91_in;
logic cond_wire91_out;
logic cond92_in;
logic cond92_write_en;
logic cond92_clk;
logic cond92_reset;
logic cond92_out;
logic cond92_done;
logic cond_wire92_in;
logic cond_wire92_out;
logic cond93_in;
logic cond93_write_en;
logic cond93_clk;
logic cond93_reset;
logic cond93_out;
logic cond93_done;
logic cond_wire93_in;
logic cond_wire93_out;
logic cond94_in;
logic cond94_write_en;
logic cond94_clk;
logic cond94_reset;
logic cond94_out;
logic cond94_done;
logic cond_wire94_in;
logic cond_wire94_out;
logic cond95_in;
logic cond95_write_en;
logic cond95_clk;
logic cond95_reset;
logic cond95_out;
logic cond95_done;
logic cond_wire95_in;
logic cond_wire95_out;
logic cond96_in;
logic cond96_write_en;
logic cond96_clk;
logic cond96_reset;
logic cond96_out;
logic cond96_done;
logic cond_wire96_in;
logic cond_wire96_out;
logic cond97_in;
logic cond97_write_en;
logic cond97_clk;
logic cond97_reset;
logic cond97_out;
logic cond97_done;
logic cond_wire97_in;
logic cond_wire97_out;
logic cond98_in;
logic cond98_write_en;
logic cond98_clk;
logic cond98_reset;
logic cond98_out;
logic cond98_done;
logic cond_wire98_in;
logic cond_wire98_out;
logic cond99_in;
logic cond99_write_en;
logic cond99_clk;
logic cond99_reset;
logic cond99_out;
logic cond99_done;
logic cond_wire99_in;
logic cond_wire99_out;
logic cond100_in;
logic cond100_write_en;
logic cond100_clk;
logic cond100_reset;
logic cond100_out;
logic cond100_done;
logic cond_wire100_in;
logic cond_wire100_out;
logic cond101_in;
logic cond101_write_en;
logic cond101_clk;
logic cond101_reset;
logic cond101_out;
logic cond101_done;
logic cond_wire101_in;
logic cond_wire101_out;
logic cond102_in;
logic cond102_write_en;
logic cond102_clk;
logic cond102_reset;
logic cond102_out;
logic cond102_done;
logic cond_wire102_in;
logic cond_wire102_out;
logic cond103_in;
logic cond103_write_en;
logic cond103_clk;
logic cond103_reset;
logic cond103_out;
logic cond103_done;
logic cond_wire103_in;
logic cond_wire103_out;
logic cond104_in;
logic cond104_write_en;
logic cond104_clk;
logic cond104_reset;
logic cond104_out;
logic cond104_done;
logic cond_wire104_in;
logic cond_wire104_out;
logic cond105_in;
logic cond105_write_en;
logic cond105_clk;
logic cond105_reset;
logic cond105_out;
logic cond105_done;
logic cond_wire105_in;
logic cond_wire105_out;
logic cond106_in;
logic cond106_write_en;
logic cond106_clk;
logic cond106_reset;
logic cond106_out;
logic cond106_done;
logic cond_wire106_in;
logic cond_wire106_out;
logic cond107_in;
logic cond107_write_en;
logic cond107_clk;
logic cond107_reset;
logic cond107_out;
logic cond107_done;
logic cond_wire107_in;
logic cond_wire107_out;
logic cond108_in;
logic cond108_write_en;
logic cond108_clk;
logic cond108_reset;
logic cond108_out;
logic cond108_done;
logic cond_wire108_in;
logic cond_wire108_out;
logic cond109_in;
logic cond109_write_en;
logic cond109_clk;
logic cond109_reset;
logic cond109_out;
logic cond109_done;
logic cond_wire109_in;
logic cond_wire109_out;
logic cond110_in;
logic cond110_write_en;
logic cond110_clk;
logic cond110_reset;
logic cond110_out;
logic cond110_done;
logic cond_wire110_in;
logic cond_wire110_out;
logic cond111_in;
logic cond111_write_en;
logic cond111_clk;
logic cond111_reset;
logic cond111_out;
logic cond111_done;
logic cond_wire111_in;
logic cond_wire111_out;
logic cond112_in;
logic cond112_write_en;
logic cond112_clk;
logic cond112_reset;
logic cond112_out;
logic cond112_done;
logic cond_wire112_in;
logic cond_wire112_out;
logic cond113_in;
logic cond113_write_en;
logic cond113_clk;
logic cond113_reset;
logic cond113_out;
logic cond113_done;
logic cond_wire113_in;
logic cond_wire113_out;
logic cond114_in;
logic cond114_write_en;
logic cond114_clk;
logic cond114_reset;
logic cond114_out;
logic cond114_done;
logic cond_wire114_in;
logic cond_wire114_out;
logic cond115_in;
logic cond115_write_en;
logic cond115_clk;
logic cond115_reset;
logic cond115_out;
logic cond115_done;
logic cond_wire115_in;
logic cond_wire115_out;
logic cond116_in;
logic cond116_write_en;
logic cond116_clk;
logic cond116_reset;
logic cond116_out;
logic cond116_done;
logic cond_wire116_in;
logic cond_wire116_out;
logic cond117_in;
logic cond117_write_en;
logic cond117_clk;
logic cond117_reset;
logic cond117_out;
logic cond117_done;
logic cond_wire117_in;
logic cond_wire117_out;
logic cond118_in;
logic cond118_write_en;
logic cond118_clk;
logic cond118_reset;
logic cond118_out;
logic cond118_done;
logic cond_wire118_in;
logic cond_wire118_out;
logic cond119_in;
logic cond119_write_en;
logic cond119_clk;
logic cond119_reset;
logic cond119_out;
logic cond119_done;
logic cond_wire119_in;
logic cond_wire119_out;
logic cond120_in;
logic cond120_write_en;
logic cond120_clk;
logic cond120_reset;
logic cond120_out;
logic cond120_done;
logic cond_wire120_in;
logic cond_wire120_out;
logic cond121_in;
logic cond121_write_en;
logic cond121_clk;
logic cond121_reset;
logic cond121_out;
logic cond121_done;
logic cond_wire121_in;
logic cond_wire121_out;
logic cond122_in;
logic cond122_write_en;
logic cond122_clk;
logic cond122_reset;
logic cond122_out;
logic cond122_done;
logic cond_wire122_in;
logic cond_wire122_out;
logic cond123_in;
logic cond123_write_en;
logic cond123_clk;
logic cond123_reset;
logic cond123_out;
logic cond123_done;
logic cond_wire123_in;
logic cond_wire123_out;
logic cond124_in;
logic cond124_write_en;
logic cond124_clk;
logic cond124_reset;
logic cond124_out;
logic cond124_done;
logic cond_wire124_in;
logic cond_wire124_out;
logic cond125_in;
logic cond125_write_en;
logic cond125_clk;
logic cond125_reset;
logic cond125_out;
logic cond125_done;
logic cond_wire125_in;
logic cond_wire125_out;
logic cond126_in;
logic cond126_write_en;
logic cond126_clk;
logic cond126_reset;
logic cond126_out;
logic cond126_done;
logic cond_wire126_in;
logic cond_wire126_out;
logic cond127_in;
logic cond127_write_en;
logic cond127_clk;
logic cond127_reset;
logic cond127_out;
logic cond127_done;
logic cond_wire127_in;
logic cond_wire127_out;
logic cond128_in;
logic cond128_write_en;
logic cond128_clk;
logic cond128_reset;
logic cond128_out;
logic cond128_done;
logic cond_wire128_in;
logic cond_wire128_out;
logic cond129_in;
logic cond129_write_en;
logic cond129_clk;
logic cond129_reset;
logic cond129_out;
logic cond129_done;
logic cond_wire129_in;
logic cond_wire129_out;
logic cond130_in;
logic cond130_write_en;
logic cond130_clk;
logic cond130_reset;
logic cond130_out;
logic cond130_done;
logic cond_wire130_in;
logic cond_wire130_out;
logic cond131_in;
logic cond131_write_en;
logic cond131_clk;
logic cond131_reset;
logic cond131_out;
logic cond131_done;
logic cond_wire131_in;
logic cond_wire131_out;
logic cond132_in;
logic cond132_write_en;
logic cond132_clk;
logic cond132_reset;
logic cond132_out;
logic cond132_done;
logic cond_wire132_in;
logic cond_wire132_out;
logic cond133_in;
logic cond133_write_en;
logic cond133_clk;
logic cond133_reset;
logic cond133_out;
logic cond133_done;
logic cond_wire133_in;
logic cond_wire133_out;
logic cond134_in;
logic cond134_write_en;
logic cond134_clk;
logic cond134_reset;
logic cond134_out;
logic cond134_done;
logic cond_wire134_in;
logic cond_wire134_out;
logic cond135_in;
logic cond135_write_en;
logic cond135_clk;
logic cond135_reset;
logic cond135_out;
logic cond135_done;
logic cond_wire135_in;
logic cond_wire135_out;
logic cond136_in;
logic cond136_write_en;
logic cond136_clk;
logic cond136_reset;
logic cond136_out;
logic cond136_done;
logic cond_wire136_in;
logic cond_wire136_out;
logic cond137_in;
logic cond137_write_en;
logic cond137_clk;
logic cond137_reset;
logic cond137_out;
logic cond137_done;
logic cond_wire137_in;
logic cond_wire137_out;
logic cond138_in;
logic cond138_write_en;
logic cond138_clk;
logic cond138_reset;
logic cond138_out;
logic cond138_done;
logic cond_wire138_in;
logic cond_wire138_out;
logic cond139_in;
logic cond139_write_en;
logic cond139_clk;
logic cond139_reset;
logic cond139_out;
logic cond139_done;
logic cond_wire139_in;
logic cond_wire139_out;
logic cond140_in;
logic cond140_write_en;
logic cond140_clk;
logic cond140_reset;
logic cond140_out;
logic cond140_done;
logic cond_wire140_in;
logic cond_wire140_out;
logic cond141_in;
logic cond141_write_en;
logic cond141_clk;
logic cond141_reset;
logic cond141_out;
logic cond141_done;
logic cond_wire141_in;
logic cond_wire141_out;
logic cond142_in;
logic cond142_write_en;
logic cond142_clk;
logic cond142_reset;
logic cond142_out;
logic cond142_done;
logic cond_wire142_in;
logic cond_wire142_out;
logic cond143_in;
logic cond143_write_en;
logic cond143_clk;
logic cond143_reset;
logic cond143_out;
logic cond143_done;
logic cond_wire143_in;
logic cond_wire143_out;
logic cond144_in;
logic cond144_write_en;
logic cond144_clk;
logic cond144_reset;
logic cond144_out;
logic cond144_done;
logic cond_wire144_in;
logic cond_wire144_out;
logic cond145_in;
logic cond145_write_en;
logic cond145_clk;
logic cond145_reset;
logic cond145_out;
logic cond145_done;
logic cond_wire145_in;
logic cond_wire145_out;
logic cond146_in;
logic cond146_write_en;
logic cond146_clk;
logic cond146_reset;
logic cond146_out;
logic cond146_done;
logic cond_wire146_in;
logic cond_wire146_out;
logic cond147_in;
logic cond147_write_en;
logic cond147_clk;
logic cond147_reset;
logic cond147_out;
logic cond147_done;
logic cond_wire147_in;
logic cond_wire147_out;
logic cond148_in;
logic cond148_write_en;
logic cond148_clk;
logic cond148_reset;
logic cond148_out;
logic cond148_done;
logic cond_wire148_in;
logic cond_wire148_out;
logic cond149_in;
logic cond149_write_en;
logic cond149_clk;
logic cond149_reset;
logic cond149_out;
logic cond149_done;
logic cond_wire149_in;
logic cond_wire149_out;
logic cond150_in;
logic cond150_write_en;
logic cond150_clk;
logic cond150_reset;
logic cond150_out;
logic cond150_done;
logic cond_wire150_in;
logic cond_wire150_out;
logic cond151_in;
logic cond151_write_en;
logic cond151_clk;
logic cond151_reset;
logic cond151_out;
logic cond151_done;
logic cond_wire151_in;
logic cond_wire151_out;
logic cond152_in;
logic cond152_write_en;
logic cond152_clk;
logic cond152_reset;
logic cond152_out;
logic cond152_done;
logic cond_wire152_in;
logic cond_wire152_out;
logic cond153_in;
logic cond153_write_en;
logic cond153_clk;
logic cond153_reset;
logic cond153_out;
logic cond153_done;
logic cond_wire153_in;
logic cond_wire153_out;
logic cond154_in;
logic cond154_write_en;
logic cond154_clk;
logic cond154_reset;
logic cond154_out;
logic cond154_done;
logic cond_wire154_in;
logic cond_wire154_out;
logic cond155_in;
logic cond155_write_en;
logic cond155_clk;
logic cond155_reset;
logic cond155_out;
logic cond155_done;
logic cond_wire155_in;
logic cond_wire155_out;
logic cond156_in;
logic cond156_write_en;
logic cond156_clk;
logic cond156_reset;
logic cond156_out;
logic cond156_done;
logic cond_wire156_in;
logic cond_wire156_out;
logic cond157_in;
logic cond157_write_en;
logic cond157_clk;
logic cond157_reset;
logic cond157_out;
logic cond157_done;
logic cond_wire157_in;
logic cond_wire157_out;
logic cond158_in;
logic cond158_write_en;
logic cond158_clk;
logic cond158_reset;
logic cond158_out;
logic cond158_done;
logic cond_wire158_in;
logic cond_wire158_out;
logic cond159_in;
logic cond159_write_en;
logic cond159_clk;
logic cond159_reset;
logic cond159_out;
logic cond159_done;
logic cond_wire159_in;
logic cond_wire159_out;
logic cond160_in;
logic cond160_write_en;
logic cond160_clk;
logic cond160_reset;
logic cond160_out;
logic cond160_done;
logic cond_wire160_in;
logic cond_wire160_out;
logic cond161_in;
logic cond161_write_en;
logic cond161_clk;
logic cond161_reset;
logic cond161_out;
logic cond161_done;
logic cond_wire161_in;
logic cond_wire161_out;
logic cond162_in;
logic cond162_write_en;
logic cond162_clk;
logic cond162_reset;
logic cond162_out;
logic cond162_done;
logic cond_wire162_in;
logic cond_wire162_out;
logic cond163_in;
logic cond163_write_en;
logic cond163_clk;
logic cond163_reset;
logic cond163_out;
logic cond163_done;
logic cond_wire163_in;
logic cond_wire163_out;
logic cond164_in;
logic cond164_write_en;
logic cond164_clk;
logic cond164_reset;
logic cond164_out;
logic cond164_done;
logic cond_wire164_in;
logic cond_wire164_out;
logic cond165_in;
logic cond165_write_en;
logic cond165_clk;
logic cond165_reset;
logic cond165_out;
logic cond165_done;
logic cond_wire165_in;
logic cond_wire165_out;
logic cond166_in;
logic cond166_write_en;
logic cond166_clk;
logic cond166_reset;
logic cond166_out;
logic cond166_done;
logic cond_wire166_in;
logic cond_wire166_out;
logic cond167_in;
logic cond167_write_en;
logic cond167_clk;
logic cond167_reset;
logic cond167_out;
logic cond167_done;
logic cond_wire167_in;
logic cond_wire167_out;
logic cond168_in;
logic cond168_write_en;
logic cond168_clk;
logic cond168_reset;
logic cond168_out;
logic cond168_done;
logic cond_wire168_in;
logic cond_wire168_out;
logic cond169_in;
logic cond169_write_en;
logic cond169_clk;
logic cond169_reset;
logic cond169_out;
logic cond169_done;
logic cond_wire169_in;
logic cond_wire169_out;
logic cond170_in;
logic cond170_write_en;
logic cond170_clk;
logic cond170_reset;
logic cond170_out;
logic cond170_done;
logic cond_wire170_in;
logic cond_wire170_out;
logic cond171_in;
logic cond171_write_en;
logic cond171_clk;
logic cond171_reset;
logic cond171_out;
logic cond171_done;
logic cond_wire171_in;
logic cond_wire171_out;
logic cond172_in;
logic cond172_write_en;
logic cond172_clk;
logic cond172_reset;
logic cond172_out;
logic cond172_done;
logic cond_wire172_in;
logic cond_wire172_out;
logic cond173_in;
logic cond173_write_en;
logic cond173_clk;
logic cond173_reset;
logic cond173_out;
logic cond173_done;
logic cond_wire173_in;
logic cond_wire173_out;
logic cond174_in;
logic cond174_write_en;
logic cond174_clk;
logic cond174_reset;
logic cond174_out;
logic cond174_done;
logic cond_wire174_in;
logic cond_wire174_out;
logic cond175_in;
logic cond175_write_en;
logic cond175_clk;
logic cond175_reset;
logic cond175_out;
logic cond175_done;
logic cond_wire175_in;
logic cond_wire175_out;
logic cond176_in;
logic cond176_write_en;
logic cond176_clk;
logic cond176_reset;
logic cond176_out;
logic cond176_done;
logic cond_wire176_in;
logic cond_wire176_out;
logic cond177_in;
logic cond177_write_en;
logic cond177_clk;
logic cond177_reset;
logic cond177_out;
logic cond177_done;
logic cond_wire177_in;
logic cond_wire177_out;
logic cond178_in;
logic cond178_write_en;
logic cond178_clk;
logic cond178_reset;
logic cond178_out;
logic cond178_done;
logic cond_wire178_in;
logic cond_wire178_out;
logic cond179_in;
logic cond179_write_en;
logic cond179_clk;
logic cond179_reset;
logic cond179_out;
logic cond179_done;
logic cond_wire179_in;
logic cond_wire179_out;
logic cond180_in;
logic cond180_write_en;
logic cond180_clk;
logic cond180_reset;
logic cond180_out;
logic cond180_done;
logic cond_wire180_in;
logic cond_wire180_out;
logic cond181_in;
logic cond181_write_en;
logic cond181_clk;
logic cond181_reset;
logic cond181_out;
logic cond181_done;
logic cond_wire181_in;
logic cond_wire181_out;
logic cond182_in;
logic cond182_write_en;
logic cond182_clk;
logic cond182_reset;
logic cond182_out;
logic cond182_done;
logic cond_wire182_in;
logic cond_wire182_out;
logic cond183_in;
logic cond183_write_en;
logic cond183_clk;
logic cond183_reset;
logic cond183_out;
logic cond183_done;
logic cond_wire183_in;
logic cond_wire183_out;
logic cond184_in;
logic cond184_write_en;
logic cond184_clk;
logic cond184_reset;
logic cond184_out;
logic cond184_done;
logic cond_wire184_in;
logic cond_wire184_out;
logic cond185_in;
logic cond185_write_en;
logic cond185_clk;
logic cond185_reset;
logic cond185_out;
logic cond185_done;
logic cond_wire185_in;
logic cond_wire185_out;
logic cond186_in;
logic cond186_write_en;
logic cond186_clk;
logic cond186_reset;
logic cond186_out;
logic cond186_done;
logic cond_wire186_in;
logic cond_wire186_out;
logic cond187_in;
logic cond187_write_en;
logic cond187_clk;
logic cond187_reset;
logic cond187_out;
logic cond187_done;
logic cond_wire187_in;
logic cond_wire187_out;
logic cond188_in;
logic cond188_write_en;
logic cond188_clk;
logic cond188_reset;
logic cond188_out;
logic cond188_done;
logic cond_wire188_in;
logic cond_wire188_out;
logic cond189_in;
logic cond189_write_en;
logic cond189_clk;
logic cond189_reset;
logic cond189_out;
logic cond189_done;
logic cond_wire189_in;
logic cond_wire189_out;
logic cond190_in;
logic cond190_write_en;
logic cond190_clk;
logic cond190_reset;
logic cond190_out;
logic cond190_done;
logic cond_wire190_in;
logic cond_wire190_out;
logic cond191_in;
logic cond191_write_en;
logic cond191_clk;
logic cond191_reset;
logic cond191_out;
logic cond191_done;
logic cond_wire191_in;
logic cond_wire191_out;
logic cond192_in;
logic cond192_write_en;
logic cond192_clk;
logic cond192_reset;
logic cond192_out;
logic cond192_done;
logic cond_wire192_in;
logic cond_wire192_out;
logic cond193_in;
logic cond193_write_en;
logic cond193_clk;
logic cond193_reset;
logic cond193_out;
logic cond193_done;
logic cond_wire193_in;
logic cond_wire193_out;
logic cond194_in;
logic cond194_write_en;
logic cond194_clk;
logic cond194_reset;
logic cond194_out;
logic cond194_done;
logic cond_wire194_in;
logic cond_wire194_out;
logic cond195_in;
logic cond195_write_en;
logic cond195_clk;
logic cond195_reset;
logic cond195_out;
logic cond195_done;
logic cond_wire195_in;
logic cond_wire195_out;
logic cond196_in;
logic cond196_write_en;
logic cond196_clk;
logic cond196_reset;
logic cond196_out;
logic cond196_done;
logic cond_wire196_in;
logic cond_wire196_out;
logic cond197_in;
logic cond197_write_en;
logic cond197_clk;
logic cond197_reset;
logic cond197_out;
logic cond197_done;
logic cond_wire197_in;
logic cond_wire197_out;
logic cond198_in;
logic cond198_write_en;
logic cond198_clk;
logic cond198_reset;
logic cond198_out;
logic cond198_done;
logic cond_wire198_in;
logic cond_wire198_out;
logic cond199_in;
logic cond199_write_en;
logic cond199_clk;
logic cond199_reset;
logic cond199_out;
logic cond199_done;
logic cond_wire199_in;
logic cond_wire199_out;
logic cond200_in;
logic cond200_write_en;
logic cond200_clk;
logic cond200_reset;
logic cond200_out;
logic cond200_done;
logic cond_wire200_in;
logic cond_wire200_out;
logic cond201_in;
logic cond201_write_en;
logic cond201_clk;
logic cond201_reset;
logic cond201_out;
logic cond201_done;
logic cond_wire201_in;
logic cond_wire201_out;
logic cond202_in;
logic cond202_write_en;
logic cond202_clk;
logic cond202_reset;
logic cond202_out;
logic cond202_done;
logic cond_wire202_in;
logic cond_wire202_out;
logic cond203_in;
logic cond203_write_en;
logic cond203_clk;
logic cond203_reset;
logic cond203_out;
logic cond203_done;
logic cond_wire203_in;
logic cond_wire203_out;
logic cond204_in;
logic cond204_write_en;
logic cond204_clk;
logic cond204_reset;
logic cond204_out;
logic cond204_done;
logic cond_wire204_in;
logic cond_wire204_out;
logic cond205_in;
logic cond205_write_en;
logic cond205_clk;
logic cond205_reset;
logic cond205_out;
logic cond205_done;
logic cond_wire205_in;
logic cond_wire205_out;
logic cond206_in;
logic cond206_write_en;
logic cond206_clk;
logic cond206_reset;
logic cond206_out;
logic cond206_done;
logic cond_wire206_in;
logic cond_wire206_out;
logic cond207_in;
logic cond207_write_en;
logic cond207_clk;
logic cond207_reset;
logic cond207_out;
logic cond207_done;
logic cond_wire207_in;
logic cond_wire207_out;
logic cond208_in;
logic cond208_write_en;
logic cond208_clk;
logic cond208_reset;
logic cond208_out;
logic cond208_done;
logic cond_wire208_in;
logic cond_wire208_out;
logic cond209_in;
logic cond209_write_en;
logic cond209_clk;
logic cond209_reset;
logic cond209_out;
logic cond209_done;
logic cond_wire209_in;
logic cond_wire209_out;
logic cond210_in;
logic cond210_write_en;
logic cond210_clk;
logic cond210_reset;
logic cond210_out;
logic cond210_done;
logic cond_wire210_in;
logic cond_wire210_out;
logic cond211_in;
logic cond211_write_en;
logic cond211_clk;
logic cond211_reset;
logic cond211_out;
logic cond211_done;
logic cond_wire211_in;
logic cond_wire211_out;
logic cond212_in;
logic cond212_write_en;
logic cond212_clk;
logic cond212_reset;
logic cond212_out;
logic cond212_done;
logic cond_wire212_in;
logic cond_wire212_out;
logic cond213_in;
logic cond213_write_en;
logic cond213_clk;
logic cond213_reset;
logic cond213_out;
logic cond213_done;
logic cond_wire213_in;
logic cond_wire213_out;
logic cond214_in;
logic cond214_write_en;
logic cond214_clk;
logic cond214_reset;
logic cond214_out;
logic cond214_done;
logic cond_wire214_in;
logic cond_wire214_out;
logic cond215_in;
logic cond215_write_en;
logic cond215_clk;
logic cond215_reset;
logic cond215_out;
logic cond215_done;
logic cond_wire215_in;
logic cond_wire215_out;
logic cond216_in;
logic cond216_write_en;
logic cond216_clk;
logic cond216_reset;
logic cond216_out;
logic cond216_done;
logic cond_wire216_in;
logic cond_wire216_out;
logic cond217_in;
logic cond217_write_en;
logic cond217_clk;
logic cond217_reset;
logic cond217_out;
logic cond217_done;
logic cond_wire217_in;
logic cond_wire217_out;
logic cond218_in;
logic cond218_write_en;
logic cond218_clk;
logic cond218_reset;
logic cond218_out;
logic cond218_done;
logic cond_wire218_in;
logic cond_wire218_out;
logic cond219_in;
logic cond219_write_en;
logic cond219_clk;
logic cond219_reset;
logic cond219_out;
logic cond219_done;
logic cond_wire219_in;
logic cond_wire219_out;
logic cond220_in;
logic cond220_write_en;
logic cond220_clk;
logic cond220_reset;
logic cond220_out;
logic cond220_done;
logic cond_wire220_in;
logic cond_wire220_out;
logic cond221_in;
logic cond221_write_en;
logic cond221_clk;
logic cond221_reset;
logic cond221_out;
logic cond221_done;
logic cond_wire221_in;
logic cond_wire221_out;
logic cond222_in;
logic cond222_write_en;
logic cond222_clk;
logic cond222_reset;
logic cond222_out;
logic cond222_done;
logic cond_wire222_in;
logic cond_wire222_out;
logic cond223_in;
logic cond223_write_en;
logic cond223_clk;
logic cond223_reset;
logic cond223_out;
logic cond223_done;
logic cond_wire223_in;
logic cond_wire223_out;
logic cond224_in;
logic cond224_write_en;
logic cond224_clk;
logic cond224_reset;
logic cond224_out;
logic cond224_done;
logic cond_wire224_in;
logic cond_wire224_out;
logic cond225_in;
logic cond225_write_en;
logic cond225_clk;
logic cond225_reset;
logic cond225_out;
logic cond225_done;
logic cond_wire225_in;
logic cond_wire225_out;
logic cond226_in;
logic cond226_write_en;
logic cond226_clk;
logic cond226_reset;
logic cond226_out;
logic cond226_done;
logic cond_wire226_in;
logic cond_wire226_out;
logic cond227_in;
logic cond227_write_en;
logic cond227_clk;
logic cond227_reset;
logic cond227_out;
logic cond227_done;
logic cond_wire227_in;
logic cond_wire227_out;
logic cond228_in;
logic cond228_write_en;
logic cond228_clk;
logic cond228_reset;
logic cond228_out;
logic cond228_done;
logic cond_wire228_in;
logic cond_wire228_out;
logic cond229_in;
logic cond229_write_en;
logic cond229_clk;
logic cond229_reset;
logic cond229_out;
logic cond229_done;
logic cond_wire229_in;
logic cond_wire229_out;
logic cond230_in;
logic cond230_write_en;
logic cond230_clk;
logic cond230_reset;
logic cond230_out;
logic cond230_done;
logic cond_wire230_in;
logic cond_wire230_out;
logic cond231_in;
logic cond231_write_en;
logic cond231_clk;
logic cond231_reset;
logic cond231_out;
logic cond231_done;
logic cond_wire231_in;
logic cond_wire231_out;
logic cond232_in;
logic cond232_write_en;
logic cond232_clk;
logic cond232_reset;
logic cond232_out;
logic cond232_done;
logic cond_wire232_in;
logic cond_wire232_out;
logic cond233_in;
logic cond233_write_en;
logic cond233_clk;
logic cond233_reset;
logic cond233_out;
logic cond233_done;
logic cond_wire233_in;
logic cond_wire233_out;
logic cond234_in;
logic cond234_write_en;
logic cond234_clk;
logic cond234_reset;
logic cond234_out;
logic cond234_done;
logic cond_wire234_in;
logic cond_wire234_out;
logic cond235_in;
logic cond235_write_en;
logic cond235_clk;
logic cond235_reset;
logic cond235_out;
logic cond235_done;
logic cond_wire235_in;
logic cond_wire235_out;
logic cond236_in;
logic cond236_write_en;
logic cond236_clk;
logic cond236_reset;
logic cond236_out;
logic cond236_done;
logic cond_wire236_in;
logic cond_wire236_out;
logic cond237_in;
logic cond237_write_en;
logic cond237_clk;
logic cond237_reset;
logic cond237_out;
logic cond237_done;
logic cond_wire237_in;
logic cond_wire237_out;
logic cond238_in;
logic cond238_write_en;
logic cond238_clk;
logic cond238_reset;
logic cond238_out;
logic cond238_done;
logic cond_wire238_in;
logic cond_wire238_out;
logic cond239_in;
logic cond239_write_en;
logic cond239_clk;
logic cond239_reset;
logic cond239_out;
logic cond239_done;
logic cond_wire239_in;
logic cond_wire239_out;
logic cond240_in;
logic cond240_write_en;
logic cond240_clk;
logic cond240_reset;
logic cond240_out;
logic cond240_done;
logic cond_wire240_in;
logic cond_wire240_out;
logic cond241_in;
logic cond241_write_en;
logic cond241_clk;
logic cond241_reset;
logic cond241_out;
logic cond241_done;
logic cond_wire241_in;
logic cond_wire241_out;
logic cond242_in;
logic cond242_write_en;
logic cond242_clk;
logic cond242_reset;
logic cond242_out;
logic cond242_done;
logic cond_wire242_in;
logic cond_wire242_out;
logic cond243_in;
logic cond243_write_en;
logic cond243_clk;
logic cond243_reset;
logic cond243_out;
logic cond243_done;
logic cond_wire243_in;
logic cond_wire243_out;
logic cond244_in;
logic cond244_write_en;
logic cond244_clk;
logic cond244_reset;
logic cond244_out;
logic cond244_done;
logic cond_wire244_in;
logic cond_wire244_out;
logic cond245_in;
logic cond245_write_en;
logic cond245_clk;
logic cond245_reset;
logic cond245_out;
logic cond245_done;
logic cond_wire245_in;
logic cond_wire245_out;
logic cond246_in;
logic cond246_write_en;
logic cond246_clk;
logic cond246_reset;
logic cond246_out;
logic cond246_done;
logic cond_wire246_in;
logic cond_wire246_out;
logic cond247_in;
logic cond247_write_en;
logic cond247_clk;
logic cond247_reset;
logic cond247_out;
logic cond247_done;
logic cond_wire247_in;
logic cond_wire247_out;
logic cond248_in;
logic cond248_write_en;
logic cond248_clk;
logic cond248_reset;
logic cond248_out;
logic cond248_done;
logic cond_wire248_in;
logic cond_wire248_out;
logic cond249_in;
logic cond249_write_en;
logic cond249_clk;
logic cond249_reset;
logic cond249_out;
logic cond249_done;
logic cond_wire249_in;
logic cond_wire249_out;
logic cond250_in;
logic cond250_write_en;
logic cond250_clk;
logic cond250_reset;
logic cond250_out;
logic cond250_done;
logic cond_wire250_in;
logic cond_wire250_out;
logic cond251_in;
logic cond251_write_en;
logic cond251_clk;
logic cond251_reset;
logic cond251_out;
logic cond251_done;
logic cond_wire251_in;
logic cond_wire251_out;
logic cond252_in;
logic cond252_write_en;
logic cond252_clk;
logic cond252_reset;
logic cond252_out;
logic cond252_done;
logic cond_wire252_in;
logic cond_wire252_out;
logic cond253_in;
logic cond253_write_en;
logic cond253_clk;
logic cond253_reset;
logic cond253_out;
logic cond253_done;
logic cond_wire253_in;
logic cond_wire253_out;
logic cond254_in;
logic cond254_write_en;
logic cond254_clk;
logic cond254_reset;
logic cond254_out;
logic cond254_done;
logic cond_wire254_in;
logic cond_wire254_out;
logic cond255_in;
logic cond255_write_en;
logic cond255_clk;
logic cond255_reset;
logic cond255_out;
logic cond255_done;
logic cond_wire255_in;
logic cond_wire255_out;
logic cond256_in;
logic cond256_write_en;
logic cond256_clk;
logic cond256_reset;
logic cond256_out;
logic cond256_done;
logic cond_wire256_in;
logic cond_wire256_out;
logic cond257_in;
logic cond257_write_en;
logic cond257_clk;
logic cond257_reset;
logic cond257_out;
logic cond257_done;
logic cond_wire257_in;
logic cond_wire257_out;
logic cond258_in;
logic cond258_write_en;
logic cond258_clk;
logic cond258_reset;
logic cond258_out;
logic cond258_done;
logic cond_wire258_in;
logic cond_wire258_out;
logic cond259_in;
logic cond259_write_en;
logic cond259_clk;
logic cond259_reset;
logic cond259_out;
logic cond259_done;
logic cond_wire259_in;
logic cond_wire259_out;
logic cond260_in;
logic cond260_write_en;
logic cond260_clk;
logic cond260_reset;
logic cond260_out;
logic cond260_done;
logic cond_wire260_in;
logic cond_wire260_out;
logic cond261_in;
logic cond261_write_en;
logic cond261_clk;
logic cond261_reset;
logic cond261_out;
logic cond261_done;
logic cond_wire261_in;
logic cond_wire261_out;
logic cond262_in;
logic cond262_write_en;
logic cond262_clk;
logic cond262_reset;
logic cond262_out;
logic cond262_done;
logic cond_wire262_in;
logic cond_wire262_out;
logic cond263_in;
logic cond263_write_en;
logic cond263_clk;
logic cond263_reset;
logic cond263_out;
logic cond263_done;
logic cond_wire263_in;
logic cond_wire263_out;
logic cond264_in;
logic cond264_write_en;
logic cond264_clk;
logic cond264_reset;
logic cond264_out;
logic cond264_done;
logic cond_wire264_in;
logic cond_wire264_out;
logic cond265_in;
logic cond265_write_en;
logic cond265_clk;
logic cond265_reset;
logic cond265_out;
logic cond265_done;
logic cond_wire265_in;
logic cond_wire265_out;
logic cond266_in;
logic cond266_write_en;
logic cond266_clk;
logic cond266_reset;
logic cond266_out;
logic cond266_done;
logic cond_wire266_in;
logic cond_wire266_out;
logic cond267_in;
logic cond267_write_en;
logic cond267_clk;
logic cond267_reset;
logic cond267_out;
logic cond267_done;
logic cond_wire267_in;
logic cond_wire267_out;
logic cond268_in;
logic cond268_write_en;
logic cond268_clk;
logic cond268_reset;
logic cond268_out;
logic cond268_done;
logic cond_wire268_in;
logic cond_wire268_out;
logic fsm_in;
logic fsm_write_en;
logic fsm_clk;
logic fsm_reset;
logic fsm_out;
logic fsm_done;
logic [4:0] fsm0_in;
logic fsm0_write_en;
logic fsm0_clk;
logic fsm0_reset;
logic [4:0] fsm0_out;
logic fsm0_done;
logic ud_out;
logic [4:0] adder_left;
logic [4:0] adder_right;
logic [4:0] adder_out;
logic ud0_out;
logic adder0_left;
logic adder0_right;
logic adder0_out;
logic signal_reg_in;
logic signal_reg_write_en;
logic signal_reg_clk;
logic signal_reg_reset;
logic signal_reg_out;
logic signal_reg_done;
logic early_reset_static_seq_go_in;
logic early_reset_static_seq_go_out;
logic early_reset_static_seq_done_in;
logic early_reset_static_seq_done_out;
logic early_reset_static_par0_go_in;
logic early_reset_static_par0_go_out;
logic early_reset_static_par0_done_in;
logic early_reset_static_par0_done_out;
logic wrapper_early_reset_static_seq_go_in;
logic wrapper_early_reset_static_seq_go_out;
logic wrapper_early_reset_static_seq_done_in;
logic wrapper_early_reset_static_seq_done_out;
mac_pe pe_0_0 (
    .clk(pe_0_0_clk),
    .done(pe_0_0_done),
    .go(pe_0_0_go),
    .left(pe_0_0_left),
    .mul_ready(pe_0_0_mul_ready),
    .out(pe_0_0_out),
    .reset(pe_0_0_reset),
    .top(pe_0_0_top)
);
std_reg # (
    .WIDTH(32)
) top_0_0 (
    .clk(top_0_0_clk),
    .done(top_0_0_done),
    .in(top_0_0_in),
    .out(top_0_0_out),
    .reset(top_0_0_reset),
    .write_en(top_0_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_0 (
    .clk(left_0_0_clk),
    .done(left_0_0_done),
    .in(left_0_0_in),
    .out(left_0_0_out),
    .reset(left_0_0_reset),
    .write_en(left_0_0_write_en)
);
mac_pe pe_0_1 (
    .clk(pe_0_1_clk),
    .done(pe_0_1_done),
    .go(pe_0_1_go),
    .left(pe_0_1_left),
    .mul_ready(pe_0_1_mul_ready),
    .out(pe_0_1_out),
    .reset(pe_0_1_reset),
    .top(pe_0_1_top)
);
std_reg # (
    .WIDTH(32)
) top_0_1 (
    .clk(top_0_1_clk),
    .done(top_0_1_done),
    .in(top_0_1_in),
    .out(top_0_1_out),
    .reset(top_0_1_reset),
    .write_en(top_0_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_1 (
    .clk(left_0_1_clk),
    .done(left_0_1_done),
    .in(left_0_1_in),
    .out(left_0_1_out),
    .reset(left_0_1_reset),
    .write_en(left_0_1_write_en)
);
mac_pe pe_0_2 (
    .clk(pe_0_2_clk),
    .done(pe_0_2_done),
    .go(pe_0_2_go),
    .left(pe_0_2_left),
    .mul_ready(pe_0_2_mul_ready),
    .out(pe_0_2_out),
    .reset(pe_0_2_reset),
    .top(pe_0_2_top)
);
std_reg # (
    .WIDTH(32)
) top_0_2 (
    .clk(top_0_2_clk),
    .done(top_0_2_done),
    .in(top_0_2_in),
    .out(top_0_2_out),
    .reset(top_0_2_reset),
    .write_en(top_0_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_2 (
    .clk(left_0_2_clk),
    .done(left_0_2_done),
    .in(left_0_2_in),
    .out(left_0_2_out),
    .reset(left_0_2_reset),
    .write_en(left_0_2_write_en)
);
mac_pe pe_0_3 (
    .clk(pe_0_3_clk),
    .done(pe_0_3_done),
    .go(pe_0_3_go),
    .left(pe_0_3_left),
    .mul_ready(pe_0_3_mul_ready),
    .out(pe_0_3_out),
    .reset(pe_0_3_reset),
    .top(pe_0_3_top)
);
std_reg # (
    .WIDTH(32)
) top_0_3 (
    .clk(top_0_3_clk),
    .done(top_0_3_done),
    .in(top_0_3_in),
    .out(top_0_3_out),
    .reset(top_0_3_reset),
    .write_en(top_0_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_3 (
    .clk(left_0_3_clk),
    .done(left_0_3_done),
    .in(left_0_3_in),
    .out(left_0_3_out),
    .reset(left_0_3_reset),
    .write_en(left_0_3_write_en)
);
mac_pe pe_0_4 (
    .clk(pe_0_4_clk),
    .done(pe_0_4_done),
    .go(pe_0_4_go),
    .left(pe_0_4_left),
    .mul_ready(pe_0_4_mul_ready),
    .out(pe_0_4_out),
    .reset(pe_0_4_reset),
    .top(pe_0_4_top)
);
std_reg # (
    .WIDTH(32)
) top_0_4 (
    .clk(top_0_4_clk),
    .done(top_0_4_done),
    .in(top_0_4_in),
    .out(top_0_4_out),
    .reset(top_0_4_reset),
    .write_en(top_0_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_4 (
    .clk(left_0_4_clk),
    .done(left_0_4_done),
    .in(left_0_4_in),
    .out(left_0_4_out),
    .reset(left_0_4_reset),
    .write_en(left_0_4_write_en)
);
mac_pe pe_0_5 (
    .clk(pe_0_5_clk),
    .done(pe_0_5_done),
    .go(pe_0_5_go),
    .left(pe_0_5_left),
    .mul_ready(pe_0_5_mul_ready),
    .out(pe_0_5_out),
    .reset(pe_0_5_reset),
    .top(pe_0_5_top)
);
std_reg # (
    .WIDTH(32)
) top_0_5 (
    .clk(top_0_5_clk),
    .done(top_0_5_done),
    .in(top_0_5_in),
    .out(top_0_5_out),
    .reset(top_0_5_reset),
    .write_en(top_0_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_5 (
    .clk(left_0_5_clk),
    .done(left_0_5_done),
    .in(left_0_5_in),
    .out(left_0_5_out),
    .reset(left_0_5_reset),
    .write_en(left_0_5_write_en)
);
mac_pe pe_0_6 (
    .clk(pe_0_6_clk),
    .done(pe_0_6_done),
    .go(pe_0_6_go),
    .left(pe_0_6_left),
    .mul_ready(pe_0_6_mul_ready),
    .out(pe_0_6_out),
    .reset(pe_0_6_reset),
    .top(pe_0_6_top)
);
std_reg # (
    .WIDTH(32)
) top_0_6 (
    .clk(top_0_6_clk),
    .done(top_0_6_done),
    .in(top_0_6_in),
    .out(top_0_6_out),
    .reset(top_0_6_reset),
    .write_en(top_0_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_6 (
    .clk(left_0_6_clk),
    .done(left_0_6_done),
    .in(left_0_6_in),
    .out(left_0_6_out),
    .reset(left_0_6_reset),
    .write_en(left_0_6_write_en)
);
mac_pe pe_0_7 (
    .clk(pe_0_7_clk),
    .done(pe_0_7_done),
    .go(pe_0_7_go),
    .left(pe_0_7_left),
    .mul_ready(pe_0_7_mul_ready),
    .out(pe_0_7_out),
    .reset(pe_0_7_reset),
    .top(pe_0_7_top)
);
std_reg # (
    .WIDTH(32)
) top_0_7 (
    .clk(top_0_7_clk),
    .done(top_0_7_done),
    .in(top_0_7_in),
    .out(top_0_7_out),
    .reset(top_0_7_reset),
    .write_en(top_0_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_7 (
    .clk(left_0_7_clk),
    .done(left_0_7_done),
    .in(left_0_7_in),
    .out(left_0_7_out),
    .reset(left_0_7_reset),
    .write_en(left_0_7_write_en)
);
mac_pe pe_1_0 (
    .clk(pe_1_0_clk),
    .done(pe_1_0_done),
    .go(pe_1_0_go),
    .left(pe_1_0_left),
    .mul_ready(pe_1_0_mul_ready),
    .out(pe_1_0_out),
    .reset(pe_1_0_reset),
    .top(pe_1_0_top)
);
std_reg # (
    .WIDTH(32)
) top_1_0 (
    .clk(top_1_0_clk),
    .done(top_1_0_done),
    .in(top_1_0_in),
    .out(top_1_0_out),
    .reset(top_1_0_reset),
    .write_en(top_1_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_0 (
    .clk(left_1_0_clk),
    .done(left_1_0_done),
    .in(left_1_0_in),
    .out(left_1_0_out),
    .reset(left_1_0_reset),
    .write_en(left_1_0_write_en)
);
mac_pe pe_1_1 (
    .clk(pe_1_1_clk),
    .done(pe_1_1_done),
    .go(pe_1_1_go),
    .left(pe_1_1_left),
    .mul_ready(pe_1_1_mul_ready),
    .out(pe_1_1_out),
    .reset(pe_1_1_reset),
    .top(pe_1_1_top)
);
std_reg # (
    .WIDTH(32)
) top_1_1 (
    .clk(top_1_1_clk),
    .done(top_1_1_done),
    .in(top_1_1_in),
    .out(top_1_1_out),
    .reset(top_1_1_reset),
    .write_en(top_1_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_1 (
    .clk(left_1_1_clk),
    .done(left_1_1_done),
    .in(left_1_1_in),
    .out(left_1_1_out),
    .reset(left_1_1_reset),
    .write_en(left_1_1_write_en)
);
mac_pe pe_1_2 (
    .clk(pe_1_2_clk),
    .done(pe_1_2_done),
    .go(pe_1_2_go),
    .left(pe_1_2_left),
    .mul_ready(pe_1_2_mul_ready),
    .out(pe_1_2_out),
    .reset(pe_1_2_reset),
    .top(pe_1_2_top)
);
std_reg # (
    .WIDTH(32)
) top_1_2 (
    .clk(top_1_2_clk),
    .done(top_1_2_done),
    .in(top_1_2_in),
    .out(top_1_2_out),
    .reset(top_1_2_reset),
    .write_en(top_1_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_2 (
    .clk(left_1_2_clk),
    .done(left_1_2_done),
    .in(left_1_2_in),
    .out(left_1_2_out),
    .reset(left_1_2_reset),
    .write_en(left_1_2_write_en)
);
mac_pe pe_1_3 (
    .clk(pe_1_3_clk),
    .done(pe_1_3_done),
    .go(pe_1_3_go),
    .left(pe_1_3_left),
    .mul_ready(pe_1_3_mul_ready),
    .out(pe_1_3_out),
    .reset(pe_1_3_reset),
    .top(pe_1_3_top)
);
std_reg # (
    .WIDTH(32)
) top_1_3 (
    .clk(top_1_3_clk),
    .done(top_1_3_done),
    .in(top_1_3_in),
    .out(top_1_3_out),
    .reset(top_1_3_reset),
    .write_en(top_1_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_3 (
    .clk(left_1_3_clk),
    .done(left_1_3_done),
    .in(left_1_3_in),
    .out(left_1_3_out),
    .reset(left_1_3_reset),
    .write_en(left_1_3_write_en)
);
mac_pe pe_1_4 (
    .clk(pe_1_4_clk),
    .done(pe_1_4_done),
    .go(pe_1_4_go),
    .left(pe_1_4_left),
    .mul_ready(pe_1_4_mul_ready),
    .out(pe_1_4_out),
    .reset(pe_1_4_reset),
    .top(pe_1_4_top)
);
std_reg # (
    .WIDTH(32)
) top_1_4 (
    .clk(top_1_4_clk),
    .done(top_1_4_done),
    .in(top_1_4_in),
    .out(top_1_4_out),
    .reset(top_1_4_reset),
    .write_en(top_1_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_4 (
    .clk(left_1_4_clk),
    .done(left_1_4_done),
    .in(left_1_4_in),
    .out(left_1_4_out),
    .reset(left_1_4_reset),
    .write_en(left_1_4_write_en)
);
mac_pe pe_1_5 (
    .clk(pe_1_5_clk),
    .done(pe_1_5_done),
    .go(pe_1_5_go),
    .left(pe_1_5_left),
    .mul_ready(pe_1_5_mul_ready),
    .out(pe_1_5_out),
    .reset(pe_1_5_reset),
    .top(pe_1_5_top)
);
std_reg # (
    .WIDTH(32)
) top_1_5 (
    .clk(top_1_5_clk),
    .done(top_1_5_done),
    .in(top_1_5_in),
    .out(top_1_5_out),
    .reset(top_1_5_reset),
    .write_en(top_1_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_5 (
    .clk(left_1_5_clk),
    .done(left_1_5_done),
    .in(left_1_5_in),
    .out(left_1_5_out),
    .reset(left_1_5_reset),
    .write_en(left_1_5_write_en)
);
mac_pe pe_1_6 (
    .clk(pe_1_6_clk),
    .done(pe_1_6_done),
    .go(pe_1_6_go),
    .left(pe_1_6_left),
    .mul_ready(pe_1_6_mul_ready),
    .out(pe_1_6_out),
    .reset(pe_1_6_reset),
    .top(pe_1_6_top)
);
std_reg # (
    .WIDTH(32)
) top_1_6 (
    .clk(top_1_6_clk),
    .done(top_1_6_done),
    .in(top_1_6_in),
    .out(top_1_6_out),
    .reset(top_1_6_reset),
    .write_en(top_1_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_6 (
    .clk(left_1_6_clk),
    .done(left_1_6_done),
    .in(left_1_6_in),
    .out(left_1_6_out),
    .reset(left_1_6_reset),
    .write_en(left_1_6_write_en)
);
mac_pe pe_1_7 (
    .clk(pe_1_7_clk),
    .done(pe_1_7_done),
    .go(pe_1_7_go),
    .left(pe_1_7_left),
    .mul_ready(pe_1_7_mul_ready),
    .out(pe_1_7_out),
    .reset(pe_1_7_reset),
    .top(pe_1_7_top)
);
std_reg # (
    .WIDTH(32)
) top_1_7 (
    .clk(top_1_7_clk),
    .done(top_1_7_done),
    .in(top_1_7_in),
    .out(top_1_7_out),
    .reset(top_1_7_reset),
    .write_en(top_1_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_7 (
    .clk(left_1_7_clk),
    .done(left_1_7_done),
    .in(left_1_7_in),
    .out(left_1_7_out),
    .reset(left_1_7_reset),
    .write_en(left_1_7_write_en)
);
mac_pe pe_2_0 (
    .clk(pe_2_0_clk),
    .done(pe_2_0_done),
    .go(pe_2_0_go),
    .left(pe_2_0_left),
    .mul_ready(pe_2_0_mul_ready),
    .out(pe_2_0_out),
    .reset(pe_2_0_reset),
    .top(pe_2_0_top)
);
std_reg # (
    .WIDTH(32)
) top_2_0 (
    .clk(top_2_0_clk),
    .done(top_2_0_done),
    .in(top_2_0_in),
    .out(top_2_0_out),
    .reset(top_2_0_reset),
    .write_en(top_2_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_0 (
    .clk(left_2_0_clk),
    .done(left_2_0_done),
    .in(left_2_0_in),
    .out(left_2_0_out),
    .reset(left_2_0_reset),
    .write_en(left_2_0_write_en)
);
mac_pe pe_2_1 (
    .clk(pe_2_1_clk),
    .done(pe_2_1_done),
    .go(pe_2_1_go),
    .left(pe_2_1_left),
    .mul_ready(pe_2_1_mul_ready),
    .out(pe_2_1_out),
    .reset(pe_2_1_reset),
    .top(pe_2_1_top)
);
std_reg # (
    .WIDTH(32)
) top_2_1 (
    .clk(top_2_1_clk),
    .done(top_2_1_done),
    .in(top_2_1_in),
    .out(top_2_1_out),
    .reset(top_2_1_reset),
    .write_en(top_2_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_1 (
    .clk(left_2_1_clk),
    .done(left_2_1_done),
    .in(left_2_1_in),
    .out(left_2_1_out),
    .reset(left_2_1_reset),
    .write_en(left_2_1_write_en)
);
mac_pe pe_2_2 (
    .clk(pe_2_2_clk),
    .done(pe_2_2_done),
    .go(pe_2_2_go),
    .left(pe_2_2_left),
    .mul_ready(pe_2_2_mul_ready),
    .out(pe_2_2_out),
    .reset(pe_2_2_reset),
    .top(pe_2_2_top)
);
std_reg # (
    .WIDTH(32)
) top_2_2 (
    .clk(top_2_2_clk),
    .done(top_2_2_done),
    .in(top_2_2_in),
    .out(top_2_2_out),
    .reset(top_2_2_reset),
    .write_en(top_2_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_2 (
    .clk(left_2_2_clk),
    .done(left_2_2_done),
    .in(left_2_2_in),
    .out(left_2_2_out),
    .reset(left_2_2_reset),
    .write_en(left_2_2_write_en)
);
mac_pe pe_2_3 (
    .clk(pe_2_3_clk),
    .done(pe_2_3_done),
    .go(pe_2_3_go),
    .left(pe_2_3_left),
    .mul_ready(pe_2_3_mul_ready),
    .out(pe_2_3_out),
    .reset(pe_2_3_reset),
    .top(pe_2_3_top)
);
std_reg # (
    .WIDTH(32)
) top_2_3 (
    .clk(top_2_3_clk),
    .done(top_2_3_done),
    .in(top_2_3_in),
    .out(top_2_3_out),
    .reset(top_2_3_reset),
    .write_en(top_2_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_3 (
    .clk(left_2_3_clk),
    .done(left_2_3_done),
    .in(left_2_3_in),
    .out(left_2_3_out),
    .reset(left_2_3_reset),
    .write_en(left_2_3_write_en)
);
mac_pe pe_2_4 (
    .clk(pe_2_4_clk),
    .done(pe_2_4_done),
    .go(pe_2_4_go),
    .left(pe_2_4_left),
    .mul_ready(pe_2_4_mul_ready),
    .out(pe_2_4_out),
    .reset(pe_2_4_reset),
    .top(pe_2_4_top)
);
std_reg # (
    .WIDTH(32)
) top_2_4 (
    .clk(top_2_4_clk),
    .done(top_2_4_done),
    .in(top_2_4_in),
    .out(top_2_4_out),
    .reset(top_2_4_reset),
    .write_en(top_2_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_4 (
    .clk(left_2_4_clk),
    .done(left_2_4_done),
    .in(left_2_4_in),
    .out(left_2_4_out),
    .reset(left_2_4_reset),
    .write_en(left_2_4_write_en)
);
mac_pe pe_2_5 (
    .clk(pe_2_5_clk),
    .done(pe_2_5_done),
    .go(pe_2_5_go),
    .left(pe_2_5_left),
    .mul_ready(pe_2_5_mul_ready),
    .out(pe_2_5_out),
    .reset(pe_2_5_reset),
    .top(pe_2_5_top)
);
std_reg # (
    .WIDTH(32)
) top_2_5 (
    .clk(top_2_5_clk),
    .done(top_2_5_done),
    .in(top_2_5_in),
    .out(top_2_5_out),
    .reset(top_2_5_reset),
    .write_en(top_2_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_5 (
    .clk(left_2_5_clk),
    .done(left_2_5_done),
    .in(left_2_5_in),
    .out(left_2_5_out),
    .reset(left_2_5_reset),
    .write_en(left_2_5_write_en)
);
mac_pe pe_2_6 (
    .clk(pe_2_6_clk),
    .done(pe_2_6_done),
    .go(pe_2_6_go),
    .left(pe_2_6_left),
    .mul_ready(pe_2_6_mul_ready),
    .out(pe_2_6_out),
    .reset(pe_2_6_reset),
    .top(pe_2_6_top)
);
std_reg # (
    .WIDTH(32)
) top_2_6 (
    .clk(top_2_6_clk),
    .done(top_2_6_done),
    .in(top_2_6_in),
    .out(top_2_6_out),
    .reset(top_2_6_reset),
    .write_en(top_2_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_6 (
    .clk(left_2_6_clk),
    .done(left_2_6_done),
    .in(left_2_6_in),
    .out(left_2_6_out),
    .reset(left_2_6_reset),
    .write_en(left_2_6_write_en)
);
mac_pe pe_2_7 (
    .clk(pe_2_7_clk),
    .done(pe_2_7_done),
    .go(pe_2_7_go),
    .left(pe_2_7_left),
    .mul_ready(pe_2_7_mul_ready),
    .out(pe_2_7_out),
    .reset(pe_2_7_reset),
    .top(pe_2_7_top)
);
std_reg # (
    .WIDTH(32)
) top_2_7 (
    .clk(top_2_7_clk),
    .done(top_2_7_done),
    .in(top_2_7_in),
    .out(top_2_7_out),
    .reset(top_2_7_reset),
    .write_en(top_2_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_7 (
    .clk(left_2_7_clk),
    .done(left_2_7_done),
    .in(left_2_7_in),
    .out(left_2_7_out),
    .reset(left_2_7_reset),
    .write_en(left_2_7_write_en)
);
mac_pe pe_3_0 (
    .clk(pe_3_0_clk),
    .done(pe_3_0_done),
    .go(pe_3_0_go),
    .left(pe_3_0_left),
    .mul_ready(pe_3_0_mul_ready),
    .out(pe_3_0_out),
    .reset(pe_3_0_reset),
    .top(pe_3_0_top)
);
std_reg # (
    .WIDTH(32)
) top_3_0 (
    .clk(top_3_0_clk),
    .done(top_3_0_done),
    .in(top_3_0_in),
    .out(top_3_0_out),
    .reset(top_3_0_reset),
    .write_en(top_3_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_0 (
    .clk(left_3_0_clk),
    .done(left_3_0_done),
    .in(left_3_0_in),
    .out(left_3_0_out),
    .reset(left_3_0_reset),
    .write_en(left_3_0_write_en)
);
mac_pe pe_3_1 (
    .clk(pe_3_1_clk),
    .done(pe_3_1_done),
    .go(pe_3_1_go),
    .left(pe_3_1_left),
    .mul_ready(pe_3_1_mul_ready),
    .out(pe_3_1_out),
    .reset(pe_3_1_reset),
    .top(pe_3_1_top)
);
std_reg # (
    .WIDTH(32)
) top_3_1 (
    .clk(top_3_1_clk),
    .done(top_3_1_done),
    .in(top_3_1_in),
    .out(top_3_1_out),
    .reset(top_3_1_reset),
    .write_en(top_3_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_1 (
    .clk(left_3_1_clk),
    .done(left_3_1_done),
    .in(left_3_1_in),
    .out(left_3_1_out),
    .reset(left_3_1_reset),
    .write_en(left_3_1_write_en)
);
mac_pe pe_3_2 (
    .clk(pe_3_2_clk),
    .done(pe_3_2_done),
    .go(pe_3_2_go),
    .left(pe_3_2_left),
    .mul_ready(pe_3_2_mul_ready),
    .out(pe_3_2_out),
    .reset(pe_3_2_reset),
    .top(pe_3_2_top)
);
std_reg # (
    .WIDTH(32)
) top_3_2 (
    .clk(top_3_2_clk),
    .done(top_3_2_done),
    .in(top_3_2_in),
    .out(top_3_2_out),
    .reset(top_3_2_reset),
    .write_en(top_3_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_2 (
    .clk(left_3_2_clk),
    .done(left_3_2_done),
    .in(left_3_2_in),
    .out(left_3_2_out),
    .reset(left_3_2_reset),
    .write_en(left_3_2_write_en)
);
mac_pe pe_3_3 (
    .clk(pe_3_3_clk),
    .done(pe_3_3_done),
    .go(pe_3_3_go),
    .left(pe_3_3_left),
    .mul_ready(pe_3_3_mul_ready),
    .out(pe_3_3_out),
    .reset(pe_3_3_reset),
    .top(pe_3_3_top)
);
std_reg # (
    .WIDTH(32)
) top_3_3 (
    .clk(top_3_3_clk),
    .done(top_3_3_done),
    .in(top_3_3_in),
    .out(top_3_3_out),
    .reset(top_3_3_reset),
    .write_en(top_3_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_3 (
    .clk(left_3_3_clk),
    .done(left_3_3_done),
    .in(left_3_3_in),
    .out(left_3_3_out),
    .reset(left_3_3_reset),
    .write_en(left_3_3_write_en)
);
mac_pe pe_3_4 (
    .clk(pe_3_4_clk),
    .done(pe_3_4_done),
    .go(pe_3_4_go),
    .left(pe_3_4_left),
    .mul_ready(pe_3_4_mul_ready),
    .out(pe_3_4_out),
    .reset(pe_3_4_reset),
    .top(pe_3_4_top)
);
std_reg # (
    .WIDTH(32)
) top_3_4 (
    .clk(top_3_4_clk),
    .done(top_3_4_done),
    .in(top_3_4_in),
    .out(top_3_4_out),
    .reset(top_3_4_reset),
    .write_en(top_3_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_4 (
    .clk(left_3_4_clk),
    .done(left_3_4_done),
    .in(left_3_4_in),
    .out(left_3_4_out),
    .reset(left_3_4_reset),
    .write_en(left_3_4_write_en)
);
mac_pe pe_3_5 (
    .clk(pe_3_5_clk),
    .done(pe_3_5_done),
    .go(pe_3_5_go),
    .left(pe_3_5_left),
    .mul_ready(pe_3_5_mul_ready),
    .out(pe_3_5_out),
    .reset(pe_3_5_reset),
    .top(pe_3_5_top)
);
std_reg # (
    .WIDTH(32)
) top_3_5 (
    .clk(top_3_5_clk),
    .done(top_3_5_done),
    .in(top_3_5_in),
    .out(top_3_5_out),
    .reset(top_3_5_reset),
    .write_en(top_3_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_5 (
    .clk(left_3_5_clk),
    .done(left_3_5_done),
    .in(left_3_5_in),
    .out(left_3_5_out),
    .reset(left_3_5_reset),
    .write_en(left_3_5_write_en)
);
mac_pe pe_3_6 (
    .clk(pe_3_6_clk),
    .done(pe_3_6_done),
    .go(pe_3_6_go),
    .left(pe_3_6_left),
    .mul_ready(pe_3_6_mul_ready),
    .out(pe_3_6_out),
    .reset(pe_3_6_reset),
    .top(pe_3_6_top)
);
std_reg # (
    .WIDTH(32)
) top_3_6 (
    .clk(top_3_6_clk),
    .done(top_3_6_done),
    .in(top_3_6_in),
    .out(top_3_6_out),
    .reset(top_3_6_reset),
    .write_en(top_3_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_6 (
    .clk(left_3_6_clk),
    .done(left_3_6_done),
    .in(left_3_6_in),
    .out(left_3_6_out),
    .reset(left_3_6_reset),
    .write_en(left_3_6_write_en)
);
mac_pe pe_3_7 (
    .clk(pe_3_7_clk),
    .done(pe_3_7_done),
    .go(pe_3_7_go),
    .left(pe_3_7_left),
    .mul_ready(pe_3_7_mul_ready),
    .out(pe_3_7_out),
    .reset(pe_3_7_reset),
    .top(pe_3_7_top)
);
std_reg # (
    .WIDTH(32)
) top_3_7 (
    .clk(top_3_7_clk),
    .done(top_3_7_done),
    .in(top_3_7_in),
    .out(top_3_7_out),
    .reset(top_3_7_reset),
    .write_en(top_3_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_7 (
    .clk(left_3_7_clk),
    .done(left_3_7_done),
    .in(left_3_7_in),
    .out(left_3_7_out),
    .reset(left_3_7_reset),
    .write_en(left_3_7_write_en)
);
mac_pe pe_4_0 (
    .clk(pe_4_0_clk),
    .done(pe_4_0_done),
    .go(pe_4_0_go),
    .left(pe_4_0_left),
    .mul_ready(pe_4_0_mul_ready),
    .out(pe_4_0_out),
    .reset(pe_4_0_reset),
    .top(pe_4_0_top)
);
std_reg # (
    .WIDTH(32)
) top_4_0 (
    .clk(top_4_0_clk),
    .done(top_4_0_done),
    .in(top_4_0_in),
    .out(top_4_0_out),
    .reset(top_4_0_reset),
    .write_en(top_4_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_0 (
    .clk(left_4_0_clk),
    .done(left_4_0_done),
    .in(left_4_0_in),
    .out(left_4_0_out),
    .reset(left_4_0_reset),
    .write_en(left_4_0_write_en)
);
mac_pe pe_4_1 (
    .clk(pe_4_1_clk),
    .done(pe_4_1_done),
    .go(pe_4_1_go),
    .left(pe_4_1_left),
    .mul_ready(pe_4_1_mul_ready),
    .out(pe_4_1_out),
    .reset(pe_4_1_reset),
    .top(pe_4_1_top)
);
std_reg # (
    .WIDTH(32)
) top_4_1 (
    .clk(top_4_1_clk),
    .done(top_4_1_done),
    .in(top_4_1_in),
    .out(top_4_1_out),
    .reset(top_4_1_reset),
    .write_en(top_4_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_1 (
    .clk(left_4_1_clk),
    .done(left_4_1_done),
    .in(left_4_1_in),
    .out(left_4_1_out),
    .reset(left_4_1_reset),
    .write_en(left_4_1_write_en)
);
mac_pe pe_4_2 (
    .clk(pe_4_2_clk),
    .done(pe_4_2_done),
    .go(pe_4_2_go),
    .left(pe_4_2_left),
    .mul_ready(pe_4_2_mul_ready),
    .out(pe_4_2_out),
    .reset(pe_4_2_reset),
    .top(pe_4_2_top)
);
std_reg # (
    .WIDTH(32)
) top_4_2 (
    .clk(top_4_2_clk),
    .done(top_4_2_done),
    .in(top_4_2_in),
    .out(top_4_2_out),
    .reset(top_4_2_reset),
    .write_en(top_4_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_2 (
    .clk(left_4_2_clk),
    .done(left_4_2_done),
    .in(left_4_2_in),
    .out(left_4_2_out),
    .reset(left_4_2_reset),
    .write_en(left_4_2_write_en)
);
mac_pe pe_4_3 (
    .clk(pe_4_3_clk),
    .done(pe_4_3_done),
    .go(pe_4_3_go),
    .left(pe_4_3_left),
    .mul_ready(pe_4_3_mul_ready),
    .out(pe_4_3_out),
    .reset(pe_4_3_reset),
    .top(pe_4_3_top)
);
std_reg # (
    .WIDTH(32)
) top_4_3 (
    .clk(top_4_3_clk),
    .done(top_4_3_done),
    .in(top_4_3_in),
    .out(top_4_3_out),
    .reset(top_4_3_reset),
    .write_en(top_4_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_3 (
    .clk(left_4_3_clk),
    .done(left_4_3_done),
    .in(left_4_3_in),
    .out(left_4_3_out),
    .reset(left_4_3_reset),
    .write_en(left_4_3_write_en)
);
mac_pe pe_4_4 (
    .clk(pe_4_4_clk),
    .done(pe_4_4_done),
    .go(pe_4_4_go),
    .left(pe_4_4_left),
    .mul_ready(pe_4_4_mul_ready),
    .out(pe_4_4_out),
    .reset(pe_4_4_reset),
    .top(pe_4_4_top)
);
std_reg # (
    .WIDTH(32)
) top_4_4 (
    .clk(top_4_4_clk),
    .done(top_4_4_done),
    .in(top_4_4_in),
    .out(top_4_4_out),
    .reset(top_4_4_reset),
    .write_en(top_4_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_4 (
    .clk(left_4_4_clk),
    .done(left_4_4_done),
    .in(left_4_4_in),
    .out(left_4_4_out),
    .reset(left_4_4_reset),
    .write_en(left_4_4_write_en)
);
mac_pe pe_4_5 (
    .clk(pe_4_5_clk),
    .done(pe_4_5_done),
    .go(pe_4_5_go),
    .left(pe_4_5_left),
    .mul_ready(pe_4_5_mul_ready),
    .out(pe_4_5_out),
    .reset(pe_4_5_reset),
    .top(pe_4_5_top)
);
std_reg # (
    .WIDTH(32)
) top_4_5 (
    .clk(top_4_5_clk),
    .done(top_4_5_done),
    .in(top_4_5_in),
    .out(top_4_5_out),
    .reset(top_4_5_reset),
    .write_en(top_4_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_5 (
    .clk(left_4_5_clk),
    .done(left_4_5_done),
    .in(left_4_5_in),
    .out(left_4_5_out),
    .reset(left_4_5_reset),
    .write_en(left_4_5_write_en)
);
mac_pe pe_4_6 (
    .clk(pe_4_6_clk),
    .done(pe_4_6_done),
    .go(pe_4_6_go),
    .left(pe_4_6_left),
    .mul_ready(pe_4_6_mul_ready),
    .out(pe_4_6_out),
    .reset(pe_4_6_reset),
    .top(pe_4_6_top)
);
std_reg # (
    .WIDTH(32)
) top_4_6 (
    .clk(top_4_6_clk),
    .done(top_4_6_done),
    .in(top_4_6_in),
    .out(top_4_6_out),
    .reset(top_4_6_reset),
    .write_en(top_4_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_6 (
    .clk(left_4_6_clk),
    .done(left_4_6_done),
    .in(left_4_6_in),
    .out(left_4_6_out),
    .reset(left_4_6_reset),
    .write_en(left_4_6_write_en)
);
mac_pe pe_4_7 (
    .clk(pe_4_7_clk),
    .done(pe_4_7_done),
    .go(pe_4_7_go),
    .left(pe_4_7_left),
    .mul_ready(pe_4_7_mul_ready),
    .out(pe_4_7_out),
    .reset(pe_4_7_reset),
    .top(pe_4_7_top)
);
std_reg # (
    .WIDTH(32)
) top_4_7 (
    .clk(top_4_7_clk),
    .done(top_4_7_done),
    .in(top_4_7_in),
    .out(top_4_7_out),
    .reset(top_4_7_reset),
    .write_en(top_4_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_7 (
    .clk(left_4_7_clk),
    .done(left_4_7_done),
    .in(left_4_7_in),
    .out(left_4_7_out),
    .reset(left_4_7_reset),
    .write_en(left_4_7_write_en)
);
mac_pe pe_5_0 (
    .clk(pe_5_0_clk),
    .done(pe_5_0_done),
    .go(pe_5_0_go),
    .left(pe_5_0_left),
    .mul_ready(pe_5_0_mul_ready),
    .out(pe_5_0_out),
    .reset(pe_5_0_reset),
    .top(pe_5_0_top)
);
std_reg # (
    .WIDTH(32)
) top_5_0 (
    .clk(top_5_0_clk),
    .done(top_5_0_done),
    .in(top_5_0_in),
    .out(top_5_0_out),
    .reset(top_5_0_reset),
    .write_en(top_5_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_0 (
    .clk(left_5_0_clk),
    .done(left_5_0_done),
    .in(left_5_0_in),
    .out(left_5_0_out),
    .reset(left_5_0_reset),
    .write_en(left_5_0_write_en)
);
mac_pe pe_5_1 (
    .clk(pe_5_1_clk),
    .done(pe_5_1_done),
    .go(pe_5_1_go),
    .left(pe_5_1_left),
    .mul_ready(pe_5_1_mul_ready),
    .out(pe_5_1_out),
    .reset(pe_5_1_reset),
    .top(pe_5_1_top)
);
std_reg # (
    .WIDTH(32)
) top_5_1 (
    .clk(top_5_1_clk),
    .done(top_5_1_done),
    .in(top_5_1_in),
    .out(top_5_1_out),
    .reset(top_5_1_reset),
    .write_en(top_5_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_1 (
    .clk(left_5_1_clk),
    .done(left_5_1_done),
    .in(left_5_1_in),
    .out(left_5_1_out),
    .reset(left_5_1_reset),
    .write_en(left_5_1_write_en)
);
mac_pe pe_5_2 (
    .clk(pe_5_2_clk),
    .done(pe_5_2_done),
    .go(pe_5_2_go),
    .left(pe_5_2_left),
    .mul_ready(pe_5_2_mul_ready),
    .out(pe_5_2_out),
    .reset(pe_5_2_reset),
    .top(pe_5_2_top)
);
std_reg # (
    .WIDTH(32)
) top_5_2 (
    .clk(top_5_2_clk),
    .done(top_5_2_done),
    .in(top_5_2_in),
    .out(top_5_2_out),
    .reset(top_5_2_reset),
    .write_en(top_5_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_2 (
    .clk(left_5_2_clk),
    .done(left_5_2_done),
    .in(left_5_2_in),
    .out(left_5_2_out),
    .reset(left_5_2_reset),
    .write_en(left_5_2_write_en)
);
mac_pe pe_5_3 (
    .clk(pe_5_3_clk),
    .done(pe_5_3_done),
    .go(pe_5_3_go),
    .left(pe_5_3_left),
    .mul_ready(pe_5_3_mul_ready),
    .out(pe_5_3_out),
    .reset(pe_5_3_reset),
    .top(pe_5_3_top)
);
std_reg # (
    .WIDTH(32)
) top_5_3 (
    .clk(top_5_3_clk),
    .done(top_5_3_done),
    .in(top_5_3_in),
    .out(top_5_3_out),
    .reset(top_5_3_reset),
    .write_en(top_5_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_3 (
    .clk(left_5_3_clk),
    .done(left_5_3_done),
    .in(left_5_3_in),
    .out(left_5_3_out),
    .reset(left_5_3_reset),
    .write_en(left_5_3_write_en)
);
mac_pe pe_5_4 (
    .clk(pe_5_4_clk),
    .done(pe_5_4_done),
    .go(pe_5_4_go),
    .left(pe_5_4_left),
    .mul_ready(pe_5_4_mul_ready),
    .out(pe_5_4_out),
    .reset(pe_5_4_reset),
    .top(pe_5_4_top)
);
std_reg # (
    .WIDTH(32)
) top_5_4 (
    .clk(top_5_4_clk),
    .done(top_5_4_done),
    .in(top_5_4_in),
    .out(top_5_4_out),
    .reset(top_5_4_reset),
    .write_en(top_5_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_4 (
    .clk(left_5_4_clk),
    .done(left_5_4_done),
    .in(left_5_4_in),
    .out(left_5_4_out),
    .reset(left_5_4_reset),
    .write_en(left_5_4_write_en)
);
mac_pe pe_5_5 (
    .clk(pe_5_5_clk),
    .done(pe_5_5_done),
    .go(pe_5_5_go),
    .left(pe_5_5_left),
    .mul_ready(pe_5_5_mul_ready),
    .out(pe_5_5_out),
    .reset(pe_5_5_reset),
    .top(pe_5_5_top)
);
std_reg # (
    .WIDTH(32)
) top_5_5 (
    .clk(top_5_5_clk),
    .done(top_5_5_done),
    .in(top_5_5_in),
    .out(top_5_5_out),
    .reset(top_5_5_reset),
    .write_en(top_5_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_5 (
    .clk(left_5_5_clk),
    .done(left_5_5_done),
    .in(left_5_5_in),
    .out(left_5_5_out),
    .reset(left_5_5_reset),
    .write_en(left_5_5_write_en)
);
mac_pe pe_5_6 (
    .clk(pe_5_6_clk),
    .done(pe_5_6_done),
    .go(pe_5_6_go),
    .left(pe_5_6_left),
    .mul_ready(pe_5_6_mul_ready),
    .out(pe_5_6_out),
    .reset(pe_5_6_reset),
    .top(pe_5_6_top)
);
std_reg # (
    .WIDTH(32)
) top_5_6 (
    .clk(top_5_6_clk),
    .done(top_5_6_done),
    .in(top_5_6_in),
    .out(top_5_6_out),
    .reset(top_5_6_reset),
    .write_en(top_5_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_6 (
    .clk(left_5_6_clk),
    .done(left_5_6_done),
    .in(left_5_6_in),
    .out(left_5_6_out),
    .reset(left_5_6_reset),
    .write_en(left_5_6_write_en)
);
mac_pe pe_5_7 (
    .clk(pe_5_7_clk),
    .done(pe_5_7_done),
    .go(pe_5_7_go),
    .left(pe_5_7_left),
    .mul_ready(pe_5_7_mul_ready),
    .out(pe_5_7_out),
    .reset(pe_5_7_reset),
    .top(pe_5_7_top)
);
std_reg # (
    .WIDTH(32)
) top_5_7 (
    .clk(top_5_7_clk),
    .done(top_5_7_done),
    .in(top_5_7_in),
    .out(top_5_7_out),
    .reset(top_5_7_reset),
    .write_en(top_5_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_7 (
    .clk(left_5_7_clk),
    .done(left_5_7_done),
    .in(left_5_7_in),
    .out(left_5_7_out),
    .reset(left_5_7_reset),
    .write_en(left_5_7_write_en)
);
mac_pe pe_6_0 (
    .clk(pe_6_0_clk),
    .done(pe_6_0_done),
    .go(pe_6_0_go),
    .left(pe_6_0_left),
    .mul_ready(pe_6_0_mul_ready),
    .out(pe_6_0_out),
    .reset(pe_6_0_reset),
    .top(pe_6_0_top)
);
std_reg # (
    .WIDTH(32)
) top_6_0 (
    .clk(top_6_0_clk),
    .done(top_6_0_done),
    .in(top_6_0_in),
    .out(top_6_0_out),
    .reset(top_6_0_reset),
    .write_en(top_6_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_0 (
    .clk(left_6_0_clk),
    .done(left_6_0_done),
    .in(left_6_0_in),
    .out(left_6_0_out),
    .reset(left_6_0_reset),
    .write_en(left_6_0_write_en)
);
mac_pe pe_6_1 (
    .clk(pe_6_1_clk),
    .done(pe_6_1_done),
    .go(pe_6_1_go),
    .left(pe_6_1_left),
    .mul_ready(pe_6_1_mul_ready),
    .out(pe_6_1_out),
    .reset(pe_6_1_reset),
    .top(pe_6_1_top)
);
std_reg # (
    .WIDTH(32)
) top_6_1 (
    .clk(top_6_1_clk),
    .done(top_6_1_done),
    .in(top_6_1_in),
    .out(top_6_1_out),
    .reset(top_6_1_reset),
    .write_en(top_6_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_1 (
    .clk(left_6_1_clk),
    .done(left_6_1_done),
    .in(left_6_1_in),
    .out(left_6_1_out),
    .reset(left_6_1_reset),
    .write_en(left_6_1_write_en)
);
mac_pe pe_6_2 (
    .clk(pe_6_2_clk),
    .done(pe_6_2_done),
    .go(pe_6_2_go),
    .left(pe_6_2_left),
    .mul_ready(pe_6_2_mul_ready),
    .out(pe_6_2_out),
    .reset(pe_6_2_reset),
    .top(pe_6_2_top)
);
std_reg # (
    .WIDTH(32)
) top_6_2 (
    .clk(top_6_2_clk),
    .done(top_6_2_done),
    .in(top_6_2_in),
    .out(top_6_2_out),
    .reset(top_6_2_reset),
    .write_en(top_6_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_2 (
    .clk(left_6_2_clk),
    .done(left_6_2_done),
    .in(left_6_2_in),
    .out(left_6_2_out),
    .reset(left_6_2_reset),
    .write_en(left_6_2_write_en)
);
mac_pe pe_6_3 (
    .clk(pe_6_3_clk),
    .done(pe_6_3_done),
    .go(pe_6_3_go),
    .left(pe_6_3_left),
    .mul_ready(pe_6_3_mul_ready),
    .out(pe_6_3_out),
    .reset(pe_6_3_reset),
    .top(pe_6_3_top)
);
std_reg # (
    .WIDTH(32)
) top_6_3 (
    .clk(top_6_3_clk),
    .done(top_6_3_done),
    .in(top_6_3_in),
    .out(top_6_3_out),
    .reset(top_6_3_reset),
    .write_en(top_6_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_3 (
    .clk(left_6_3_clk),
    .done(left_6_3_done),
    .in(left_6_3_in),
    .out(left_6_3_out),
    .reset(left_6_3_reset),
    .write_en(left_6_3_write_en)
);
mac_pe pe_6_4 (
    .clk(pe_6_4_clk),
    .done(pe_6_4_done),
    .go(pe_6_4_go),
    .left(pe_6_4_left),
    .mul_ready(pe_6_4_mul_ready),
    .out(pe_6_4_out),
    .reset(pe_6_4_reset),
    .top(pe_6_4_top)
);
std_reg # (
    .WIDTH(32)
) top_6_4 (
    .clk(top_6_4_clk),
    .done(top_6_4_done),
    .in(top_6_4_in),
    .out(top_6_4_out),
    .reset(top_6_4_reset),
    .write_en(top_6_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_4 (
    .clk(left_6_4_clk),
    .done(left_6_4_done),
    .in(left_6_4_in),
    .out(left_6_4_out),
    .reset(left_6_4_reset),
    .write_en(left_6_4_write_en)
);
mac_pe pe_6_5 (
    .clk(pe_6_5_clk),
    .done(pe_6_5_done),
    .go(pe_6_5_go),
    .left(pe_6_5_left),
    .mul_ready(pe_6_5_mul_ready),
    .out(pe_6_5_out),
    .reset(pe_6_5_reset),
    .top(pe_6_5_top)
);
std_reg # (
    .WIDTH(32)
) top_6_5 (
    .clk(top_6_5_clk),
    .done(top_6_5_done),
    .in(top_6_5_in),
    .out(top_6_5_out),
    .reset(top_6_5_reset),
    .write_en(top_6_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_5 (
    .clk(left_6_5_clk),
    .done(left_6_5_done),
    .in(left_6_5_in),
    .out(left_6_5_out),
    .reset(left_6_5_reset),
    .write_en(left_6_5_write_en)
);
mac_pe pe_6_6 (
    .clk(pe_6_6_clk),
    .done(pe_6_6_done),
    .go(pe_6_6_go),
    .left(pe_6_6_left),
    .mul_ready(pe_6_6_mul_ready),
    .out(pe_6_6_out),
    .reset(pe_6_6_reset),
    .top(pe_6_6_top)
);
std_reg # (
    .WIDTH(32)
) top_6_6 (
    .clk(top_6_6_clk),
    .done(top_6_6_done),
    .in(top_6_6_in),
    .out(top_6_6_out),
    .reset(top_6_6_reset),
    .write_en(top_6_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_6 (
    .clk(left_6_6_clk),
    .done(left_6_6_done),
    .in(left_6_6_in),
    .out(left_6_6_out),
    .reset(left_6_6_reset),
    .write_en(left_6_6_write_en)
);
mac_pe pe_6_7 (
    .clk(pe_6_7_clk),
    .done(pe_6_7_done),
    .go(pe_6_7_go),
    .left(pe_6_7_left),
    .mul_ready(pe_6_7_mul_ready),
    .out(pe_6_7_out),
    .reset(pe_6_7_reset),
    .top(pe_6_7_top)
);
std_reg # (
    .WIDTH(32)
) top_6_7 (
    .clk(top_6_7_clk),
    .done(top_6_7_done),
    .in(top_6_7_in),
    .out(top_6_7_out),
    .reset(top_6_7_reset),
    .write_en(top_6_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_7 (
    .clk(left_6_7_clk),
    .done(left_6_7_done),
    .in(left_6_7_in),
    .out(left_6_7_out),
    .reset(left_6_7_reset),
    .write_en(left_6_7_write_en)
);
mac_pe pe_7_0 (
    .clk(pe_7_0_clk),
    .done(pe_7_0_done),
    .go(pe_7_0_go),
    .left(pe_7_0_left),
    .mul_ready(pe_7_0_mul_ready),
    .out(pe_7_0_out),
    .reset(pe_7_0_reset),
    .top(pe_7_0_top)
);
std_reg # (
    .WIDTH(32)
) top_7_0 (
    .clk(top_7_0_clk),
    .done(top_7_0_done),
    .in(top_7_0_in),
    .out(top_7_0_out),
    .reset(top_7_0_reset),
    .write_en(top_7_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_0 (
    .clk(left_7_0_clk),
    .done(left_7_0_done),
    .in(left_7_0_in),
    .out(left_7_0_out),
    .reset(left_7_0_reset),
    .write_en(left_7_0_write_en)
);
mac_pe pe_7_1 (
    .clk(pe_7_1_clk),
    .done(pe_7_1_done),
    .go(pe_7_1_go),
    .left(pe_7_1_left),
    .mul_ready(pe_7_1_mul_ready),
    .out(pe_7_1_out),
    .reset(pe_7_1_reset),
    .top(pe_7_1_top)
);
std_reg # (
    .WIDTH(32)
) top_7_1 (
    .clk(top_7_1_clk),
    .done(top_7_1_done),
    .in(top_7_1_in),
    .out(top_7_1_out),
    .reset(top_7_1_reset),
    .write_en(top_7_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_1 (
    .clk(left_7_1_clk),
    .done(left_7_1_done),
    .in(left_7_1_in),
    .out(left_7_1_out),
    .reset(left_7_1_reset),
    .write_en(left_7_1_write_en)
);
mac_pe pe_7_2 (
    .clk(pe_7_2_clk),
    .done(pe_7_2_done),
    .go(pe_7_2_go),
    .left(pe_7_2_left),
    .mul_ready(pe_7_2_mul_ready),
    .out(pe_7_2_out),
    .reset(pe_7_2_reset),
    .top(pe_7_2_top)
);
std_reg # (
    .WIDTH(32)
) top_7_2 (
    .clk(top_7_2_clk),
    .done(top_7_2_done),
    .in(top_7_2_in),
    .out(top_7_2_out),
    .reset(top_7_2_reset),
    .write_en(top_7_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_2 (
    .clk(left_7_2_clk),
    .done(left_7_2_done),
    .in(left_7_2_in),
    .out(left_7_2_out),
    .reset(left_7_2_reset),
    .write_en(left_7_2_write_en)
);
mac_pe pe_7_3 (
    .clk(pe_7_3_clk),
    .done(pe_7_3_done),
    .go(pe_7_3_go),
    .left(pe_7_3_left),
    .mul_ready(pe_7_3_mul_ready),
    .out(pe_7_3_out),
    .reset(pe_7_3_reset),
    .top(pe_7_3_top)
);
std_reg # (
    .WIDTH(32)
) top_7_3 (
    .clk(top_7_3_clk),
    .done(top_7_3_done),
    .in(top_7_3_in),
    .out(top_7_3_out),
    .reset(top_7_3_reset),
    .write_en(top_7_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_3 (
    .clk(left_7_3_clk),
    .done(left_7_3_done),
    .in(left_7_3_in),
    .out(left_7_3_out),
    .reset(left_7_3_reset),
    .write_en(left_7_3_write_en)
);
mac_pe pe_7_4 (
    .clk(pe_7_4_clk),
    .done(pe_7_4_done),
    .go(pe_7_4_go),
    .left(pe_7_4_left),
    .mul_ready(pe_7_4_mul_ready),
    .out(pe_7_4_out),
    .reset(pe_7_4_reset),
    .top(pe_7_4_top)
);
std_reg # (
    .WIDTH(32)
) top_7_4 (
    .clk(top_7_4_clk),
    .done(top_7_4_done),
    .in(top_7_4_in),
    .out(top_7_4_out),
    .reset(top_7_4_reset),
    .write_en(top_7_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_4 (
    .clk(left_7_4_clk),
    .done(left_7_4_done),
    .in(left_7_4_in),
    .out(left_7_4_out),
    .reset(left_7_4_reset),
    .write_en(left_7_4_write_en)
);
mac_pe pe_7_5 (
    .clk(pe_7_5_clk),
    .done(pe_7_5_done),
    .go(pe_7_5_go),
    .left(pe_7_5_left),
    .mul_ready(pe_7_5_mul_ready),
    .out(pe_7_5_out),
    .reset(pe_7_5_reset),
    .top(pe_7_5_top)
);
std_reg # (
    .WIDTH(32)
) top_7_5 (
    .clk(top_7_5_clk),
    .done(top_7_5_done),
    .in(top_7_5_in),
    .out(top_7_5_out),
    .reset(top_7_5_reset),
    .write_en(top_7_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_5 (
    .clk(left_7_5_clk),
    .done(left_7_5_done),
    .in(left_7_5_in),
    .out(left_7_5_out),
    .reset(left_7_5_reset),
    .write_en(left_7_5_write_en)
);
mac_pe pe_7_6 (
    .clk(pe_7_6_clk),
    .done(pe_7_6_done),
    .go(pe_7_6_go),
    .left(pe_7_6_left),
    .mul_ready(pe_7_6_mul_ready),
    .out(pe_7_6_out),
    .reset(pe_7_6_reset),
    .top(pe_7_6_top)
);
std_reg # (
    .WIDTH(32)
) top_7_6 (
    .clk(top_7_6_clk),
    .done(top_7_6_done),
    .in(top_7_6_in),
    .out(top_7_6_out),
    .reset(top_7_6_reset),
    .write_en(top_7_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_6 (
    .clk(left_7_6_clk),
    .done(left_7_6_done),
    .in(left_7_6_in),
    .out(left_7_6_out),
    .reset(left_7_6_reset),
    .write_en(left_7_6_write_en)
);
mac_pe pe_7_7 (
    .clk(pe_7_7_clk),
    .done(pe_7_7_done),
    .go(pe_7_7_go),
    .left(pe_7_7_left),
    .mul_ready(pe_7_7_mul_ready),
    .out(pe_7_7_out),
    .reset(pe_7_7_reset),
    .top(pe_7_7_top)
);
std_reg # (
    .WIDTH(32)
) top_7_7 (
    .clk(top_7_7_clk),
    .done(top_7_7_done),
    .in(top_7_7_in),
    .out(top_7_7_out),
    .reset(top_7_7_reset),
    .write_en(top_7_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_7 (
    .clk(left_7_7_clk),
    .done(left_7_7_done),
    .in(left_7_7_in),
    .out(left_7_7_out),
    .reset(left_7_7_reset),
    .write_en(left_7_7_write_en)
);
std_reg # (
    .WIDTH(4)
) t0_idx (
    .clk(t0_idx_clk),
    .done(t0_idx_done),
    .in(t0_idx_in),
    .out(t0_idx_out),
    .reset(t0_idx_reset),
    .write_en(t0_idx_write_en)
);
std_add # (
    .WIDTH(4)
) t0_add (
    .left(t0_add_left),
    .out(t0_add_out),
    .right(t0_add_right)
);
std_reg # (
    .WIDTH(4)
) t1_idx (
    .clk(t1_idx_clk),
    .done(t1_idx_done),
    .in(t1_idx_in),
    .out(t1_idx_out),
    .reset(t1_idx_reset),
    .write_en(t1_idx_write_en)
);
std_add # (
    .WIDTH(4)
) t1_add (
    .left(t1_add_left),
    .out(t1_add_out),
    .right(t1_add_right)
);
std_reg # (
    .WIDTH(4)
) t2_idx (
    .clk(t2_idx_clk),
    .done(t2_idx_done),
    .in(t2_idx_in),
    .out(t2_idx_out),
    .reset(t2_idx_reset),
    .write_en(t2_idx_write_en)
);
std_add # (
    .WIDTH(4)
) t2_add (
    .left(t2_add_left),
    .out(t2_add_out),
    .right(t2_add_right)
);
std_reg # (
    .WIDTH(4)
) t3_idx (
    .clk(t3_idx_clk),
    .done(t3_idx_done),
    .in(t3_idx_in),
    .out(t3_idx_out),
    .reset(t3_idx_reset),
    .write_en(t3_idx_write_en)
);
std_add # (
    .WIDTH(4)
) t3_add (
    .left(t3_add_left),
    .out(t3_add_out),
    .right(t3_add_right)
);
std_reg # (
    .WIDTH(4)
) t4_idx (
    .clk(t4_idx_clk),
    .done(t4_idx_done),
    .in(t4_idx_in),
    .out(t4_idx_out),
    .reset(t4_idx_reset),
    .write_en(t4_idx_write_en)
);
std_add # (
    .WIDTH(4)
) t4_add (
    .left(t4_add_left),
    .out(t4_add_out),
    .right(t4_add_right)
);
std_reg # (
    .WIDTH(4)
) t5_idx (
    .clk(t5_idx_clk),
    .done(t5_idx_done),
    .in(t5_idx_in),
    .out(t5_idx_out),
    .reset(t5_idx_reset),
    .write_en(t5_idx_write_en)
);
std_add # (
    .WIDTH(4)
) t5_add (
    .left(t5_add_left),
    .out(t5_add_out),
    .right(t5_add_right)
);
std_reg # (
    .WIDTH(4)
) t6_idx (
    .clk(t6_idx_clk),
    .done(t6_idx_done),
    .in(t6_idx_in),
    .out(t6_idx_out),
    .reset(t6_idx_reset),
    .write_en(t6_idx_write_en)
);
std_add # (
    .WIDTH(4)
) t6_add (
    .left(t6_add_left),
    .out(t6_add_out),
    .right(t6_add_right)
);
std_reg # (
    .WIDTH(4)
) t7_idx (
    .clk(t7_idx_clk),
    .done(t7_idx_done),
    .in(t7_idx_in),
    .out(t7_idx_out),
    .reset(t7_idx_reset),
    .write_en(t7_idx_write_en)
);
std_add # (
    .WIDTH(4)
) t7_add (
    .left(t7_add_left),
    .out(t7_add_out),
    .right(t7_add_right)
);
std_reg # (
    .WIDTH(4)
) l0_idx (
    .clk(l0_idx_clk),
    .done(l0_idx_done),
    .in(l0_idx_in),
    .out(l0_idx_out),
    .reset(l0_idx_reset),
    .write_en(l0_idx_write_en)
);
std_add # (
    .WIDTH(4)
) l0_add (
    .left(l0_add_left),
    .out(l0_add_out),
    .right(l0_add_right)
);
std_reg # (
    .WIDTH(4)
) l1_idx (
    .clk(l1_idx_clk),
    .done(l1_idx_done),
    .in(l1_idx_in),
    .out(l1_idx_out),
    .reset(l1_idx_reset),
    .write_en(l1_idx_write_en)
);
std_add # (
    .WIDTH(4)
) l1_add (
    .left(l1_add_left),
    .out(l1_add_out),
    .right(l1_add_right)
);
std_reg # (
    .WIDTH(4)
) l2_idx (
    .clk(l2_idx_clk),
    .done(l2_idx_done),
    .in(l2_idx_in),
    .out(l2_idx_out),
    .reset(l2_idx_reset),
    .write_en(l2_idx_write_en)
);
std_add # (
    .WIDTH(4)
) l2_add (
    .left(l2_add_left),
    .out(l2_add_out),
    .right(l2_add_right)
);
std_reg # (
    .WIDTH(4)
) l3_idx (
    .clk(l3_idx_clk),
    .done(l3_idx_done),
    .in(l3_idx_in),
    .out(l3_idx_out),
    .reset(l3_idx_reset),
    .write_en(l3_idx_write_en)
);
std_add # (
    .WIDTH(4)
) l3_add (
    .left(l3_add_left),
    .out(l3_add_out),
    .right(l3_add_right)
);
std_reg # (
    .WIDTH(4)
) l4_idx (
    .clk(l4_idx_clk),
    .done(l4_idx_done),
    .in(l4_idx_in),
    .out(l4_idx_out),
    .reset(l4_idx_reset),
    .write_en(l4_idx_write_en)
);
std_add # (
    .WIDTH(4)
) l4_add (
    .left(l4_add_left),
    .out(l4_add_out),
    .right(l4_add_right)
);
std_reg # (
    .WIDTH(4)
) l5_idx (
    .clk(l5_idx_clk),
    .done(l5_idx_done),
    .in(l5_idx_in),
    .out(l5_idx_out),
    .reset(l5_idx_reset),
    .write_en(l5_idx_write_en)
);
std_add # (
    .WIDTH(4)
) l5_add (
    .left(l5_add_left),
    .out(l5_add_out),
    .right(l5_add_right)
);
std_reg # (
    .WIDTH(4)
) l6_idx (
    .clk(l6_idx_clk),
    .done(l6_idx_done),
    .in(l6_idx_in),
    .out(l6_idx_out),
    .reset(l6_idx_reset),
    .write_en(l6_idx_write_en)
);
std_add # (
    .WIDTH(4)
) l6_add (
    .left(l6_add_left),
    .out(l6_add_out),
    .right(l6_add_right)
);
std_reg # (
    .WIDTH(4)
) l7_idx (
    .clk(l7_idx_clk),
    .done(l7_idx_done),
    .in(l7_idx_in),
    .out(l7_idx_out),
    .reset(l7_idx_reset),
    .write_en(l7_idx_write_en)
);
std_add # (
    .WIDTH(4)
) l7_add (
    .left(l7_add_left),
    .out(l7_add_out),
    .right(l7_add_right)
);
std_reg # (
    .WIDTH(5)
) idx (
    .clk(idx_clk),
    .done(idx_done),
    .in(idx_in),
    .out(idx_out),
    .reset(idx_reset),
    .write_en(idx_write_en)
);
std_add # (
    .WIDTH(5)
) idx_add (
    .left(idx_add_left),
    .out(idx_add_out),
    .right(idx_add_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_18_26_reg (
    .clk(idx_between_18_26_reg_clk),
    .done(idx_between_18_26_reg_done),
    .in(idx_between_18_26_reg_in),
    .out(idx_between_18_26_reg_out),
    .reset(idx_between_18_26_reg_reset),
    .write_en(idx_between_18_26_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_26 (
    .left(index_lt_26_left),
    .out(index_lt_26_out),
    .right(index_lt_26_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_18 (
    .left(index_ge_18_left),
    .out(index_ge_18_out),
    .right(index_ge_18_right)
);
std_and # (
    .WIDTH(1)
) idx_between_18_26_comb (
    .left(idx_between_18_26_comb_left),
    .out(idx_between_18_26_comb_out),
    .right(idx_between_18_26_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_3_7_reg (
    .clk(idx_between_3_7_reg_clk),
    .done(idx_between_3_7_reg_done),
    .in(idx_between_3_7_reg_in),
    .out(idx_between_3_7_reg_out),
    .reset(idx_between_3_7_reg_reset),
    .write_en(idx_between_3_7_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_7 (
    .left(index_lt_7_left),
    .out(index_lt_7_out),
    .right(index_lt_7_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_3 (
    .left(index_ge_3_left),
    .out(index_ge_3_out),
    .right(index_ge_3_right)
);
std_and # (
    .WIDTH(1)
) idx_between_3_7_comb (
    .left(idx_between_3_7_comb_left),
    .out(idx_between_3_7_comb_out),
    .right(idx_between_3_7_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_12_16_reg (
    .clk(idx_between_12_16_reg_clk),
    .done(idx_between_12_16_reg_done),
    .in(idx_between_12_16_reg_in),
    .out(idx_between_12_16_reg_out),
    .reset(idx_between_12_16_reg_reset),
    .write_en(idx_between_12_16_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_16 (
    .left(index_lt_16_left),
    .out(index_lt_16_out),
    .right(index_lt_16_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_12 (
    .left(index_ge_12_left),
    .out(index_ge_12_out),
    .right(index_ge_12_right)
);
std_and # (
    .WIDTH(1)
) idx_between_12_16_comb (
    .left(idx_between_12_16_comb_left),
    .out(idx_between_12_16_comb_out),
    .right(idx_between_12_16_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_26_27_reg (
    .clk(idx_between_26_27_reg_clk),
    .done(idx_between_26_27_reg_done),
    .in(idx_between_26_27_reg_in),
    .out(idx_between_26_27_reg_out),
    .reset(idx_between_26_27_reg_reset),
    .write_en(idx_between_26_27_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_27 (
    .left(index_lt_27_left),
    .out(index_lt_27_out),
    .right(index_lt_27_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_26 (
    .left(index_ge_26_left),
    .out(index_ge_26_out),
    .right(index_ge_26_right)
);
std_and # (
    .WIDTH(1)
) idx_between_26_27_comb (
    .left(idx_between_26_27_comb_left),
    .out(idx_between_26_27_comb_out),
    .right(idx_between_26_27_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_4_12_reg (
    .clk(idx_between_4_12_reg_clk),
    .done(idx_between_4_12_reg_done),
    .in(idx_between_4_12_reg_in),
    .out(idx_between_4_12_reg_out),
    .reset(idx_between_4_12_reg_reset),
    .write_en(idx_between_4_12_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_12 (
    .left(index_lt_12_left),
    .out(index_lt_12_out),
    .right(index_lt_12_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_4 (
    .left(index_ge_4_left),
    .out(index_ge_4_out),
    .right(index_ge_4_right)
);
std_and # (
    .WIDTH(1)
) idx_between_4_12_comb (
    .left(idx_between_4_12_comb_left),
    .out(idx_between_4_12_comb_out),
    .right(idx_between_4_12_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_21_22_reg (
    .clk(idx_between_21_22_reg_clk),
    .done(idx_between_21_22_reg_done),
    .in(idx_between_21_22_reg_in),
    .out(idx_between_21_22_reg_out),
    .reset(idx_between_21_22_reg_reset),
    .write_en(idx_between_21_22_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_22 (
    .left(index_lt_22_left),
    .out(index_lt_22_out),
    .right(index_lt_22_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_21 (
    .left(index_ge_21_left),
    .out(index_ge_21_out),
    .right(index_ge_21_right)
);
std_and # (
    .WIDTH(1)
) idx_between_21_22_comb (
    .left(idx_between_21_22_comb_left),
    .out(idx_between_21_22_comb_out),
    .right(idx_between_21_22_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_5_13_reg (
    .clk(idx_between_5_13_reg_clk),
    .done(idx_between_5_13_reg_done),
    .in(idx_between_5_13_reg_in),
    .out(idx_between_5_13_reg_out),
    .reset(idx_between_5_13_reg_reset),
    .write_en(idx_between_5_13_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_13 (
    .left(index_lt_13_left),
    .out(index_lt_13_out),
    .right(index_lt_13_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_5 (
    .left(index_ge_5_left),
    .out(index_ge_5_out),
    .right(index_ge_5_right)
);
std_and # (
    .WIDTH(1)
) idx_between_5_13_comb (
    .left(idx_between_5_13_comb_left),
    .out(idx_between_5_13_comb_out),
    .right(idx_between_5_13_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_22_23_reg (
    .clk(idx_between_22_23_reg_clk),
    .done(idx_between_22_23_reg_done),
    .in(idx_between_22_23_reg_in),
    .out(idx_between_22_23_reg_out),
    .reset(idx_between_22_23_reg_reset),
    .write_en(idx_between_22_23_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_23 (
    .left(index_lt_23_left),
    .out(index_lt_23_out),
    .right(index_lt_23_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_22 (
    .left(index_ge_22_left),
    .out(index_ge_22_out),
    .right(index_ge_22_right)
);
std_and # (
    .WIDTH(1)
) idx_between_22_23_comb (
    .left(idx_between_22_23_comb_left),
    .out(idx_between_22_23_comb_out),
    .right(idx_between_22_23_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_14_22_reg (
    .clk(idx_between_14_22_reg_clk),
    .done(idx_between_14_22_reg_done),
    .in(idx_between_14_22_reg_in),
    .out(idx_between_14_22_reg_out),
    .reset(idx_between_14_22_reg_reset),
    .write_en(idx_between_14_22_reg_write_en)
);
std_ge # (
    .WIDTH(5)
) index_ge_14 (
    .left(index_ge_14_left),
    .out(index_ge_14_out),
    .right(index_ge_14_right)
);
std_and # (
    .WIDTH(1)
) idx_between_14_22_comb (
    .left(idx_between_14_22_comb_left),
    .out(idx_between_14_22_comb_out),
    .right(idx_between_14_22_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_8_12_reg (
    .clk(idx_between_8_12_reg_clk),
    .done(idx_between_8_12_reg_done),
    .in(idx_between_8_12_reg_in),
    .out(idx_between_8_12_reg_out),
    .reset(idx_between_8_12_reg_reset),
    .write_en(idx_between_8_12_reg_write_en)
);
std_ge # (
    .WIDTH(5)
) index_ge_8 (
    .left(index_ge_8_left),
    .out(index_ge_8_out),
    .right(index_ge_8_right)
);
std_and # (
    .WIDTH(1)
) idx_between_8_12_comb (
    .left(idx_between_8_12_comb_left),
    .out(idx_between_8_12_comb_out),
    .right(idx_between_8_12_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_9_17_reg (
    .clk(idx_between_9_17_reg_clk),
    .done(idx_between_9_17_reg_done),
    .in(idx_between_9_17_reg_in),
    .out(idx_between_9_17_reg_out),
    .reset(idx_between_9_17_reg_reset),
    .write_en(idx_between_9_17_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_17 (
    .left(index_lt_17_left),
    .out(index_lt_17_out),
    .right(index_lt_17_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_9 (
    .left(index_ge_9_left),
    .out(index_ge_9_out),
    .right(index_ge_9_right)
);
std_and # (
    .WIDTH(1)
) idx_between_9_17_comb (
    .left(idx_between_9_17_comb_left),
    .out(idx_between_9_17_comb_out),
    .right(idx_between_9_17_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_0_8_reg (
    .clk(idx_between_0_8_reg_clk),
    .done(idx_between_0_8_reg_done),
    .in(idx_between_0_8_reg_in),
    .out(idx_between_0_8_reg_out),
    .reset(idx_between_0_8_reg_reset),
    .write_en(idx_between_0_8_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_8 (
    .left(index_lt_8_left),
    .out(index_lt_8_out),
    .right(index_lt_8_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_17_18_reg (
    .clk(idx_between_17_18_reg_clk),
    .done(idx_between_17_18_reg_done),
    .in(idx_between_17_18_reg_in),
    .out(idx_between_17_18_reg_out),
    .reset(idx_between_17_18_reg_reset),
    .write_en(idx_between_17_18_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_18 (
    .left(index_lt_18_left),
    .out(index_lt_18_out),
    .right(index_lt_18_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_17 (
    .left(index_ge_17_left),
    .out(index_ge_17_out),
    .right(index_ge_17_right)
);
std_and # (
    .WIDTH(1)
) idx_between_17_18_comb (
    .left(idx_between_17_18_comb_left),
    .out(idx_between_17_18_comb_out),
    .right(idx_between_17_18_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_1_9_reg (
    .clk(idx_between_1_9_reg_clk),
    .done(idx_between_1_9_reg_done),
    .in(idx_between_1_9_reg_in),
    .out(idx_between_1_9_reg_out),
    .reset(idx_between_1_9_reg_reset),
    .write_en(idx_between_1_9_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_9 (
    .left(index_lt_9_left),
    .out(index_lt_9_out),
    .right(index_lt_9_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_1 (
    .left(index_ge_1_left),
    .out(index_ge_1_out),
    .right(index_ge_1_right)
);
std_and # (
    .WIDTH(1)
) idx_between_1_9_comb (
    .left(idx_between_1_9_comb_left),
    .out(idx_between_1_9_comb_out),
    .right(idx_between_1_9_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_10_18_reg (
    .clk(idx_between_10_18_reg_clk),
    .done(idx_between_10_18_reg_done),
    .in(idx_between_10_18_reg_in),
    .out(idx_between_10_18_reg_out),
    .reset(idx_between_10_18_reg_reset),
    .write_en(idx_between_10_18_reg_write_en)
);
std_ge # (
    .WIDTH(5)
) index_ge_10 (
    .left(index_ge_10_left),
    .out(index_ge_10_out),
    .right(index_ge_10_right)
);
std_and # (
    .WIDTH(1)
) idx_between_10_18_comb (
    .left(idx_between_10_18_comb_left),
    .out(idx_between_10_18_comb_out),
    .right(idx_between_10_18_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_25_26_reg (
    .clk(idx_between_25_26_reg_clk),
    .done(idx_between_25_26_reg_done),
    .in(idx_between_25_26_reg_in),
    .out(idx_between_25_26_reg_out),
    .reset(idx_between_25_26_reg_reset),
    .write_en(idx_between_25_26_reg_write_en)
);
std_ge # (
    .WIDTH(5)
) index_ge_25 (
    .left(index_ge_25_left),
    .out(index_ge_25_out),
    .right(index_ge_25_right)
);
std_and # (
    .WIDTH(1)
) idx_between_25_26_comb (
    .left(idx_between_25_26_comb_left),
    .out(idx_between_25_26_comb_out),
    .right(idx_between_25_26_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_27_28_reg (
    .clk(idx_between_27_28_reg_clk),
    .done(idx_between_27_28_reg_done),
    .in(idx_between_27_28_reg_in),
    .out(idx_between_27_28_reg_out),
    .reset(idx_between_27_28_reg_reset),
    .write_en(idx_between_27_28_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_28 (
    .left(index_lt_28_left),
    .out(index_lt_28_out),
    .right(index_lt_28_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_27 (
    .left(index_ge_27_left),
    .out(index_ge_27_out),
    .right(index_ge_27_right)
);
std_and # (
    .WIDTH(1)
) idx_between_27_28_comb (
    .left(idx_between_27_28_comb_left),
    .out(idx_between_27_28_comb_out),
    .right(idx_between_27_28_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_13_14_reg (
    .clk(idx_between_13_14_reg_clk),
    .done(idx_between_13_14_reg_done),
    .in(idx_between_13_14_reg_in),
    .out(idx_between_13_14_reg_out),
    .reset(idx_between_13_14_reg_reset),
    .write_en(idx_between_13_14_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_14 (
    .left(index_lt_14_left),
    .out(index_lt_14_out),
    .right(index_lt_14_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_13 (
    .left(index_ge_13_left),
    .out(index_ge_13_out),
    .right(index_ge_13_right)
);
std_and # (
    .WIDTH(1)
) idx_between_13_14_comb (
    .left(idx_between_13_14_comb_left),
    .out(idx_between_13_14_comb_out),
    .right(idx_between_13_14_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_19_27_reg (
    .clk(idx_between_19_27_reg_clk),
    .done(idx_between_19_27_reg_done),
    .in(idx_between_19_27_reg_in),
    .out(idx_between_19_27_reg_out),
    .reset(idx_between_19_27_reg_reset),
    .write_en(idx_between_19_27_reg_write_en)
);
std_ge # (
    .WIDTH(5)
) index_ge_19 (
    .left(index_ge_19_left),
    .out(index_ge_19_out),
    .right(index_ge_19_right)
);
std_and # (
    .WIDTH(1)
) idx_between_19_27_comb (
    .left(idx_between_19_27_comb_left),
    .out(idx_between_19_27_comb_out),
    .right(idx_between_19_27_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_13_17_reg (
    .clk(idx_between_13_17_reg_clk),
    .done(idx_between_13_17_reg_done),
    .in(idx_between_13_17_reg_in),
    .out(idx_between_13_17_reg_out),
    .reset(idx_between_13_17_reg_reset),
    .write_en(idx_between_13_17_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_13_17_comb (
    .left(idx_between_13_17_comb_left),
    .out(idx_between_13_17_comb_out),
    .right(idx_between_13_17_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_6_14_reg (
    .clk(idx_between_6_14_reg_clk),
    .done(idx_between_6_14_reg_done),
    .in(idx_between_6_14_reg_in),
    .out(idx_between_6_14_reg_out),
    .reset(idx_between_6_14_reg_reset),
    .write_en(idx_between_6_14_reg_write_en)
);
std_ge # (
    .WIDTH(5)
) index_ge_6 (
    .left(index_ge_6_left),
    .out(index_ge_6_out),
    .right(index_ge_6_right)
);
std_and # (
    .WIDTH(1)
) idx_between_6_14_comb (
    .left(idx_between_6_14_comb_left),
    .out(idx_between_6_14_comb_out),
    .right(idx_between_6_14_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_15_23_reg (
    .clk(idx_between_15_23_reg_clk),
    .done(idx_between_15_23_reg_done),
    .in(idx_between_15_23_reg_in),
    .out(idx_between_15_23_reg_out),
    .reset(idx_between_15_23_reg_reset),
    .write_en(idx_between_15_23_reg_write_en)
);
std_ge # (
    .WIDTH(5)
) index_ge_15 (
    .left(index_ge_15_left),
    .out(index_ge_15_out),
    .right(index_ge_15_right)
);
std_and # (
    .WIDTH(1)
) idx_between_15_23_comb (
    .left(idx_between_15_23_comb_left),
    .out(idx_between_15_23_comb_out),
    .right(idx_between_15_23_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_18_19_reg (
    .clk(idx_between_18_19_reg_clk),
    .done(idx_between_18_19_reg_done),
    .in(idx_between_18_19_reg_in),
    .out(idx_between_18_19_reg_out),
    .reset(idx_between_18_19_reg_reset),
    .write_en(idx_between_18_19_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_19 (
    .left(index_lt_19_left),
    .out(index_lt_19_out),
    .right(index_lt_19_right)
);
std_and # (
    .WIDTH(1)
) idx_between_18_19_comb (
    .left(idx_between_18_19_comb_left),
    .out(idx_between_18_19_comb_out),
    .right(idx_between_18_19_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_4_8_reg (
    .clk(idx_between_4_8_reg_clk),
    .done(idx_between_4_8_reg_done),
    .in(idx_between_4_8_reg_in),
    .out(idx_between_4_8_reg_out),
    .reset(idx_between_4_8_reg_reset),
    .write_en(idx_between_4_8_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_4_8_comb (
    .left(idx_between_4_8_comb_left),
    .out(idx_between_4_8_comb_out),
    .right(idx_between_4_8_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_5_9_reg (
    .clk(idx_between_5_9_reg_clk),
    .done(idx_between_5_9_reg_done),
    .in(idx_between_5_9_reg_in),
    .out(idx_between_5_9_reg_out),
    .reset(idx_between_5_9_reg_reset),
    .write_en(idx_between_5_9_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_5_9_comb (
    .left(idx_between_5_9_comb_left),
    .out(idx_between_5_9_comb_out),
    .right(idx_between_5_9_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_14_18_reg (
    .clk(idx_between_14_18_reg_clk),
    .done(idx_between_14_18_reg_done),
    .in(idx_between_14_18_reg_in),
    .out(idx_between_14_18_reg_out),
    .reset(idx_between_14_18_reg_reset),
    .write_en(idx_between_14_18_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_14_18_comb (
    .left(idx_between_14_18_comb_left),
    .out(idx_between_14_18_comb_out),
    .right(idx_between_14_18_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_14_15_reg (
    .clk(idx_between_14_15_reg_clk),
    .done(idx_between_14_15_reg_done),
    .in(idx_between_14_15_reg_in),
    .out(idx_between_14_15_reg_out),
    .reset(idx_between_14_15_reg_reset),
    .write_en(idx_between_14_15_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_15 (
    .left(index_lt_15_left),
    .out(index_lt_15_out),
    .right(index_lt_15_right)
);
std_and # (
    .WIDTH(1)
) idx_between_14_15_comb (
    .left(idx_between_14_15_comb_left),
    .out(idx_between_14_15_comb_out),
    .right(idx_between_14_15_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_23_24_reg (
    .clk(idx_between_23_24_reg_clk),
    .done(idx_between_23_24_reg_done),
    .in(idx_between_23_24_reg_in),
    .out(idx_between_23_24_reg_out),
    .reset(idx_between_23_24_reg_reset),
    .write_en(idx_between_23_24_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_24 (
    .left(index_lt_24_left),
    .out(index_lt_24_out),
    .right(index_lt_24_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_23 (
    .left(index_ge_23_left),
    .out(index_ge_23_out),
    .right(index_ge_23_right)
);
std_and # (
    .WIDTH(1)
) idx_between_23_24_comb (
    .left(idx_between_23_24_comb_left),
    .out(idx_between_23_24_comb_out),
    .right(idx_between_23_24_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_9_13_reg (
    .clk(idx_between_9_13_reg_clk),
    .done(idx_between_9_13_reg_done),
    .in(idx_between_9_13_reg_in),
    .out(idx_between_9_13_reg_out),
    .reset(idx_between_9_13_reg_reset),
    .write_en(idx_between_9_13_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_9_13_comb (
    .left(idx_between_9_13_comb_left),
    .out(idx_between_9_13_comb_out),
    .right(idx_between_9_13_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_1_5_reg (
    .clk(idx_between_1_5_reg_clk),
    .done(idx_between_1_5_reg_done),
    .in(idx_between_1_5_reg_in),
    .out(idx_between_1_5_reg_out),
    .reset(idx_between_1_5_reg_reset),
    .write_en(idx_between_1_5_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_5 (
    .left(index_lt_5_left),
    .out(index_lt_5_out),
    .right(index_lt_5_right)
);
std_and # (
    .WIDTH(1)
) idx_between_1_5_comb (
    .left(idx_between_1_5_comb_left),
    .out(idx_between_1_5_comb_out),
    .right(idx_between_1_5_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_10_14_reg (
    .clk(idx_between_10_14_reg_clk),
    .done(idx_between_10_14_reg_done),
    .in(idx_between_10_14_reg_in),
    .out(idx_between_10_14_reg_out),
    .reset(idx_between_10_14_reg_reset),
    .write_en(idx_between_10_14_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_10_14_comb (
    .left(idx_between_10_14_comb_left),
    .out(idx_between_10_14_comb_out),
    .right(idx_between_10_14_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_2_10_reg (
    .clk(idx_between_2_10_reg_clk),
    .done(idx_between_2_10_reg_done),
    .in(idx_between_2_10_reg_in),
    .out(idx_between_2_10_reg_out),
    .reset(idx_between_2_10_reg_reset),
    .write_en(idx_between_2_10_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_10 (
    .left(index_lt_10_left),
    .out(index_lt_10_out),
    .right(index_lt_10_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_2 (
    .left(index_ge_2_left),
    .out(index_ge_2_out),
    .right(index_ge_2_right)
);
std_and # (
    .WIDTH(1)
) idx_between_2_10_comb (
    .left(idx_between_2_10_comb_left),
    .out(idx_between_2_10_comb_out),
    .right(idx_between_2_10_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_11_19_reg (
    .clk(idx_between_11_19_reg_clk),
    .done(idx_between_11_19_reg_done),
    .in(idx_between_11_19_reg_in),
    .out(idx_between_11_19_reg_out),
    .reset(idx_between_11_19_reg_reset),
    .write_en(idx_between_11_19_reg_write_en)
);
std_ge # (
    .WIDTH(5)
) index_ge_11 (
    .left(index_ge_11_left),
    .out(index_ge_11_out),
    .right(index_ge_11_right)
);
std_and # (
    .WIDTH(1)
) idx_between_11_19_comb (
    .left(idx_between_11_19_comb_left),
    .out(idx_between_11_19_comb_out),
    .right(idx_between_11_19_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_19_20_reg (
    .clk(idx_between_19_20_reg_clk),
    .done(idx_between_19_20_reg_done),
    .in(idx_between_19_20_reg_in),
    .out(idx_between_19_20_reg_out),
    .reset(idx_between_19_20_reg_reset),
    .write_en(idx_between_19_20_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_20 (
    .left(index_lt_20_left),
    .out(index_lt_20_out),
    .right(index_lt_20_right)
);
std_and # (
    .WIDTH(1)
) idx_between_19_20_comb (
    .left(idx_between_19_20_comb_left),
    .out(idx_between_19_20_comb_out),
    .right(idx_between_19_20_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_15_16_reg (
    .clk(idx_between_15_16_reg_clk),
    .done(idx_between_15_16_reg_done),
    .in(idx_between_15_16_reg_in),
    .out(idx_between_15_16_reg_out),
    .reset(idx_between_15_16_reg_reset),
    .write_en(idx_between_15_16_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_15_16_comb (
    .left(idx_between_15_16_comb_left),
    .out(idx_between_15_16_comb_out),
    .right(idx_between_15_16_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_24_25_reg (
    .clk(idx_between_24_25_reg_clk),
    .done(idx_between_24_25_reg_done),
    .in(idx_between_24_25_reg_in),
    .out(idx_between_24_25_reg_out),
    .reset(idx_between_24_25_reg_reset),
    .write_en(idx_between_24_25_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_25 (
    .left(index_lt_25_left),
    .out(index_lt_25_out),
    .right(index_lt_25_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_24 (
    .left(index_ge_24_left),
    .out(index_ge_24_out),
    .right(index_ge_24_right)
);
std_and # (
    .WIDTH(1)
) idx_between_24_25_comb (
    .left(idx_between_24_25_comb_left),
    .out(idx_between_24_25_comb_out),
    .right(idx_between_24_25_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_6_10_reg (
    .clk(idx_between_6_10_reg_clk),
    .done(idx_between_6_10_reg_done),
    .in(idx_between_6_10_reg_in),
    .out(idx_between_6_10_reg_out),
    .reset(idx_between_6_10_reg_reset),
    .write_en(idx_between_6_10_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_6_10_comb (
    .left(idx_between_6_10_comb_left),
    .out(idx_between_6_10_comb_out),
    .right(idx_between_6_10_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_15_19_reg (
    .clk(idx_between_15_19_reg_clk),
    .done(idx_between_15_19_reg_done),
    .in(idx_between_15_19_reg_in),
    .out(idx_between_15_19_reg_out),
    .reset(idx_between_15_19_reg_reset),
    .write_en(idx_between_15_19_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_15_19_comb (
    .left(idx_between_15_19_comb_left),
    .out(idx_between_15_19_comb_out),
    .right(idx_between_15_19_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_7_15_reg (
    .clk(idx_between_7_15_reg_clk),
    .done(idx_between_7_15_reg_done),
    .in(idx_between_7_15_reg_in),
    .out(idx_between_7_15_reg_out),
    .reset(idx_between_7_15_reg_reset),
    .write_en(idx_between_7_15_reg_write_en)
);
std_ge # (
    .WIDTH(5)
) index_ge_7 (
    .left(index_ge_7_left),
    .out(index_ge_7_out),
    .right(index_ge_7_right)
);
std_and # (
    .WIDTH(1)
) idx_between_7_15_comb (
    .left(idx_between_7_15_comb_left),
    .out(idx_between_7_15_comb_out),
    .right(idx_between_7_15_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_16_24_reg (
    .clk(idx_between_16_24_reg_clk),
    .done(idx_between_16_24_reg_done),
    .in(idx_between_16_24_reg_in),
    .out(idx_between_16_24_reg_out),
    .reset(idx_between_16_24_reg_reset),
    .write_en(idx_between_16_24_reg_write_en)
);
std_ge # (
    .WIDTH(5)
) index_ge_16 (
    .left(index_ge_16_left),
    .out(index_ge_16_out),
    .right(index_ge_16_right)
);
std_and # (
    .WIDTH(1)
) idx_between_16_24_comb (
    .left(idx_between_16_24_comb_left),
    .out(idx_between_16_24_comb_out),
    .right(idx_between_16_24_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_3_11_reg (
    .clk(idx_between_3_11_reg_clk),
    .done(idx_between_3_11_reg_done),
    .in(idx_between_3_11_reg_in),
    .out(idx_between_3_11_reg_out),
    .reset(idx_between_3_11_reg_reset),
    .write_en(idx_between_3_11_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_11 (
    .left(index_lt_11_left),
    .out(index_lt_11_out),
    .right(index_lt_11_right)
);
std_and # (
    .WIDTH(1)
) idx_between_3_11_comb (
    .left(idx_between_3_11_comb_left),
    .out(idx_between_3_11_comb_out),
    .right(idx_between_3_11_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_20_21_reg (
    .clk(idx_between_20_21_reg_clk),
    .done(idx_between_20_21_reg_done),
    .in(idx_between_20_21_reg_in),
    .out(idx_between_20_21_reg_out),
    .reset(idx_between_20_21_reg_reset),
    .write_en(idx_between_20_21_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_21 (
    .left(index_lt_21_left),
    .out(index_lt_21_out),
    .right(index_lt_21_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_20 (
    .left(index_ge_20_left),
    .out(index_ge_20_out),
    .right(index_ge_20_right)
);
std_and # (
    .WIDTH(1)
) idx_between_20_21_comb (
    .left(idx_between_20_21_comb_left),
    .out(idx_between_20_21_comb_out),
    .right(idx_between_20_21_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_12_20_reg (
    .clk(idx_between_12_20_reg_clk),
    .done(idx_between_12_20_reg_done),
    .in(idx_between_12_20_reg_in),
    .out(idx_between_12_20_reg_out),
    .reset(idx_between_12_20_reg_reset),
    .write_en(idx_between_12_20_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_12_20_comb (
    .left(idx_between_12_20_comb_left),
    .out(idx_between_12_20_comb_out),
    .right(idx_between_12_20_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_8_16_reg (
    .clk(idx_between_8_16_reg_clk),
    .done(idx_between_8_16_reg_done),
    .in(idx_between_8_16_reg_in),
    .out(idx_between_8_16_reg_out),
    .reset(idx_between_8_16_reg_reset),
    .write_en(idx_between_8_16_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_8_16_comb (
    .left(idx_between_8_16_comb_left),
    .out(idx_between_8_16_comb_out),
    .right(idx_between_8_16_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_7_11_reg (
    .clk(idx_between_7_11_reg_clk),
    .done(idx_between_7_11_reg_done),
    .in(idx_between_7_11_reg_in),
    .out(idx_between_7_11_reg_out),
    .reset(idx_between_7_11_reg_reset),
    .write_en(idx_between_7_11_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_7_11_comb (
    .left(idx_between_7_11_comb_left),
    .out(idx_between_7_11_comb_out),
    .right(idx_between_7_11_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_2_6_reg (
    .clk(idx_between_2_6_reg_clk),
    .done(idx_between_2_6_reg_done),
    .in(idx_between_2_6_reg_in),
    .out(idx_between_2_6_reg_out),
    .reset(idx_between_2_6_reg_reset),
    .write_en(idx_between_2_6_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_6 (
    .left(index_lt_6_left),
    .out(index_lt_6_out),
    .right(index_lt_6_right)
);
std_and # (
    .WIDTH(1)
) idx_between_2_6_comb (
    .left(idx_between_2_6_comb_left),
    .out(idx_between_2_6_comb_out),
    .right(idx_between_2_6_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_11_15_reg (
    .clk(idx_between_11_15_reg_clk),
    .done(idx_between_11_15_reg_done),
    .in(idx_between_11_15_reg_in),
    .out(idx_between_11_15_reg_out),
    .reset(idx_between_11_15_reg_reset),
    .write_en(idx_between_11_15_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_11_15_comb (
    .left(idx_between_11_15_comb_left),
    .out(idx_between_11_15_comb_out),
    .right(idx_between_11_15_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_17_25_reg (
    .clk(idx_between_17_25_reg_clk),
    .done(idx_between_17_25_reg_done),
    .in(idx_between_17_25_reg_in),
    .out(idx_between_17_25_reg_out),
    .reset(idx_between_17_25_reg_reset),
    .write_en(idx_between_17_25_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_17_25_comb (
    .left(idx_between_17_25_comb_left),
    .out(idx_between_17_25_comb_out),
    .right(idx_between_17_25_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_13_21_reg (
    .clk(idx_between_13_21_reg_clk),
    .done(idx_between_13_21_reg_done),
    .in(idx_between_13_21_reg_in),
    .out(idx_between_13_21_reg_out),
    .reset(idx_between_13_21_reg_reset),
    .write_en(idx_between_13_21_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_13_21_comb (
    .left(idx_between_13_21_comb_left),
    .out(idx_between_13_21_comb_out),
    .right(idx_between_13_21_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_16_17_reg (
    .clk(idx_between_16_17_reg_clk),
    .done(idx_between_16_17_reg_done),
    .in(idx_between_16_17_reg_in),
    .out(idx_between_16_17_reg_out),
    .reset(idx_between_16_17_reg_reset),
    .write_en(idx_between_16_17_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_16_17_comb (
    .left(idx_between_16_17_comb_left),
    .out(idx_between_16_17_comb_out),
    .right(idx_between_16_17_comb_right)
);
std_reg # (
    .WIDTH(1)
) cond (
    .clk(cond_clk),
    .done(cond_done),
    .in(cond_in),
    .out(cond_out),
    .reset(cond_reset),
    .write_en(cond_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire (
    .in(cond_wire_in),
    .out(cond_wire_out)
);
std_reg # (
    .WIDTH(1)
) cond0 (
    .clk(cond0_clk),
    .done(cond0_done),
    .in(cond0_in),
    .out(cond0_out),
    .reset(cond0_reset),
    .write_en(cond0_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire0 (
    .in(cond_wire0_in),
    .out(cond_wire0_out)
);
std_reg # (
    .WIDTH(1)
) cond1 (
    .clk(cond1_clk),
    .done(cond1_done),
    .in(cond1_in),
    .out(cond1_out),
    .reset(cond1_reset),
    .write_en(cond1_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1 (
    .in(cond_wire1_in),
    .out(cond_wire1_out)
);
std_reg # (
    .WIDTH(1)
) cond2 (
    .clk(cond2_clk),
    .done(cond2_done),
    .in(cond2_in),
    .out(cond2_out),
    .reset(cond2_reset),
    .write_en(cond2_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire2 (
    .in(cond_wire2_in),
    .out(cond_wire2_out)
);
std_reg # (
    .WIDTH(1)
) cond3 (
    .clk(cond3_clk),
    .done(cond3_done),
    .in(cond3_in),
    .out(cond3_out),
    .reset(cond3_reset),
    .write_en(cond3_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire3 (
    .in(cond_wire3_in),
    .out(cond_wire3_out)
);
std_reg # (
    .WIDTH(1)
) cond4 (
    .clk(cond4_clk),
    .done(cond4_done),
    .in(cond4_in),
    .out(cond4_out),
    .reset(cond4_reset),
    .write_en(cond4_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire4 (
    .in(cond_wire4_in),
    .out(cond_wire4_out)
);
std_reg # (
    .WIDTH(1)
) cond5 (
    .clk(cond5_clk),
    .done(cond5_done),
    .in(cond5_in),
    .out(cond5_out),
    .reset(cond5_reset),
    .write_en(cond5_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire5 (
    .in(cond_wire5_in),
    .out(cond_wire5_out)
);
std_reg # (
    .WIDTH(1)
) cond6 (
    .clk(cond6_clk),
    .done(cond6_done),
    .in(cond6_in),
    .out(cond6_out),
    .reset(cond6_reset),
    .write_en(cond6_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire6 (
    .in(cond_wire6_in),
    .out(cond_wire6_out)
);
std_reg # (
    .WIDTH(1)
) cond7 (
    .clk(cond7_clk),
    .done(cond7_done),
    .in(cond7_in),
    .out(cond7_out),
    .reset(cond7_reset),
    .write_en(cond7_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire7 (
    .in(cond_wire7_in),
    .out(cond_wire7_out)
);
std_reg # (
    .WIDTH(1)
) cond8 (
    .clk(cond8_clk),
    .done(cond8_done),
    .in(cond8_in),
    .out(cond8_out),
    .reset(cond8_reset),
    .write_en(cond8_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire8 (
    .in(cond_wire8_in),
    .out(cond_wire8_out)
);
std_reg # (
    .WIDTH(1)
) cond9 (
    .clk(cond9_clk),
    .done(cond9_done),
    .in(cond9_in),
    .out(cond9_out),
    .reset(cond9_reset),
    .write_en(cond9_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire9 (
    .in(cond_wire9_in),
    .out(cond_wire9_out)
);
std_reg # (
    .WIDTH(1)
) cond10 (
    .clk(cond10_clk),
    .done(cond10_done),
    .in(cond10_in),
    .out(cond10_out),
    .reset(cond10_reset),
    .write_en(cond10_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire10 (
    .in(cond_wire10_in),
    .out(cond_wire10_out)
);
std_reg # (
    .WIDTH(1)
) cond11 (
    .clk(cond11_clk),
    .done(cond11_done),
    .in(cond11_in),
    .out(cond11_out),
    .reset(cond11_reset),
    .write_en(cond11_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire11 (
    .in(cond_wire11_in),
    .out(cond_wire11_out)
);
std_reg # (
    .WIDTH(1)
) cond12 (
    .clk(cond12_clk),
    .done(cond12_done),
    .in(cond12_in),
    .out(cond12_out),
    .reset(cond12_reset),
    .write_en(cond12_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire12 (
    .in(cond_wire12_in),
    .out(cond_wire12_out)
);
std_reg # (
    .WIDTH(1)
) cond13 (
    .clk(cond13_clk),
    .done(cond13_done),
    .in(cond13_in),
    .out(cond13_out),
    .reset(cond13_reset),
    .write_en(cond13_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire13 (
    .in(cond_wire13_in),
    .out(cond_wire13_out)
);
std_reg # (
    .WIDTH(1)
) cond14 (
    .clk(cond14_clk),
    .done(cond14_done),
    .in(cond14_in),
    .out(cond14_out),
    .reset(cond14_reset),
    .write_en(cond14_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire14 (
    .in(cond_wire14_in),
    .out(cond_wire14_out)
);
std_reg # (
    .WIDTH(1)
) cond15 (
    .clk(cond15_clk),
    .done(cond15_done),
    .in(cond15_in),
    .out(cond15_out),
    .reset(cond15_reset),
    .write_en(cond15_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire15 (
    .in(cond_wire15_in),
    .out(cond_wire15_out)
);
std_reg # (
    .WIDTH(1)
) cond16 (
    .clk(cond16_clk),
    .done(cond16_done),
    .in(cond16_in),
    .out(cond16_out),
    .reset(cond16_reset),
    .write_en(cond16_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire16 (
    .in(cond_wire16_in),
    .out(cond_wire16_out)
);
std_reg # (
    .WIDTH(1)
) cond17 (
    .clk(cond17_clk),
    .done(cond17_done),
    .in(cond17_in),
    .out(cond17_out),
    .reset(cond17_reset),
    .write_en(cond17_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire17 (
    .in(cond_wire17_in),
    .out(cond_wire17_out)
);
std_reg # (
    .WIDTH(1)
) cond18 (
    .clk(cond18_clk),
    .done(cond18_done),
    .in(cond18_in),
    .out(cond18_out),
    .reset(cond18_reset),
    .write_en(cond18_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire18 (
    .in(cond_wire18_in),
    .out(cond_wire18_out)
);
std_reg # (
    .WIDTH(1)
) cond19 (
    .clk(cond19_clk),
    .done(cond19_done),
    .in(cond19_in),
    .out(cond19_out),
    .reset(cond19_reset),
    .write_en(cond19_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire19 (
    .in(cond_wire19_in),
    .out(cond_wire19_out)
);
std_reg # (
    .WIDTH(1)
) cond20 (
    .clk(cond20_clk),
    .done(cond20_done),
    .in(cond20_in),
    .out(cond20_out),
    .reset(cond20_reset),
    .write_en(cond20_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire20 (
    .in(cond_wire20_in),
    .out(cond_wire20_out)
);
std_reg # (
    .WIDTH(1)
) cond21 (
    .clk(cond21_clk),
    .done(cond21_done),
    .in(cond21_in),
    .out(cond21_out),
    .reset(cond21_reset),
    .write_en(cond21_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire21 (
    .in(cond_wire21_in),
    .out(cond_wire21_out)
);
std_reg # (
    .WIDTH(1)
) cond22 (
    .clk(cond22_clk),
    .done(cond22_done),
    .in(cond22_in),
    .out(cond22_out),
    .reset(cond22_reset),
    .write_en(cond22_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire22 (
    .in(cond_wire22_in),
    .out(cond_wire22_out)
);
std_reg # (
    .WIDTH(1)
) cond23 (
    .clk(cond23_clk),
    .done(cond23_done),
    .in(cond23_in),
    .out(cond23_out),
    .reset(cond23_reset),
    .write_en(cond23_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire23 (
    .in(cond_wire23_in),
    .out(cond_wire23_out)
);
std_reg # (
    .WIDTH(1)
) cond24 (
    .clk(cond24_clk),
    .done(cond24_done),
    .in(cond24_in),
    .out(cond24_out),
    .reset(cond24_reset),
    .write_en(cond24_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire24 (
    .in(cond_wire24_in),
    .out(cond_wire24_out)
);
std_reg # (
    .WIDTH(1)
) cond25 (
    .clk(cond25_clk),
    .done(cond25_done),
    .in(cond25_in),
    .out(cond25_out),
    .reset(cond25_reset),
    .write_en(cond25_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire25 (
    .in(cond_wire25_in),
    .out(cond_wire25_out)
);
std_reg # (
    .WIDTH(1)
) cond26 (
    .clk(cond26_clk),
    .done(cond26_done),
    .in(cond26_in),
    .out(cond26_out),
    .reset(cond26_reset),
    .write_en(cond26_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire26 (
    .in(cond_wire26_in),
    .out(cond_wire26_out)
);
std_reg # (
    .WIDTH(1)
) cond27 (
    .clk(cond27_clk),
    .done(cond27_done),
    .in(cond27_in),
    .out(cond27_out),
    .reset(cond27_reset),
    .write_en(cond27_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire27 (
    .in(cond_wire27_in),
    .out(cond_wire27_out)
);
std_reg # (
    .WIDTH(1)
) cond28 (
    .clk(cond28_clk),
    .done(cond28_done),
    .in(cond28_in),
    .out(cond28_out),
    .reset(cond28_reset),
    .write_en(cond28_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire28 (
    .in(cond_wire28_in),
    .out(cond_wire28_out)
);
std_reg # (
    .WIDTH(1)
) cond29 (
    .clk(cond29_clk),
    .done(cond29_done),
    .in(cond29_in),
    .out(cond29_out),
    .reset(cond29_reset),
    .write_en(cond29_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire29 (
    .in(cond_wire29_in),
    .out(cond_wire29_out)
);
std_reg # (
    .WIDTH(1)
) cond30 (
    .clk(cond30_clk),
    .done(cond30_done),
    .in(cond30_in),
    .out(cond30_out),
    .reset(cond30_reset),
    .write_en(cond30_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire30 (
    .in(cond_wire30_in),
    .out(cond_wire30_out)
);
std_reg # (
    .WIDTH(1)
) cond31 (
    .clk(cond31_clk),
    .done(cond31_done),
    .in(cond31_in),
    .out(cond31_out),
    .reset(cond31_reset),
    .write_en(cond31_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire31 (
    .in(cond_wire31_in),
    .out(cond_wire31_out)
);
std_reg # (
    .WIDTH(1)
) cond32 (
    .clk(cond32_clk),
    .done(cond32_done),
    .in(cond32_in),
    .out(cond32_out),
    .reset(cond32_reset),
    .write_en(cond32_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire32 (
    .in(cond_wire32_in),
    .out(cond_wire32_out)
);
std_reg # (
    .WIDTH(1)
) cond33 (
    .clk(cond33_clk),
    .done(cond33_done),
    .in(cond33_in),
    .out(cond33_out),
    .reset(cond33_reset),
    .write_en(cond33_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire33 (
    .in(cond_wire33_in),
    .out(cond_wire33_out)
);
std_reg # (
    .WIDTH(1)
) cond34 (
    .clk(cond34_clk),
    .done(cond34_done),
    .in(cond34_in),
    .out(cond34_out),
    .reset(cond34_reset),
    .write_en(cond34_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire34 (
    .in(cond_wire34_in),
    .out(cond_wire34_out)
);
std_reg # (
    .WIDTH(1)
) cond35 (
    .clk(cond35_clk),
    .done(cond35_done),
    .in(cond35_in),
    .out(cond35_out),
    .reset(cond35_reset),
    .write_en(cond35_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire35 (
    .in(cond_wire35_in),
    .out(cond_wire35_out)
);
std_reg # (
    .WIDTH(1)
) cond36 (
    .clk(cond36_clk),
    .done(cond36_done),
    .in(cond36_in),
    .out(cond36_out),
    .reset(cond36_reset),
    .write_en(cond36_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire36 (
    .in(cond_wire36_in),
    .out(cond_wire36_out)
);
std_reg # (
    .WIDTH(1)
) cond37 (
    .clk(cond37_clk),
    .done(cond37_done),
    .in(cond37_in),
    .out(cond37_out),
    .reset(cond37_reset),
    .write_en(cond37_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire37 (
    .in(cond_wire37_in),
    .out(cond_wire37_out)
);
std_reg # (
    .WIDTH(1)
) cond38 (
    .clk(cond38_clk),
    .done(cond38_done),
    .in(cond38_in),
    .out(cond38_out),
    .reset(cond38_reset),
    .write_en(cond38_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire38 (
    .in(cond_wire38_in),
    .out(cond_wire38_out)
);
std_reg # (
    .WIDTH(1)
) cond39 (
    .clk(cond39_clk),
    .done(cond39_done),
    .in(cond39_in),
    .out(cond39_out),
    .reset(cond39_reset),
    .write_en(cond39_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire39 (
    .in(cond_wire39_in),
    .out(cond_wire39_out)
);
std_reg # (
    .WIDTH(1)
) cond40 (
    .clk(cond40_clk),
    .done(cond40_done),
    .in(cond40_in),
    .out(cond40_out),
    .reset(cond40_reset),
    .write_en(cond40_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire40 (
    .in(cond_wire40_in),
    .out(cond_wire40_out)
);
std_reg # (
    .WIDTH(1)
) cond41 (
    .clk(cond41_clk),
    .done(cond41_done),
    .in(cond41_in),
    .out(cond41_out),
    .reset(cond41_reset),
    .write_en(cond41_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire41 (
    .in(cond_wire41_in),
    .out(cond_wire41_out)
);
std_reg # (
    .WIDTH(1)
) cond42 (
    .clk(cond42_clk),
    .done(cond42_done),
    .in(cond42_in),
    .out(cond42_out),
    .reset(cond42_reset),
    .write_en(cond42_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire42 (
    .in(cond_wire42_in),
    .out(cond_wire42_out)
);
std_reg # (
    .WIDTH(1)
) cond43 (
    .clk(cond43_clk),
    .done(cond43_done),
    .in(cond43_in),
    .out(cond43_out),
    .reset(cond43_reset),
    .write_en(cond43_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire43 (
    .in(cond_wire43_in),
    .out(cond_wire43_out)
);
std_reg # (
    .WIDTH(1)
) cond44 (
    .clk(cond44_clk),
    .done(cond44_done),
    .in(cond44_in),
    .out(cond44_out),
    .reset(cond44_reset),
    .write_en(cond44_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire44 (
    .in(cond_wire44_in),
    .out(cond_wire44_out)
);
std_reg # (
    .WIDTH(1)
) cond45 (
    .clk(cond45_clk),
    .done(cond45_done),
    .in(cond45_in),
    .out(cond45_out),
    .reset(cond45_reset),
    .write_en(cond45_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire45 (
    .in(cond_wire45_in),
    .out(cond_wire45_out)
);
std_reg # (
    .WIDTH(1)
) cond46 (
    .clk(cond46_clk),
    .done(cond46_done),
    .in(cond46_in),
    .out(cond46_out),
    .reset(cond46_reset),
    .write_en(cond46_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire46 (
    .in(cond_wire46_in),
    .out(cond_wire46_out)
);
std_reg # (
    .WIDTH(1)
) cond47 (
    .clk(cond47_clk),
    .done(cond47_done),
    .in(cond47_in),
    .out(cond47_out),
    .reset(cond47_reset),
    .write_en(cond47_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire47 (
    .in(cond_wire47_in),
    .out(cond_wire47_out)
);
std_reg # (
    .WIDTH(1)
) cond48 (
    .clk(cond48_clk),
    .done(cond48_done),
    .in(cond48_in),
    .out(cond48_out),
    .reset(cond48_reset),
    .write_en(cond48_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire48 (
    .in(cond_wire48_in),
    .out(cond_wire48_out)
);
std_reg # (
    .WIDTH(1)
) cond49 (
    .clk(cond49_clk),
    .done(cond49_done),
    .in(cond49_in),
    .out(cond49_out),
    .reset(cond49_reset),
    .write_en(cond49_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire49 (
    .in(cond_wire49_in),
    .out(cond_wire49_out)
);
std_reg # (
    .WIDTH(1)
) cond50 (
    .clk(cond50_clk),
    .done(cond50_done),
    .in(cond50_in),
    .out(cond50_out),
    .reset(cond50_reset),
    .write_en(cond50_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire50 (
    .in(cond_wire50_in),
    .out(cond_wire50_out)
);
std_reg # (
    .WIDTH(1)
) cond51 (
    .clk(cond51_clk),
    .done(cond51_done),
    .in(cond51_in),
    .out(cond51_out),
    .reset(cond51_reset),
    .write_en(cond51_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire51 (
    .in(cond_wire51_in),
    .out(cond_wire51_out)
);
std_reg # (
    .WIDTH(1)
) cond52 (
    .clk(cond52_clk),
    .done(cond52_done),
    .in(cond52_in),
    .out(cond52_out),
    .reset(cond52_reset),
    .write_en(cond52_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire52 (
    .in(cond_wire52_in),
    .out(cond_wire52_out)
);
std_reg # (
    .WIDTH(1)
) cond53 (
    .clk(cond53_clk),
    .done(cond53_done),
    .in(cond53_in),
    .out(cond53_out),
    .reset(cond53_reset),
    .write_en(cond53_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire53 (
    .in(cond_wire53_in),
    .out(cond_wire53_out)
);
std_reg # (
    .WIDTH(1)
) cond54 (
    .clk(cond54_clk),
    .done(cond54_done),
    .in(cond54_in),
    .out(cond54_out),
    .reset(cond54_reset),
    .write_en(cond54_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire54 (
    .in(cond_wire54_in),
    .out(cond_wire54_out)
);
std_reg # (
    .WIDTH(1)
) cond55 (
    .clk(cond55_clk),
    .done(cond55_done),
    .in(cond55_in),
    .out(cond55_out),
    .reset(cond55_reset),
    .write_en(cond55_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire55 (
    .in(cond_wire55_in),
    .out(cond_wire55_out)
);
std_reg # (
    .WIDTH(1)
) cond56 (
    .clk(cond56_clk),
    .done(cond56_done),
    .in(cond56_in),
    .out(cond56_out),
    .reset(cond56_reset),
    .write_en(cond56_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire56 (
    .in(cond_wire56_in),
    .out(cond_wire56_out)
);
std_reg # (
    .WIDTH(1)
) cond57 (
    .clk(cond57_clk),
    .done(cond57_done),
    .in(cond57_in),
    .out(cond57_out),
    .reset(cond57_reset),
    .write_en(cond57_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire57 (
    .in(cond_wire57_in),
    .out(cond_wire57_out)
);
std_reg # (
    .WIDTH(1)
) cond58 (
    .clk(cond58_clk),
    .done(cond58_done),
    .in(cond58_in),
    .out(cond58_out),
    .reset(cond58_reset),
    .write_en(cond58_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire58 (
    .in(cond_wire58_in),
    .out(cond_wire58_out)
);
std_reg # (
    .WIDTH(1)
) cond59 (
    .clk(cond59_clk),
    .done(cond59_done),
    .in(cond59_in),
    .out(cond59_out),
    .reset(cond59_reset),
    .write_en(cond59_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire59 (
    .in(cond_wire59_in),
    .out(cond_wire59_out)
);
std_reg # (
    .WIDTH(1)
) cond60 (
    .clk(cond60_clk),
    .done(cond60_done),
    .in(cond60_in),
    .out(cond60_out),
    .reset(cond60_reset),
    .write_en(cond60_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire60 (
    .in(cond_wire60_in),
    .out(cond_wire60_out)
);
std_reg # (
    .WIDTH(1)
) cond61 (
    .clk(cond61_clk),
    .done(cond61_done),
    .in(cond61_in),
    .out(cond61_out),
    .reset(cond61_reset),
    .write_en(cond61_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire61 (
    .in(cond_wire61_in),
    .out(cond_wire61_out)
);
std_reg # (
    .WIDTH(1)
) cond62 (
    .clk(cond62_clk),
    .done(cond62_done),
    .in(cond62_in),
    .out(cond62_out),
    .reset(cond62_reset),
    .write_en(cond62_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire62 (
    .in(cond_wire62_in),
    .out(cond_wire62_out)
);
std_reg # (
    .WIDTH(1)
) cond63 (
    .clk(cond63_clk),
    .done(cond63_done),
    .in(cond63_in),
    .out(cond63_out),
    .reset(cond63_reset),
    .write_en(cond63_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire63 (
    .in(cond_wire63_in),
    .out(cond_wire63_out)
);
std_reg # (
    .WIDTH(1)
) cond64 (
    .clk(cond64_clk),
    .done(cond64_done),
    .in(cond64_in),
    .out(cond64_out),
    .reset(cond64_reset),
    .write_en(cond64_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire64 (
    .in(cond_wire64_in),
    .out(cond_wire64_out)
);
std_reg # (
    .WIDTH(1)
) cond65 (
    .clk(cond65_clk),
    .done(cond65_done),
    .in(cond65_in),
    .out(cond65_out),
    .reset(cond65_reset),
    .write_en(cond65_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire65 (
    .in(cond_wire65_in),
    .out(cond_wire65_out)
);
std_reg # (
    .WIDTH(1)
) cond66 (
    .clk(cond66_clk),
    .done(cond66_done),
    .in(cond66_in),
    .out(cond66_out),
    .reset(cond66_reset),
    .write_en(cond66_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire66 (
    .in(cond_wire66_in),
    .out(cond_wire66_out)
);
std_reg # (
    .WIDTH(1)
) cond67 (
    .clk(cond67_clk),
    .done(cond67_done),
    .in(cond67_in),
    .out(cond67_out),
    .reset(cond67_reset),
    .write_en(cond67_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire67 (
    .in(cond_wire67_in),
    .out(cond_wire67_out)
);
std_reg # (
    .WIDTH(1)
) cond68 (
    .clk(cond68_clk),
    .done(cond68_done),
    .in(cond68_in),
    .out(cond68_out),
    .reset(cond68_reset),
    .write_en(cond68_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire68 (
    .in(cond_wire68_in),
    .out(cond_wire68_out)
);
std_reg # (
    .WIDTH(1)
) cond69 (
    .clk(cond69_clk),
    .done(cond69_done),
    .in(cond69_in),
    .out(cond69_out),
    .reset(cond69_reset),
    .write_en(cond69_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire69 (
    .in(cond_wire69_in),
    .out(cond_wire69_out)
);
std_reg # (
    .WIDTH(1)
) cond70 (
    .clk(cond70_clk),
    .done(cond70_done),
    .in(cond70_in),
    .out(cond70_out),
    .reset(cond70_reset),
    .write_en(cond70_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire70 (
    .in(cond_wire70_in),
    .out(cond_wire70_out)
);
std_reg # (
    .WIDTH(1)
) cond71 (
    .clk(cond71_clk),
    .done(cond71_done),
    .in(cond71_in),
    .out(cond71_out),
    .reset(cond71_reset),
    .write_en(cond71_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire71 (
    .in(cond_wire71_in),
    .out(cond_wire71_out)
);
std_reg # (
    .WIDTH(1)
) cond72 (
    .clk(cond72_clk),
    .done(cond72_done),
    .in(cond72_in),
    .out(cond72_out),
    .reset(cond72_reset),
    .write_en(cond72_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire72 (
    .in(cond_wire72_in),
    .out(cond_wire72_out)
);
std_reg # (
    .WIDTH(1)
) cond73 (
    .clk(cond73_clk),
    .done(cond73_done),
    .in(cond73_in),
    .out(cond73_out),
    .reset(cond73_reset),
    .write_en(cond73_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire73 (
    .in(cond_wire73_in),
    .out(cond_wire73_out)
);
std_reg # (
    .WIDTH(1)
) cond74 (
    .clk(cond74_clk),
    .done(cond74_done),
    .in(cond74_in),
    .out(cond74_out),
    .reset(cond74_reset),
    .write_en(cond74_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire74 (
    .in(cond_wire74_in),
    .out(cond_wire74_out)
);
std_reg # (
    .WIDTH(1)
) cond75 (
    .clk(cond75_clk),
    .done(cond75_done),
    .in(cond75_in),
    .out(cond75_out),
    .reset(cond75_reset),
    .write_en(cond75_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire75 (
    .in(cond_wire75_in),
    .out(cond_wire75_out)
);
std_reg # (
    .WIDTH(1)
) cond76 (
    .clk(cond76_clk),
    .done(cond76_done),
    .in(cond76_in),
    .out(cond76_out),
    .reset(cond76_reset),
    .write_en(cond76_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire76 (
    .in(cond_wire76_in),
    .out(cond_wire76_out)
);
std_reg # (
    .WIDTH(1)
) cond77 (
    .clk(cond77_clk),
    .done(cond77_done),
    .in(cond77_in),
    .out(cond77_out),
    .reset(cond77_reset),
    .write_en(cond77_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire77 (
    .in(cond_wire77_in),
    .out(cond_wire77_out)
);
std_reg # (
    .WIDTH(1)
) cond78 (
    .clk(cond78_clk),
    .done(cond78_done),
    .in(cond78_in),
    .out(cond78_out),
    .reset(cond78_reset),
    .write_en(cond78_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire78 (
    .in(cond_wire78_in),
    .out(cond_wire78_out)
);
std_reg # (
    .WIDTH(1)
) cond79 (
    .clk(cond79_clk),
    .done(cond79_done),
    .in(cond79_in),
    .out(cond79_out),
    .reset(cond79_reset),
    .write_en(cond79_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire79 (
    .in(cond_wire79_in),
    .out(cond_wire79_out)
);
std_reg # (
    .WIDTH(1)
) cond80 (
    .clk(cond80_clk),
    .done(cond80_done),
    .in(cond80_in),
    .out(cond80_out),
    .reset(cond80_reset),
    .write_en(cond80_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire80 (
    .in(cond_wire80_in),
    .out(cond_wire80_out)
);
std_reg # (
    .WIDTH(1)
) cond81 (
    .clk(cond81_clk),
    .done(cond81_done),
    .in(cond81_in),
    .out(cond81_out),
    .reset(cond81_reset),
    .write_en(cond81_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire81 (
    .in(cond_wire81_in),
    .out(cond_wire81_out)
);
std_reg # (
    .WIDTH(1)
) cond82 (
    .clk(cond82_clk),
    .done(cond82_done),
    .in(cond82_in),
    .out(cond82_out),
    .reset(cond82_reset),
    .write_en(cond82_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire82 (
    .in(cond_wire82_in),
    .out(cond_wire82_out)
);
std_reg # (
    .WIDTH(1)
) cond83 (
    .clk(cond83_clk),
    .done(cond83_done),
    .in(cond83_in),
    .out(cond83_out),
    .reset(cond83_reset),
    .write_en(cond83_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire83 (
    .in(cond_wire83_in),
    .out(cond_wire83_out)
);
std_reg # (
    .WIDTH(1)
) cond84 (
    .clk(cond84_clk),
    .done(cond84_done),
    .in(cond84_in),
    .out(cond84_out),
    .reset(cond84_reset),
    .write_en(cond84_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire84 (
    .in(cond_wire84_in),
    .out(cond_wire84_out)
);
std_reg # (
    .WIDTH(1)
) cond85 (
    .clk(cond85_clk),
    .done(cond85_done),
    .in(cond85_in),
    .out(cond85_out),
    .reset(cond85_reset),
    .write_en(cond85_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire85 (
    .in(cond_wire85_in),
    .out(cond_wire85_out)
);
std_reg # (
    .WIDTH(1)
) cond86 (
    .clk(cond86_clk),
    .done(cond86_done),
    .in(cond86_in),
    .out(cond86_out),
    .reset(cond86_reset),
    .write_en(cond86_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire86 (
    .in(cond_wire86_in),
    .out(cond_wire86_out)
);
std_reg # (
    .WIDTH(1)
) cond87 (
    .clk(cond87_clk),
    .done(cond87_done),
    .in(cond87_in),
    .out(cond87_out),
    .reset(cond87_reset),
    .write_en(cond87_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire87 (
    .in(cond_wire87_in),
    .out(cond_wire87_out)
);
std_reg # (
    .WIDTH(1)
) cond88 (
    .clk(cond88_clk),
    .done(cond88_done),
    .in(cond88_in),
    .out(cond88_out),
    .reset(cond88_reset),
    .write_en(cond88_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire88 (
    .in(cond_wire88_in),
    .out(cond_wire88_out)
);
std_reg # (
    .WIDTH(1)
) cond89 (
    .clk(cond89_clk),
    .done(cond89_done),
    .in(cond89_in),
    .out(cond89_out),
    .reset(cond89_reset),
    .write_en(cond89_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire89 (
    .in(cond_wire89_in),
    .out(cond_wire89_out)
);
std_reg # (
    .WIDTH(1)
) cond90 (
    .clk(cond90_clk),
    .done(cond90_done),
    .in(cond90_in),
    .out(cond90_out),
    .reset(cond90_reset),
    .write_en(cond90_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire90 (
    .in(cond_wire90_in),
    .out(cond_wire90_out)
);
std_reg # (
    .WIDTH(1)
) cond91 (
    .clk(cond91_clk),
    .done(cond91_done),
    .in(cond91_in),
    .out(cond91_out),
    .reset(cond91_reset),
    .write_en(cond91_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire91 (
    .in(cond_wire91_in),
    .out(cond_wire91_out)
);
std_reg # (
    .WIDTH(1)
) cond92 (
    .clk(cond92_clk),
    .done(cond92_done),
    .in(cond92_in),
    .out(cond92_out),
    .reset(cond92_reset),
    .write_en(cond92_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire92 (
    .in(cond_wire92_in),
    .out(cond_wire92_out)
);
std_reg # (
    .WIDTH(1)
) cond93 (
    .clk(cond93_clk),
    .done(cond93_done),
    .in(cond93_in),
    .out(cond93_out),
    .reset(cond93_reset),
    .write_en(cond93_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire93 (
    .in(cond_wire93_in),
    .out(cond_wire93_out)
);
std_reg # (
    .WIDTH(1)
) cond94 (
    .clk(cond94_clk),
    .done(cond94_done),
    .in(cond94_in),
    .out(cond94_out),
    .reset(cond94_reset),
    .write_en(cond94_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire94 (
    .in(cond_wire94_in),
    .out(cond_wire94_out)
);
std_reg # (
    .WIDTH(1)
) cond95 (
    .clk(cond95_clk),
    .done(cond95_done),
    .in(cond95_in),
    .out(cond95_out),
    .reset(cond95_reset),
    .write_en(cond95_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire95 (
    .in(cond_wire95_in),
    .out(cond_wire95_out)
);
std_reg # (
    .WIDTH(1)
) cond96 (
    .clk(cond96_clk),
    .done(cond96_done),
    .in(cond96_in),
    .out(cond96_out),
    .reset(cond96_reset),
    .write_en(cond96_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire96 (
    .in(cond_wire96_in),
    .out(cond_wire96_out)
);
std_reg # (
    .WIDTH(1)
) cond97 (
    .clk(cond97_clk),
    .done(cond97_done),
    .in(cond97_in),
    .out(cond97_out),
    .reset(cond97_reset),
    .write_en(cond97_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire97 (
    .in(cond_wire97_in),
    .out(cond_wire97_out)
);
std_reg # (
    .WIDTH(1)
) cond98 (
    .clk(cond98_clk),
    .done(cond98_done),
    .in(cond98_in),
    .out(cond98_out),
    .reset(cond98_reset),
    .write_en(cond98_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire98 (
    .in(cond_wire98_in),
    .out(cond_wire98_out)
);
std_reg # (
    .WIDTH(1)
) cond99 (
    .clk(cond99_clk),
    .done(cond99_done),
    .in(cond99_in),
    .out(cond99_out),
    .reset(cond99_reset),
    .write_en(cond99_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire99 (
    .in(cond_wire99_in),
    .out(cond_wire99_out)
);
std_reg # (
    .WIDTH(1)
) cond100 (
    .clk(cond100_clk),
    .done(cond100_done),
    .in(cond100_in),
    .out(cond100_out),
    .reset(cond100_reset),
    .write_en(cond100_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire100 (
    .in(cond_wire100_in),
    .out(cond_wire100_out)
);
std_reg # (
    .WIDTH(1)
) cond101 (
    .clk(cond101_clk),
    .done(cond101_done),
    .in(cond101_in),
    .out(cond101_out),
    .reset(cond101_reset),
    .write_en(cond101_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire101 (
    .in(cond_wire101_in),
    .out(cond_wire101_out)
);
std_reg # (
    .WIDTH(1)
) cond102 (
    .clk(cond102_clk),
    .done(cond102_done),
    .in(cond102_in),
    .out(cond102_out),
    .reset(cond102_reset),
    .write_en(cond102_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire102 (
    .in(cond_wire102_in),
    .out(cond_wire102_out)
);
std_reg # (
    .WIDTH(1)
) cond103 (
    .clk(cond103_clk),
    .done(cond103_done),
    .in(cond103_in),
    .out(cond103_out),
    .reset(cond103_reset),
    .write_en(cond103_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire103 (
    .in(cond_wire103_in),
    .out(cond_wire103_out)
);
std_reg # (
    .WIDTH(1)
) cond104 (
    .clk(cond104_clk),
    .done(cond104_done),
    .in(cond104_in),
    .out(cond104_out),
    .reset(cond104_reset),
    .write_en(cond104_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire104 (
    .in(cond_wire104_in),
    .out(cond_wire104_out)
);
std_reg # (
    .WIDTH(1)
) cond105 (
    .clk(cond105_clk),
    .done(cond105_done),
    .in(cond105_in),
    .out(cond105_out),
    .reset(cond105_reset),
    .write_en(cond105_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire105 (
    .in(cond_wire105_in),
    .out(cond_wire105_out)
);
std_reg # (
    .WIDTH(1)
) cond106 (
    .clk(cond106_clk),
    .done(cond106_done),
    .in(cond106_in),
    .out(cond106_out),
    .reset(cond106_reset),
    .write_en(cond106_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire106 (
    .in(cond_wire106_in),
    .out(cond_wire106_out)
);
std_reg # (
    .WIDTH(1)
) cond107 (
    .clk(cond107_clk),
    .done(cond107_done),
    .in(cond107_in),
    .out(cond107_out),
    .reset(cond107_reset),
    .write_en(cond107_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire107 (
    .in(cond_wire107_in),
    .out(cond_wire107_out)
);
std_reg # (
    .WIDTH(1)
) cond108 (
    .clk(cond108_clk),
    .done(cond108_done),
    .in(cond108_in),
    .out(cond108_out),
    .reset(cond108_reset),
    .write_en(cond108_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire108 (
    .in(cond_wire108_in),
    .out(cond_wire108_out)
);
std_reg # (
    .WIDTH(1)
) cond109 (
    .clk(cond109_clk),
    .done(cond109_done),
    .in(cond109_in),
    .out(cond109_out),
    .reset(cond109_reset),
    .write_en(cond109_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire109 (
    .in(cond_wire109_in),
    .out(cond_wire109_out)
);
std_reg # (
    .WIDTH(1)
) cond110 (
    .clk(cond110_clk),
    .done(cond110_done),
    .in(cond110_in),
    .out(cond110_out),
    .reset(cond110_reset),
    .write_en(cond110_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire110 (
    .in(cond_wire110_in),
    .out(cond_wire110_out)
);
std_reg # (
    .WIDTH(1)
) cond111 (
    .clk(cond111_clk),
    .done(cond111_done),
    .in(cond111_in),
    .out(cond111_out),
    .reset(cond111_reset),
    .write_en(cond111_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire111 (
    .in(cond_wire111_in),
    .out(cond_wire111_out)
);
std_reg # (
    .WIDTH(1)
) cond112 (
    .clk(cond112_clk),
    .done(cond112_done),
    .in(cond112_in),
    .out(cond112_out),
    .reset(cond112_reset),
    .write_en(cond112_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire112 (
    .in(cond_wire112_in),
    .out(cond_wire112_out)
);
std_reg # (
    .WIDTH(1)
) cond113 (
    .clk(cond113_clk),
    .done(cond113_done),
    .in(cond113_in),
    .out(cond113_out),
    .reset(cond113_reset),
    .write_en(cond113_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire113 (
    .in(cond_wire113_in),
    .out(cond_wire113_out)
);
std_reg # (
    .WIDTH(1)
) cond114 (
    .clk(cond114_clk),
    .done(cond114_done),
    .in(cond114_in),
    .out(cond114_out),
    .reset(cond114_reset),
    .write_en(cond114_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire114 (
    .in(cond_wire114_in),
    .out(cond_wire114_out)
);
std_reg # (
    .WIDTH(1)
) cond115 (
    .clk(cond115_clk),
    .done(cond115_done),
    .in(cond115_in),
    .out(cond115_out),
    .reset(cond115_reset),
    .write_en(cond115_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire115 (
    .in(cond_wire115_in),
    .out(cond_wire115_out)
);
std_reg # (
    .WIDTH(1)
) cond116 (
    .clk(cond116_clk),
    .done(cond116_done),
    .in(cond116_in),
    .out(cond116_out),
    .reset(cond116_reset),
    .write_en(cond116_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire116 (
    .in(cond_wire116_in),
    .out(cond_wire116_out)
);
std_reg # (
    .WIDTH(1)
) cond117 (
    .clk(cond117_clk),
    .done(cond117_done),
    .in(cond117_in),
    .out(cond117_out),
    .reset(cond117_reset),
    .write_en(cond117_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire117 (
    .in(cond_wire117_in),
    .out(cond_wire117_out)
);
std_reg # (
    .WIDTH(1)
) cond118 (
    .clk(cond118_clk),
    .done(cond118_done),
    .in(cond118_in),
    .out(cond118_out),
    .reset(cond118_reset),
    .write_en(cond118_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire118 (
    .in(cond_wire118_in),
    .out(cond_wire118_out)
);
std_reg # (
    .WIDTH(1)
) cond119 (
    .clk(cond119_clk),
    .done(cond119_done),
    .in(cond119_in),
    .out(cond119_out),
    .reset(cond119_reset),
    .write_en(cond119_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire119 (
    .in(cond_wire119_in),
    .out(cond_wire119_out)
);
std_reg # (
    .WIDTH(1)
) cond120 (
    .clk(cond120_clk),
    .done(cond120_done),
    .in(cond120_in),
    .out(cond120_out),
    .reset(cond120_reset),
    .write_en(cond120_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire120 (
    .in(cond_wire120_in),
    .out(cond_wire120_out)
);
std_reg # (
    .WIDTH(1)
) cond121 (
    .clk(cond121_clk),
    .done(cond121_done),
    .in(cond121_in),
    .out(cond121_out),
    .reset(cond121_reset),
    .write_en(cond121_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire121 (
    .in(cond_wire121_in),
    .out(cond_wire121_out)
);
std_reg # (
    .WIDTH(1)
) cond122 (
    .clk(cond122_clk),
    .done(cond122_done),
    .in(cond122_in),
    .out(cond122_out),
    .reset(cond122_reset),
    .write_en(cond122_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire122 (
    .in(cond_wire122_in),
    .out(cond_wire122_out)
);
std_reg # (
    .WIDTH(1)
) cond123 (
    .clk(cond123_clk),
    .done(cond123_done),
    .in(cond123_in),
    .out(cond123_out),
    .reset(cond123_reset),
    .write_en(cond123_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire123 (
    .in(cond_wire123_in),
    .out(cond_wire123_out)
);
std_reg # (
    .WIDTH(1)
) cond124 (
    .clk(cond124_clk),
    .done(cond124_done),
    .in(cond124_in),
    .out(cond124_out),
    .reset(cond124_reset),
    .write_en(cond124_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire124 (
    .in(cond_wire124_in),
    .out(cond_wire124_out)
);
std_reg # (
    .WIDTH(1)
) cond125 (
    .clk(cond125_clk),
    .done(cond125_done),
    .in(cond125_in),
    .out(cond125_out),
    .reset(cond125_reset),
    .write_en(cond125_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire125 (
    .in(cond_wire125_in),
    .out(cond_wire125_out)
);
std_reg # (
    .WIDTH(1)
) cond126 (
    .clk(cond126_clk),
    .done(cond126_done),
    .in(cond126_in),
    .out(cond126_out),
    .reset(cond126_reset),
    .write_en(cond126_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire126 (
    .in(cond_wire126_in),
    .out(cond_wire126_out)
);
std_reg # (
    .WIDTH(1)
) cond127 (
    .clk(cond127_clk),
    .done(cond127_done),
    .in(cond127_in),
    .out(cond127_out),
    .reset(cond127_reset),
    .write_en(cond127_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire127 (
    .in(cond_wire127_in),
    .out(cond_wire127_out)
);
std_reg # (
    .WIDTH(1)
) cond128 (
    .clk(cond128_clk),
    .done(cond128_done),
    .in(cond128_in),
    .out(cond128_out),
    .reset(cond128_reset),
    .write_en(cond128_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire128 (
    .in(cond_wire128_in),
    .out(cond_wire128_out)
);
std_reg # (
    .WIDTH(1)
) cond129 (
    .clk(cond129_clk),
    .done(cond129_done),
    .in(cond129_in),
    .out(cond129_out),
    .reset(cond129_reset),
    .write_en(cond129_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire129 (
    .in(cond_wire129_in),
    .out(cond_wire129_out)
);
std_reg # (
    .WIDTH(1)
) cond130 (
    .clk(cond130_clk),
    .done(cond130_done),
    .in(cond130_in),
    .out(cond130_out),
    .reset(cond130_reset),
    .write_en(cond130_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire130 (
    .in(cond_wire130_in),
    .out(cond_wire130_out)
);
std_reg # (
    .WIDTH(1)
) cond131 (
    .clk(cond131_clk),
    .done(cond131_done),
    .in(cond131_in),
    .out(cond131_out),
    .reset(cond131_reset),
    .write_en(cond131_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire131 (
    .in(cond_wire131_in),
    .out(cond_wire131_out)
);
std_reg # (
    .WIDTH(1)
) cond132 (
    .clk(cond132_clk),
    .done(cond132_done),
    .in(cond132_in),
    .out(cond132_out),
    .reset(cond132_reset),
    .write_en(cond132_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire132 (
    .in(cond_wire132_in),
    .out(cond_wire132_out)
);
std_reg # (
    .WIDTH(1)
) cond133 (
    .clk(cond133_clk),
    .done(cond133_done),
    .in(cond133_in),
    .out(cond133_out),
    .reset(cond133_reset),
    .write_en(cond133_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire133 (
    .in(cond_wire133_in),
    .out(cond_wire133_out)
);
std_reg # (
    .WIDTH(1)
) cond134 (
    .clk(cond134_clk),
    .done(cond134_done),
    .in(cond134_in),
    .out(cond134_out),
    .reset(cond134_reset),
    .write_en(cond134_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire134 (
    .in(cond_wire134_in),
    .out(cond_wire134_out)
);
std_reg # (
    .WIDTH(1)
) cond135 (
    .clk(cond135_clk),
    .done(cond135_done),
    .in(cond135_in),
    .out(cond135_out),
    .reset(cond135_reset),
    .write_en(cond135_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire135 (
    .in(cond_wire135_in),
    .out(cond_wire135_out)
);
std_reg # (
    .WIDTH(1)
) cond136 (
    .clk(cond136_clk),
    .done(cond136_done),
    .in(cond136_in),
    .out(cond136_out),
    .reset(cond136_reset),
    .write_en(cond136_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire136 (
    .in(cond_wire136_in),
    .out(cond_wire136_out)
);
std_reg # (
    .WIDTH(1)
) cond137 (
    .clk(cond137_clk),
    .done(cond137_done),
    .in(cond137_in),
    .out(cond137_out),
    .reset(cond137_reset),
    .write_en(cond137_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire137 (
    .in(cond_wire137_in),
    .out(cond_wire137_out)
);
std_reg # (
    .WIDTH(1)
) cond138 (
    .clk(cond138_clk),
    .done(cond138_done),
    .in(cond138_in),
    .out(cond138_out),
    .reset(cond138_reset),
    .write_en(cond138_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire138 (
    .in(cond_wire138_in),
    .out(cond_wire138_out)
);
std_reg # (
    .WIDTH(1)
) cond139 (
    .clk(cond139_clk),
    .done(cond139_done),
    .in(cond139_in),
    .out(cond139_out),
    .reset(cond139_reset),
    .write_en(cond139_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire139 (
    .in(cond_wire139_in),
    .out(cond_wire139_out)
);
std_reg # (
    .WIDTH(1)
) cond140 (
    .clk(cond140_clk),
    .done(cond140_done),
    .in(cond140_in),
    .out(cond140_out),
    .reset(cond140_reset),
    .write_en(cond140_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire140 (
    .in(cond_wire140_in),
    .out(cond_wire140_out)
);
std_reg # (
    .WIDTH(1)
) cond141 (
    .clk(cond141_clk),
    .done(cond141_done),
    .in(cond141_in),
    .out(cond141_out),
    .reset(cond141_reset),
    .write_en(cond141_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire141 (
    .in(cond_wire141_in),
    .out(cond_wire141_out)
);
std_reg # (
    .WIDTH(1)
) cond142 (
    .clk(cond142_clk),
    .done(cond142_done),
    .in(cond142_in),
    .out(cond142_out),
    .reset(cond142_reset),
    .write_en(cond142_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire142 (
    .in(cond_wire142_in),
    .out(cond_wire142_out)
);
std_reg # (
    .WIDTH(1)
) cond143 (
    .clk(cond143_clk),
    .done(cond143_done),
    .in(cond143_in),
    .out(cond143_out),
    .reset(cond143_reset),
    .write_en(cond143_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire143 (
    .in(cond_wire143_in),
    .out(cond_wire143_out)
);
std_reg # (
    .WIDTH(1)
) cond144 (
    .clk(cond144_clk),
    .done(cond144_done),
    .in(cond144_in),
    .out(cond144_out),
    .reset(cond144_reset),
    .write_en(cond144_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire144 (
    .in(cond_wire144_in),
    .out(cond_wire144_out)
);
std_reg # (
    .WIDTH(1)
) cond145 (
    .clk(cond145_clk),
    .done(cond145_done),
    .in(cond145_in),
    .out(cond145_out),
    .reset(cond145_reset),
    .write_en(cond145_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire145 (
    .in(cond_wire145_in),
    .out(cond_wire145_out)
);
std_reg # (
    .WIDTH(1)
) cond146 (
    .clk(cond146_clk),
    .done(cond146_done),
    .in(cond146_in),
    .out(cond146_out),
    .reset(cond146_reset),
    .write_en(cond146_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire146 (
    .in(cond_wire146_in),
    .out(cond_wire146_out)
);
std_reg # (
    .WIDTH(1)
) cond147 (
    .clk(cond147_clk),
    .done(cond147_done),
    .in(cond147_in),
    .out(cond147_out),
    .reset(cond147_reset),
    .write_en(cond147_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire147 (
    .in(cond_wire147_in),
    .out(cond_wire147_out)
);
std_reg # (
    .WIDTH(1)
) cond148 (
    .clk(cond148_clk),
    .done(cond148_done),
    .in(cond148_in),
    .out(cond148_out),
    .reset(cond148_reset),
    .write_en(cond148_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire148 (
    .in(cond_wire148_in),
    .out(cond_wire148_out)
);
std_reg # (
    .WIDTH(1)
) cond149 (
    .clk(cond149_clk),
    .done(cond149_done),
    .in(cond149_in),
    .out(cond149_out),
    .reset(cond149_reset),
    .write_en(cond149_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire149 (
    .in(cond_wire149_in),
    .out(cond_wire149_out)
);
std_reg # (
    .WIDTH(1)
) cond150 (
    .clk(cond150_clk),
    .done(cond150_done),
    .in(cond150_in),
    .out(cond150_out),
    .reset(cond150_reset),
    .write_en(cond150_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire150 (
    .in(cond_wire150_in),
    .out(cond_wire150_out)
);
std_reg # (
    .WIDTH(1)
) cond151 (
    .clk(cond151_clk),
    .done(cond151_done),
    .in(cond151_in),
    .out(cond151_out),
    .reset(cond151_reset),
    .write_en(cond151_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire151 (
    .in(cond_wire151_in),
    .out(cond_wire151_out)
);
std_reg # (
    .WIDTH(1)
) cond152 (
    .clk(cond152_clk),
    .done(cond152_done),
    .in(cond152_in),
    .out(cond152_out),
    .reset(cond152_reset),
    .write_en(cond152_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire152 (
    .in(cond_wire152_in),
    .out(cond_wire152_out)
);
std_reg # (
    .WIDTH(1)
) cond153 (
    .clk(cond153_clk),
    .done(cond153_done),
    .in(cond153_in),
    .out(cond153_out),
    .reset(cond153_reset),
    .write_en(cond153_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire153 (
    .in(cond_wire153_in),
    .out(cond_wire153_out)
);
std_reg # (
    .WIDTH(1)
) cond154 (
    .clk(cond154_clk),
    .done(cond154_done),
    .in(cond154_in),
    .out(cond154_out),
    .reset(cond154_reset),
    .write_en(cond154_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire154 (
    .in(cond_wire154_in),
    .out(cond_wire154_out)
);
std_reg # (
    .WIDTH(1)
) cond155 (
    .clk(cond155_clk),
    .done(cond155_done),
    .in(cond155_in),
    .out(cond155_out),
    .reset(cond155_reset),
    .write_en(cond155_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire155 (
    .in(cond_wire155_in),
    .out(cond_wire155_out)
);
std_reg # (
    .WIDTH(1)
) cond156 (
    .clk(cond156_clk),
    .done(cond156_done),
    .in(cond156_in),
    .out(cond156_out),
    .reset(cond156_reset),
    .write_en(cond156_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire156 (
    .in(cond_wire156_in),
    .out(cond_wire156_out)
);
std_reg # (
    .WIDTH(1)
) cond157 (
    .clk(cond157_clk),
    .done(cond157_done),
    .in(cond157_in),
    .out(cond157_out),
    .reset(cond157_reset),
    .write_en(cond157_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire157 (
    .in(cond_wire157_in),
    .out(cond_wire157_out)
);
std_reg # (
    .WIDTH(1)
) cond158 (
    .clk(cond158_clk),
    .done(cond158_done),
    .in(cond158_in),
    .out(cond158_out),
    .reset(cond158_reset),
    .write_en(cond158_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire158 (
    .in(cond_wire158_in),
    .out(cond_wire158_out)
);
std_reg # (
    .WIDTH(1)
) cond159 (
    .clk(cond159_clk),
    .done(cond159_done),
    .in(cond159_in),
    .out(cond159_out),
    .reset(cond159_reset),
    .write_en(cond159_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire159 (
    .in(cond_wire159_in),
    .out(cond_wire159_out)
);
std_reg # (
    .WIDTH(1)
) cond160 (
    .clk(cond160_clk),
    .done(cond160_done),
    .in(cond160_in),
    .out(cond160_out),
    .reset(cond160_reset),
    .write_en(cond160_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire160 (
    .in(cond_wire160_in),
    .out(cond_wire160_out)
);
std_reg # (
    .WIDTH(1)
) cond161 (
    .clk(cond161_clk),
    .done(cond161_done),
    .in(cond161_in),
    .out(cond161_out),
    .reset(cond161_reset),
    .write_en(cond161_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire161 (
    .in(cond_wire161_in),
    .out(cond_wire161_out)
);
std_reg # (
    .WIDTH(1)
) cond162 (
    .clk(cond162_clk),
    .done(cond162_done),
    .in(cond162_in),
    .out(cond162_out),
    .reset(cond162_reset),
    .write_en(cond162_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire162 (
    .in(cond_wire162_in),
    .out(cond_wire162_out)
);
std_reg # (
    .WIDTH(1)
) cond163 (
    .clk(cond163_clk),
    .done(cond163_done),
    .in(cond163_in),
    .out(cond163_out),
    .reset(cond163_reset),
    .write_en(cond163_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire163 (
    .in(cond_wire163_in),
    .out(cond_wire163_out)
);
std_reg # (
    .WIDTH(1)
) cond164 (
    .clk(cond164_clk),
    .done(cond164_done),
    .in(cond164_in),
    .out(cond164_out),
    .reset(cond164_reset),
    .write_en(cond164_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire164 (
    .in(cond_wire164_in),
    .out(cond_wire164_out)
);
std_reg # (
    .WIDTH(1)
) cond165 (
    .clk(cond165_clk),
    .done(cond165_done),
    .in(cond165_in),
    .out(cond165_out),
    .reset(cond165_reset),
    .write_en(cond165_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire165 (
    .in(cond_wire165_in),
    .out(cond_wire165_out)
);
std_reg # (
    .WIDTH(1)
) cond166 (
    .clk(cond166_clk),
    .done(cond166_done),
    .in(cond166_in),
    .out(cond166_out),
    .reset(cond166_reset),
    .write_en(cond166_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire166 (
    .in(cond_wire166_in),
    .out(cond_wire166_out)
);
std_reg # (
    .WIDTH(1)
) cond167 (
    .clk(cond167_clk),
    .done(cond167_done),
    .in(cond167_in),
    .out(cond167_out),
    .reset(cond167_reset),
    .write_en(cond167_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire167 (
    .in(cond_wire167_in),
    .out(cond_wire167_out)
);
std_reg # (
    .WIDTH(1)
) cond168 (
    .clk(cond168_clk),
    .done(cond168_done),
    .in(cond168_in),
    .out(cond168_out),
    .reset(cond168_reset),
    .write_en(cond168_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire168 (
    .in(cond_wire168_in),
    .out(cond_wire168_out)
);
std_reg # (
    .WIDTH(1)
) cond169 (
    .clk(cond169_clk),
    .done(cond169_done),
    .in(cond169_in),
    .out(cond169_out),
    .reset(cond169_reset),
    .write_en(cond169_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire169 (
    .in(cond_wire169_in),
    .out(cond_wire169_out)
);
std_reg # (
    .WIDTH(1)
) cond170 (
    .clk(cond170_clk),
    .done(cond170_done),
    .in(cond170_in),
    .out(cond170_out),
    .reset(cond170_reset),
    .write_en(cond170_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire170 (
    .in(cond_wire170_in),
    .out(cond_wire170_out)
);
std_reg # (
    .WIDTH(1)
) cond171 (
    .clk(cond171_clk),
    .done(cond171_done),
    .in(cond171_in),
    .out(cond171_out),
    .reset(cond171_reset),
    .write_en(cond171_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire171 (
    .in(cond_wire171_in),
    .out(cond_wire171_out)
);
std_reg # (
    .WIDTH(1)
) cond172 (
    .clk(cond172_clk),
    .done(cond172_done),
    .in(cond172_in),
    .out(cond172_out),
    .reset(cond172_reset),
    .write_en(cond172_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire172 (
    .in(cond_wire172_in),
    .out(cond_wire172_out)
);
std_reg # (
    .WIDTH(1)
) cond173 (
    .clk(cond173_clk),
    .done(cond173_done),
    .in(cond173_in),
    .out(cond173_out),
    .reset(cond173_reset),
    .write_en(cond173_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire173 (
    .in(cond_wire173_in),
    .out(cond_wire173_out)
);
std_reg # (
    .WIDTH(1)
) cond174 (
    .clk(cond174_clk),
    .done(cond174_done),
    .in(cond174_in),
    .out(cond174_out),
    .reset(cond174_reset),
    .write_en(cond174_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire174 (
    .in(cond_wire174_in),
    .out(cond_wire174_out)
);
std_reg # (
    .WIDTH(1)
) cond175 (
    .clk(cond175_clk),
    .done(cond175_done),
    .in(cond175_in),
    .out(cond175_out),
    .reset(cond175_reset),
    .write_en(cond175_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire175 (
    .in(cond_wire175_in),
    .out(cond_wire175_out)
);
std_reg # (
    .WIDTH(1)
) cond176 (
    .clk(cond176_clk),
    .done(cond176_done),
    .in(cond176_in),
    .out(cond176_out),
    .reset(cond176_reset),
    .write_en(cond176_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire176 (
    .in(cond_wire176_in),
    .out(cond_wire176_out)
);
std_reg # (
    .WIDTH(1)
) cond177 (
    .clk(cond177_clk),
    .done(cond177_done),
    .in(cond177_in),
    .out(cond177_out),
    .reset(cond177_reset),
    .write_en(cond177_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire177 (
    .in(cond_wire177_in),
    .out(cond_wire177_out)
);
std_reg # (
    .WIDTH(1)
) cond178 (
    .clk(cond178_clk),
    .done(cond178_done),
    .in(cond178_in),
    .out(cond178_out),
    .reset(cond178_reset),
    .write_en(cond178_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire178 (
    .in(cond_wire178_in),
    .out(cond_wire178_out)
);
std_reg # (
    .WIDTH(1)
) cond179 (
    .clk(cond179_clk),
    .done(cond179_done),
    .in(cond179_in),
    .out(cond179_out),
    .reset(cond179_reset),
    .write_en(cond179_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire179 (
    .in(cond_wire179_in),
    .out(cond_wire179_out)
);
std_reg # (
    .WIDTH(1)
) cond180 (
    .clk(cond180_clk),
    .done(cond180_done),
    .in(cond180_in),
    .out(cond180_out),
    .reset(cond180_reset),
    .write_en(cond180_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire180 (
    .in(cond_wire180_in),
    .out(cond_wire180_out)
);
std_reg # (
    .WIDTH(1)
) cond181 (
    .clk(cond181_clk),
    .done(cond181_done),
    .in(cond181_in),
    .out(cond181_out),
    .reset(cond181_reset),
    .write_en(cond181_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire181 (
    .in(cond_wire181_in),
    .out(cond_wire181_out)
);
std_reg # (
    .WIDTH(1)
) cond182 (
    .clk(cond182_clk),
    .done(cond182_done),
    .in(cond182_in),
    .out(cond182_out),
    .reset(cond182_reset),
    .write_en(cond182_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire182 (
    .in(cond_wire182_in),
    .out(cond_wire182_out)
);
std_reg # (
    .WIDTH(1)
) cond183 (
    .clk(cond183_clk),
    .done(cond183_done),
    .in(cond183_in),
    .out(cond183_out),
    .reset(cond183_reset),
    .write_en(cond183_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire183 (
    .in(cond_wire183_in),
    .out(cond_wire183_out)
);
std_reg # (
    .WIDTH(1)
) cond184 (
    .clk(cond184_clk),
    .done(cond184_done),
    .in(cond184_in),
    .out(cond184_out),
    .reset(cond184_reset),
    .write_en(cond184_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire184 (
    .in(cond_wire184_in),
    .out(cond_wire184_out)
);
std_reg # (
    .WIDTH(1)
) cond185 (
    .clk(cond185_clk),
    .done(cond185_done),
    .in(cond185_in),
    .out(cond185_out),
    .reset(cond185_reset),
    .write_en(cond185_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire185 (
    .in(cond_wire185_in),
    .out(cond_wire185_out)
);
std_reg # (
    .WIDTH(1)
) cond186 (
    .clk(cond186_clk),
    .done(cond186_done),
    .in(cond186_in),
    .out(cond186_out),
    .reset(cond186_reset),
    .write_en(cond186_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire186 (
    .in(cond_wire186_in),
    .out(cond_wire186_out)
);
std_reg # (
    .WIDTH(1)
) cond187 (
    .clk(cond187_clk),
    .done(cond187_done),
    .in(cond187_in),
    .out(cond187_out),
    .reset(cond187_reset),
    .write_en(cond187_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire187 (
    .in(cond_wire187_in),
    .out(cond_wire187_out)
);
std_reg # (
    .WIDTH(1)
) cond188 (
    .clk(cond188_clk),
    .done(cond188_done),
    .in(cond188_in),
    .out(cond188_out),
    .reset(cond188_reset),
    .write_en(cond188_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire188 (
    .in(cond_wire188_in),
    .out(cond_wire188_out)
);
std_reg # (
    .WIDTH(1)
) cond189 (
    .clk(cond189_clk),
    .done(cond189_done),
    .in(cond189_in),
    .out(cond189_out),
    .reset(cond189_reset),
    .write_en(cond189_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire189 (
    .in(cond_wire189_in),
    .out(cond_wire189_out)
);
std_reg # (
    .WIDTH(1)
) cond190 (
    .clk(cond190_clk),
    .done(cond190_done),
    .in(cond190_in),
    .out(cond190_out),
    .reset(cond190_reset),
    .write_en(cond190_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire190 (
    .in(cond_wire190_in),
    .out(cond_wire190_out)
);
std_reg # (
    .WIDTH(1)
) cond191 (
    .clk(cond191_clk),
    .done(cond191_done),
    .in(cond191_in),
    .out(cond191_out),
    .reset(cond191_reset),
    .write_en(cond191_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire191 (
    .in(cond_wire191_in),
    .out(cond_wire191_out)
);
std_reg # (
    .WIDTH(1)
) cond192 (
    .clk(cond192_clk),
    .done(cond192_done),
    .in(cond192_in),
    .out(cond192_out),
    .reset(cond192_reset),
    .write_en(cond192_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire192 (
    .in(cond_wire192_in),
    .out(cond_wire192_out)
);
std_reg # (
    .WIDTH(1)
) cond193 (
    .clk(cond193_clk),
    .done(cond193_done),
    .in(cond193_in),
    .out(cond193_out),
    .reset(cond193_reset),
    .write_en(cond193_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire193 (
    .in(cond_wire193_in),
    .out(cond_wire193_out)
);
std_reg # (
    .WIDTH(1)
) cond194 (
    .clk(cond194_clk),
    .done(cond194_done),
    .in(cond194_in),
    .out(cond194_out),
    .reset(cond194_reset),
    .write_en(cond194_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire194 (
    .in(cond_wire194_in),
    .out(cond_wire194_out)
);
std_reg # (
    .WIDTH(1)
) cond195 (
    .clk(cond195_clk),
    .done(cond195_done),
    .in(cond195_in),
    .out(cond195_out),
    .reset(cond195_reset),
    .write_en(cond195_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire195 (
    .in(cond_wire195_in),
    .out(cond_wire195_out)
);
std_reg # (
    .WIDTH(1)
) cond196 (
    .clk(cond196_clk),
    .done(cond196_done),
    .in(cond196_in),
    .out(cond196_out),
    .reset(cond196_reset),
    .write_en(cond196_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire196 (
    .in(cond_wire196_in),
    .out(cond_wire196_out)
);
std_reg # (
    .WIDTH(1)
) cond197 (
    .clk(cond197_clk),
    .done(cond197_done),
    .in(cond197_in),
    .out(cond197_out),
    .reset(cond197_reset),
    .write_en(cond197_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire197 (
    .in(cond_wire197_in),
    .out(cond_wire197_out)
);
std_reg # (
    .WIDTH(1)
) cond198 (
    .clk(cond198_clk),
    .done(cond198_done),
    .in(cond198_in),
    .out(cond198_out),
    .reset(cond198_reset),
    .write_en(cond198_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire198 (
    .in(cond_wire198_in),
    .out(cond_wire198_out)
);
std_reg # (
    .WIDTH(1)
) cond199 (
    .clk(cond199_clk),
    .done(cond199_done),
    .in(cond199_in),
    .out(cond199_out),
    .reset(cond199_reset),
    .write_en(cond199_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire199 (
    .in(cond_wire199_in),
    .out(cond_wire199_out)
);
std_reg # (
    .WIDTH(1)
) cond200 (
    .clk(cond200_clk),
    .done(cond200_done),
    .in(cond200_in),
    .out(cond200_out),
    .reset(cond200_reset),
    .write_en(cond200_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire200 (
    .in(cond_wire200_in),
    .out(cond_wire200_out)
);
std_reg # (
    .WIDTH(1)
) cond201 (
    .clk(cond201_clk),
    .done(cond201_done),
    .in(cond201_in),
    .out(cond201_out),
    .reset(cond201_reset),
    .write_en(cond201_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire201 (
    .in(cond_wire201_in),
    .out(cond_wire201_out)
);
std_reg # (
    .WIDTH(1)
) cond202 (
    .clk(cond202_clk),
    .done(cond202_done),
    .in(cond202_in),
    .out(cond202_out),
    .reset(cond202_reset),
    .write_en(cond202_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire202 (
    .in(cond_wire202_in),
    .out(cond_wire202_out)
);
std_reg # (
    .WIDTH(1)
) cond203 (
    .clk(cond203_clk),
    .done(cond203_done),
    .in(cond203_in),
    .out(cond203_out),
    .reset(cond203_reset),
    .write_en(cond203_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire203 (
    .in(cond_wire203_in),
    .out(cond_wire203_out)
);
std_reg # (
    .WIDTH(1)
) cond204 (
    .clk(cond204_clk),
    .done(cond204_done),
    .in(cond204_in),
    .out(cond204_out),
    .reset(cond204_reset),
    .write_en(cond204_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire204 (
    .in(cond_wire204_in),
    .out(cond_wire204_out)
);
std_reg # (
    .WIDTH(1)
) cond205 (
    .clk(cond205_clk),
    .done(cond205_done),
    .in(cond205_in),
    .out(cond205_out),
    .reset(cond205_reset),
    .write_en(cond205_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire205 (
    .in(cond_wire205_in),
    .out(cond_wire205_out)
);
std_reg # (
    .WIDTH(1)
) cond206 (
    .clk(cond206_clk),
    .done(cond206_done),
    .in(cond206_in),
    .out(cond206_out),
    .reset(cond206_reset),
    .write_en(cond206_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire206 (
    .in(cond_wire206_in),
    .out(cond_wire206_out)
);
std_reg # (
    .WIDTH(1)
) cond207 (
    .clk(cond207_clk),
    .done(cond207_done),
    .in(cond207_in),
    .out(cond207_out),
    .reset(cond207_reset),
    .write_en(cond207_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire207 (
    .in(cond_wire207_in),
    .out(cond_wire207_out)
);
std_reg # (
    .WIDTH(1)
) cond208 (
    .clk(cond208_clk),
    .done(cond208_done),
    .in(cond208_in),
    .out(cond208_out),
    .reset(cond208_reset),
    .write_en(cond208_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire208 (
    .in(cond_wire208_in),
    .out(cond_wire208_out)
);
std_reg # (
    .WIDTH(1)
) cond209 (
    .clk(cond209_clk),
    .done(cond209_done),
    .in(cond209_in),
    .out(cond209_out),
    .reset(cond209_reset),
    .write_en(cond209_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire209 (
    .in(cond_wire209_in),
    .out(cond_wire209_out)
);
std_reg # (
    .WIDTH(1)
) cond210 (
    .clk(cond210_clk),
    .done(cond210_done),
    .in(cond210_in),
    .out(cond210_out),
    .reset(cond210_reset),
    .write_en(cond210_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire210 (
    .in(cond_wire210_in),
    .out(cond_wire210_out)
);
std_reg # (
    .WIDTH(1)
) cond211 (
    .clk(cond211_clk),
    .done(cond211_done),
    .in(cond211_in),
    .out(cond211_out),
    .reset(cond211_reset),
    .write_en(cond211_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire211 (
    .in(cond_wire211_in),
    .out(cond_wire211_out)
);
std_reg # (
    .WIDTH(1)
) cond212 (
    .clk(cond212_clk),
    .done(cond212_done),
    .in(cond212_in),
    .out(cond212_out),
    .reset(cond212_reset),
    .write_en(cond212_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire212 (
    .in(cond_wire212_in),
    .out(cond_wire212_out)
);
std_reg # (
    .WIDTH(1)
) cond213 (
    .clk(cond213_clk),
    .done(cond213_done),
    .in(cond213_in),
    .out(cond213_out),
    .reset(cond213_reset),
    .write_en(cond213_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire213 (
    .in(cond_wire213_in),
    .out(cond_wire213_out)
);
std_reg # (
    .WIDTH(1)
) cond214 (
    .clk(cond214_clk),
    .done(cond214_done),
    .in(cond214_in),
    .out(cond214_out),
    .reset(cond214_reset),
    .write_en(cond214_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire214 (
    .in(cond_wire214_in),
    .out(cond_wire214_out)
);
std_reg # (
    .WIDTH(1)
) cond215 (
    .clk(cond215_clk),
    .done(cond215_done),
    .in(cond215_in),
    .out(cond215_out),
    .reset(cond215_reset),
    .write_en(cond215_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire215 (
    .in(cond_wire215_in),
    .out(cond_wire215_out)
);
std_reg # (
    .WIDTH(1)
) cond216 (
    .clk(cond216_clk),
    .done(cond216_done),
    .in(cond216_in),
    .out(cond216_out),
    .reset(cond216_reset),
    .write_en(cond216_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire216 (
    .in(cond_wire216_in),
    .out(cond_wire216_out)
);
std_reg # (
    .WIDTH(1)
) cond217 (
    .clk(cond217_clk),
    .done(cond217_done),
    .in(cond217_in),
    .out(cond217_out),
    .reset(cond217_reset),
    .write_en(cond217_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire217 (
    .in(cond_wire217_in),
    .out(cond_wire217_out)
);
std_reg # (
    .WIDTH(1)
) cond218 (
    .clk(cond218_clk),
    .done(cond218_done),
    .in(cond218_in),
    .out(cond218_out),
    .reset(cond218_reset),
    .write_en(cond218_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire218 (
    .in(cond_wire218_in),
    .out(cond_wire218_out)
);
std_reg # (
    .WIDTH(1)
) cond219 (
    .clk(cond219_clk),
    .done(cond219_done),
    .in(cond219_in),
    .out(cond219_out),
    .reset(cond219_reset),
    .write_en(cond219_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire219 (
    .in(cond_wire219_in),
    .out(cond_wire219_out)
);
std_reg # (
    .WIDTH(1)
) cond220 (
    .clk(cond220_clk),
    .done(cond220_done),
    .in(cond220_in),
    .out(cond220_out),
    .reset(cond220_reset),
    .write_en(cond220_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire220 (
    .in(cond_wire220_in),
    .out(cond_wire220_out)
);
std_reg # (
    .WIDTH(1)
) cond221 (
    .clk(cond221_clk),
    .done(cond221_done),
    .in(cond221_in),
    .out(cond221_out),
    .reset(cond221_reset),
    .write_en(cond221_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire221 (
    .in(cond_wire221_in),
    .out(cond_wire221_out)
);
std_reg # (
    .WIDTH(1)
) cond222 (
    .clk(cond222_clk),
    .done(cond222_done),
    .in(cond222_in),
    .out(cond222_out),
    .reset(cond222_reset),
    .write_en(cond222_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire222 (
    .in(cond_wire222_in),
    .out(cond_wire222_out)
);
std_reg # (
    .WIDTH(1)
) cond223 (
    .clk(cond223_clk),
    .done(cond223_done),
    .in(cond223_in),
    .out(cond223_out),
    .reset(cond223_reset),
    .write_en(cond223_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire223 (
    .in(cond_wire223_in),
    .out(cond_wire223_out)
);
std_reg # (
    .WIDTH(1)
) cond224 (
    .clk(cond224_clk),
    .done(cond224_done),
    .in(cond224_in),
    .out(cond224_out),
    .reset(cond224_reset),
    .write_en(cond224_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire224 (
    .in(cond_wire224_in),
    .out(cond_wire224_out)
);
std_reg # (
    .WIDTH(1)
) cond225 (
    .clk(cond225_clk),
    .done(cond225_done),
    .in(cond225_in),
    .out(cond225_out),
    .reset(cond225_reset),
    .write_en(cond225_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire225 (
    .in(cond_wire225_in),
    .out(cond_wire225_out)
);
std_reg # (
    .WIDTH(1)
) cond226 (
    .clk(cond226_clk),
    .done(cond226_done),
    .in(cond226_in),
    .out(cond226_out),
    .reset(cond226_reset),
    .write_en(cond226_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire226 (
    .in(cond_wire226_in),
    .out(cond_wire226_out)
);
std_reg # (
    .WIDTH(1)
) cond227 (
    .clk(cond227_clk),
    .done(cond227_done),
    .in(cond227_in),
    .out(cond227_out),
    .reset(cond227_reset),
    .write_en(cond227_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire227 (
    .in(cond_wire227_in),
    .out(cond_wire227_out)
);
std_reg # (
    .WIDTH(1)
) cond228 (
    .clk(cond228_clk),
    .done(cond228_done),
    .in(cond228_in),
    .out(cond228_out),
    .reset(cond228_reset),
    .write_en(cond228_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire228 (
    .in(cond_wire228_in),
    .out(cond_wire228_out)
);
std_reg # (
    .WIDTH(1)
) cond229 (
    .clk(cond229_clk),
    .done(cond229_done),
    .in(cond229_in),
    .out(cond229_out),
    .reset(cond229_reset),
    .write_en(cond229_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire229 (
    .in(cond_wire229_in),
    .out(cond_wire229_out)
);
std_reg # (
    .WIDTH(1)
) cond230 (
    .clk(cond230_clk),
    .done(cond230_done),
    .in(cond230_in),
    .out(cond230_out),
    .reset(cond230_reset),
    .write_en(cond230_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire230 (
    .in(cond_wire230_in),
    .out(cond_wire230_out)
);
std_reg # (
    .WIDTH(1)
) cond231 (
    .clk(cond231_clk),
    .done(cond231_done),
    .in(cond231_in),
    .out(cond231_out),
    .reset(cond231_reset),
    .write_en(cond231_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire231 (
    .in(cond_wire231_in),
    .out(cond_wire231_out)
);
std_reg # (
    .WIDTH(1)
) cond232 (
    .clk(cond232_clk),
    .done(cond232_done),
    .in(cond232_in),
    .out(cond232_out),
    .reset(cond232_reset),
    .write_en(cond232_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire232 (
    .in(cond_wire232_in),
    .out(cond_wire232_out)
);
std_reg # (
    .WIDTH(1)
) cond233 (
    .clk(cond233_clk),
    .done(cond233_done),
    .in(cond233_in),
    .out(cond233_out),
    .reset(cond233_reset),
    .write_en(cond233_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire233 (
    .in(cond_wire233_in),
    .out(cond_wire233_out)
);
std_reg # (
    .WIDTH(1)
) cond234 (
    .clk(cond234_clk),
    .done(cond234_done),
    .in(cond234_in),
    .out(cond234_out),
    .reset(cond234_reset),
    .write_en(cond234_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire234 (
    .in(cond_wire234_in),
    .out(cond_wire234_out)
);
std_reg # (
    .WIDTH(1)
) cond235 (
    .clk(cond235_clk),
    .done(cond235_done),
    .in(cond235_in),
    .out(cond235_out),
    .reset(cond235_reset),
    .write_en(cond235_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire235 (
    .in(cond_wire235_in),
    .out(cond_wire235_out)
);
std_reg # (
    .WIDTH(1)
) cond236 (
    .clk(cond236_clk),
    .done(cond236_done),
    .in(cond236_in),
    .out(cond236_out),
    .reset(cond236_reset),
    .write_en(cond236_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire236 (
    .in(cond_wire236_in),
    .out(cond_wire236_out)
);
std_reg # (
    .WIDTH(1)
) cond237 (
    .clk(cond237_clk),
    .done(cond237_done),
    .in(cond237_in),
    .out(cond237_out),
    .reset(cond237_reset),
    .write_en(cond237_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire237 (
    .in(cond_wire237_in),
    .out(cond_wire237_out)
);
std_reg # (
    .WIDTH(1)
) cond238 (
    .clk(cond238_clk),
    .done(cond238_done),
    .in(cond238_in),
    .out(cond238_out),
    .reset(cond238_reset),
    .write_en(cond238_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire238 (
    .in(cond_wire238_in),
    .out(cond_wire238_out)
);
std_reg # (
    .WIDTH(1)
) cond239 (
    .clk(cond239_clk),
    .done(cond239_done),
    .in(cond239_in),
    .out(cond239_out),
    .reset(cond239_reset),
    .write_en(cond239_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire239 (
    .in(cond_wire239_in),
    .out(cond_wire239_out)
);
std_reg # (
    .WIDTH(1)
) cond240 (
    .clk(cond240_clk),
    .done(cond240_done),
    .in(cond240_in),
    .out(cond240_out),
    .reset(cond240_reset),
    .write_en(cond240_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire240 (
    .in(cond_wire240_in),
    .out(cond_wire240_out)
);
std_reg # (
    .WIDTH(1)
) cond241 (
    .clk(cond241_clk),
    .done(cond241_done),
    .in(cond241_in),
    .out(cond241_out),
    .reset(cond241_reset),
    .write_en(cond241_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire241 (
    .in(cond_wire241_in),
    .out(cond_wire241_out)
);
std_reg # (
    .WIDTH(1)
) cond242 (
    .clk(cond242_clk),
    .done(cond242_done),
    .in(cond242_in),
    .out(cond242_out),
    .reset(cond242_reset),
    .write_en(cond242_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire242 (
    .in(cond_wire242_in),
    .out(cond_wire242_out)
);
std_reg # (
    .WIDTH(1)
) cond243 (
    .clk(cond243_clk),
    .done(cond243_done),
    .in(cond243_in),
    .out(cond243_out),
    .reset(cond243_reset),
    .write_en(cond243_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire243 (
    .in(cond_wire243_in),
    .out(cond_wire243_out)
);
std_reg # (
    .WIDTH(1)
) cond244 (
    .clk(cond244_clk),
    .done(cond244_done),
    .in(cond244_in),
    .out(cond244_out),
    .reset(cond244_reset),
    .write_en(cond244_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire244 (
    .in(cond_wire244_in),
    .out(cond_wire244_out)
);
std_reg # (
    .WIDTH(1)
) cond245 (
    .clk(cond245_clk),
    .done(cond245_done),
    .in(cond245_in),
    .out(cond245_out),
    .reset(cond245_reset),
    .write_en(cond245_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire245 (
    .in(cond_wire245_in),
    .out(cond_wire245_out)
);
std_reg # (
    .WIDTH(1)
) cond246 (
    .clk(cond246_clk),
    .done(cond246_done),
    .in(cond246_in),
    .out(cond246_out),
    .reset(cond246_reset),
    .write_en(cond246_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire246 (
    .in(cond_wire246_in),
    .out(cond_wire246_out)
);
std_reg # (
    .WIDTH(1)
) cond247 (
    .clk(cond247_clk),
    .done(cond247_done),
    .in(cond247_in),
    .out(cond247_out),
    .reset(cond247_reset),
    .write_en(cond247_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire247 (
    .in(cond_wire247_in),
    .out(cond_wire247_out)
);
std_reg # (
    .WIDTH(1)
) cond248 (
    .clk(cond248_clk),
    .done(cond248_done),
    .in(cond248_in),
    .out(cond248_out),
    .reset(cond248_reset),
    .write_en(cond248_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire248 (
    .in(cond_wire248_in),
    .out(cond_wire248_out)
);
std_reg # (
    .WIDTH(1)
) cond249 (
    .clk(cond249_clk),
    .done(cond249_done),
    .in(cond249_in),
    .out(cond249_out),
    .reset(cond249_reset),
    .write_en(cond249_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire249 (
    .in(cond_wire249_in),
    .out(cond_wire249_out)
);
std_reg # (
    .WIDTH(1)
) cond250 (
    .clk(cond250_clk),
    .done(cond250_done),
    .in(cond250_in),
    .out(cond250_out),
    .reset(cond250_reset),
    .write_en(cond250_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire250 (
    .in(cond_wire250_in),
    .out(cond_wire250_out)
);
std_reg # (
    .WIDTH(1)
) cond251 (
    .clk(cond251_clk),
    .done(cond251_done),
    .in(cond251_in),
    .out(cond251_out),
    .reset(cond251_reset),
    .write_en(cond251_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire251 (
    .in(cond_wire251_in),
    .out(cond_wire251_out)
);
std_reg # (
    .WIDTH(1)
) cond252 (
    .clk(cond252_clk),
    .done(cond252_done),
    .in(cond252_in),
    .out(cond252_out),
    .reset(cond252_reset),
    .write_en(cond252_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire252 (
    .in(cond_wire252_in),
    .out(cond_wire252_out)
);
std_reg # (
    .WIDTH(1)
) cond253 (
    .clk(cond253_clk),
    .done(cond253_done),
    .in(cond253_in),
    .out(cond253_out),
    .reset(cond253_reset),
    .write_en(cond253_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire253 (
    .in(cond_wire253_in),
    .out(cond_wire253_out)
);
std_reg # (
    .WIDTH(1)
) cond254 (
    .clk(cond254_clk),
    .done(cond254_done),
    .in(cond254_in),
    .out(cond254_out),
    .reset(cond254_reset),
    .write_en(cond254_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire254 (
    .in(cond_wire254_in),
    .out(cond_wire254_out)
);
std_reg # (
    .WIDTH(1)
) cond255 (
    .clk(cond255_clk),
    .done(cond255_done),
    .in(cond255_in),
    .out(cond255_out),
    .reset(cond255_reset),
    .write_en(cond255_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire255 (
    .in(cond_wire255_in),
    .out(cond_wire255_out)
);
std_reg # (
    .WIDTH(1)
) cond256 (
    .clk(cond256_clk),
    .done(cond256_done),
    .in(cond256_in),
    .out(cond256_out),
    .reset(cond256_reset),
    .write_en(cond256_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire256 (
    .in(cond_wire256_in),
    .out(cond_wire256_out)
);
std_reg # (
    .WIDTH(1)
) cond257 (
    .clk(cond257_clk),
    .done(cond257_done),
    .in(cond257_in),
    .out(cond257_out),
    .reset(cond257_reset),
    .write_en(cond257_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire257 (
    .in(cond_wire257_in),
    .out(cond_wire257_out)
);
std_reg # (
    .WIDTH(1)
) cond258 (
    .clk(cond258_clk),
    .done(cond258_done),
    .in(cond258_in),
    .out(cond258_out),
    .reset(cond258_reset),
    .write_en(cond258_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire258 (
    .in(cond_wire258_in),
    .out(cond_wire258_out)
);
std_reg # (
    .WIDTH(1)
) cond259 (
    .clk(cond259_clk),
    .done(cond259_done),
    .in(cond259_in),
    .out(cond259_out),
    .reset(cond259_reset),
    .write_en(cond259_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire259 (
    .in(cond_wire259_in),
    .out(cond_wire259_out)
);
std_reg # (
    .WIDTH(1)
) cond260 (
    .clk(cond260_clk),
    .done(cond260_done),
    .in(cond260_in),
    .out(cond260_out),
    .reset(cond260_reset),
    .write_en(cond260_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire260 (
    .in(cond_wire260_in),
    .out(cond_wire260_out)
);
std_reg # (
    .WIDTH(1)
) cond261 (
    .clk(cond261_clk),
    .done(cond261_done),
    .in(cond261_in),
    .out(cond261_out),
    .reset(cond261_reset),
    .write_en(cond261_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire261 (
    .in(cond_wire261_in),
    .out(cond_wire261_out)
);
std_reg # (
    .WIDTH(1)
) cond262 (
    .clk(cond262_clk),
    .done(cond262_done),
    .in(cond262_in),
    .out(cond262_out),
    .reset(cond262_reset),
    .write_en(cond262_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire262 (
    .in(cond_wire262_in),
    .out(cond_wire262_out)
);
std_reg # (
    .WIDTH(1)
) cond263 (
    .clk(cond263_clk),
    .done(cond263_done),
    .in(cond263_in),
    .out(cond263_out),
    .reset(cond263_reset),
    .write_en(cond263_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire263 (
    .in(cond_wire263_in),
    .out(cond_wire263_out)
);
std_reg # (
    .WIDTH(1)
) cond264 (
    .clk(cond264_clk),
    .done(cond264_done),
    .in(cond264_in),
    .out(cond264_out),
    .reset(cond264_reset),
    .write_en(cond264_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire264 (
    .in(cond_wire264_in),
    .out(cond_wire264_out)
);
std_reg # (
    .WIDTH(1)
) cond265 (
    .clk(cond265_clk),
    .done(cond265_done),
    .in(cond265_in),
    .out(cond265_out),
    .reset(cond265_reset),
    .write_en(cond265_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire265 (
    .in(cond_wire265_in),
    .out(cond_wire265_out)
);
std_reg # (
    .WIDTH(1)
) cond266 (
    .clk(cond266_clk),
    .done(cond266_done),
    .in(cond266_in),
    .out(cond266_out),
    .reset(cond266_reset),
    .write_en(cond266_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire266 (
    .in(cond_wire266_in),
    .out(cond_wire266_out)
);
std_reg # (
    .WIDTH(1)
) cond267 (
    .clk(cond267_clk),
    .done(cond267_done),
    .in(cond267_in),
    .out(cond267_out),
    .reset(cond267_reset),
    .write_en(cond267_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire267 (
    .in(cond_wire267_in),
    .out(cond_wire267_out)
);
std_reg # (
    .WIDTH(1)
) cond268 (
    .clk(cond268_clk),
    .done(cond268_done),
    .in(cond268_in),
    .out(cond268_out),
    .reset(cond268_reset),
    .write_en(cond268_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire268 (
    .in(cond_wire268_in),
    .out(cond_wire268_out)
);
std_reg # (
    .WIDTH(1)
) fsm (
    .clk(fsm_clk),
    .done(fsm_done),
    .in(fsm_in),
    .out(fsm_out),
    .reset(fsm_reset),
    .write_en(fsm_write_en)
);
std_reg # (
    .WIDTH(5)
) fsm0 (
    .clk(fsm0_clk),
    .done(fsm0_done),
    .in(fsm0_in),
    .out(fsm0_out),
    .reset(fsm0_reset),
    .write_en(fsm0_write_en)
);
undef # (
    .WIDTH(1)
) ud (
    .out(ud_out)
);
std_add # (
    .WIDTH(5)
) adder (
    .left(adder_left),
    .out(adder_out),
    .right(adder_right)
);
undef # (
    .WIDTH(1)
) ud0 (
    .out(ud0_out)
);
std_add # (
    .WIDTH(1)
) adder0 (
    .left(adder0_left),
    .out(adder0_out),
    .right(adder0_right)
);
std_reg # (
    .WIDTH(1)
) signal_reg (
    .clk(signal_reg_clk),
    .done(signal_reg_done),
    .in(signal_reg_in),
    .out(signal_reg_out),
    .reset(signal_reg_reset),
    .write_en(signal_reg_write_en)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_seq_go (
    .in(early_reset_static_seq_go_in),
    .out(early_reset_static_seq_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_seq_done (
    .in(early_reset_static_seq_done_in),
    .out(early_reset_static_seq_done_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par0_go (
    .in(early_reset_static_par0_go_in),
    .out(early_reset_static_par0_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par0_done (
    .in(early_reset_static_par0_done_in),
    .out(early_reset_static_par0_done_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_seq_go (
    .in(wrapper_early_reset_static_seq_go_in),
    .out(wrapper_early_reset_static_seq_go_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_seq_done (
    .in(wrapper_early_reset_static_seq_done_in),
    .out(wrapper_early_reset_static_seq_done_out)
);
wire _guard0 = 1;
wire _guard1 = cond_wire58_out;
wire _guard2 = early_reset_static_par0_go_out;
wire _guard3 = _guard1 & _guard2;
wire _guard4 = cond_wire56_out;
wire _guard5 = early_reset_static_par0_go_out;
wire _guard6 = _guard4 & _guard5;
wire _guard7 = fsm_out == 1'd0;
wire _guard8 = cond_wire56_out;
wire _guard9 = _guard7 & _guard8;
wire _guard10 = fsm_out == 1'd0;
wire _guard11 = _guard9 & _guard10;
wire _guard12 = fsm_out == 1'd0;
wire _guard13 = cond_wire58_out;
wire _guard14 = _guard12 & _guard13;
wire _guard15 = fsm_out == 1'd0;
wire _guard16 = _guard14 & _guard15;
wire _guard17 = _guard11 | _guard16;
wire _guard18 = early_reset_static_par0_go_out;
wire _guard19 = _guard17 & _guard18;
wire _guard20 = fsm_out == 1'd0;
wire _guard21 = cond_wire56_out;
wire _guard22 = _guard20 & _guard21;
wire _guard23 = fsm_out == 1'd0;
wire _guard24 = _guard22 & _guard23;
wire _guard25 = fsm_out == 1'd0;
wire _guard26 = cond_wire58_out;
wire _guard27 = _guard25 & _guard26;
wire _guard28 = fsm_out == 1'd0;
wire _guard29 = _guard27 & _guard28;
wire _guard30 = _guard24 | _guard29;
wire _guard31 = early_reset_static_par0_go_out;
wire _guard32 = _guard30 & _guard31;
wire _guard33 = fsm_out == 1'd0;
wire _guard34 = cond_wire56_out;
wire _guard35 = _guard33 & _guard34;
wire _guard36 = fsm_out == 1'd0;
wire _guard37 = _guard35 & _guard36;
wire _guard38 = fsm_out == 1'd0;
wire _guard39 = cond_wire58_out;
wire _guard40 = _guard38 & _guard39;
wire _guard41 = fsm_out == 1'd0;
wire _guard42 = _guard40 & _guard41;
wire _guard43 = _guard37 | _guard42;
wire _guard44 = early_reset_static_par0_go_out;
wire _guard45 = _guard43 & _guard44;
wire _guard46 = cond_wire70_out;
wire _guard47 = early_reset_static_par0_go_out;
wire _guard48 = _guard46 & _guard47;
wire _guard49 = cond_wire68_out;
wire _guard50 = early_reset_static_par0_go_out;
wire _guard51 = _guard49 & _guard50;
wire _guard52 = fsm_out == 1'd0;
wire _guard53 = cond_wire68_out;
wire _guard54 = _guard52 & _guard53;
wire _guard55 = fsm_out == 1'd0;
wire _guard56 = _guard54 & _guard55;
wire _guard57 = fsm_out == 1'd0;
wire _guard58 = cond_wire70_out;
wire _guard59 = _guard57 & _guard58;
wire _guard60 = fsm_out == 1'd0;
wire _guard61 = _guard59 & _guard60;
wire _guard62 = _guard56 | _guard61;
wire _guard63 = early_reset_static_par0_go_out;
wire _guard64 = _guard62 & _guard63;
wire _guard65 = fsm_out == 1'd0;
wire _guard66 = cond_wire68_out;
wire _guard67 = _guard65 & _guard66;
wire _guard68 = fsm_out == 1'd0;
wire _guard69 = _guard67 & _guard68;
wire _guard70 = fsm_out == 1'd0;
wire _guard71 = cond_wire70_out;
wire _guard72 = _guard70 & _guard71;
wire _guard73 = fsm_out == 1'd0;
wire _guard74 = _guard72 & _guard73;
wire _guard75 = _guard69 | _guard74;
wire _guard76 = early_reset_static_par0_go_out;
wire _guard77 = _guard75 & _guard76;
wire _guard78 = fsm_out == 1'd0;
wire _guard79 = cond_wire68_out;
wire _guard80 = _guard78 & _guard79;
wire _guard81 = fsm_out == 1'd0;
wire _guard82 = _guard80 & _guard81;
wire _guard83 = fsm_out == 1'd0;
wire _guard84 = cond_wire70_out;
wire _guard85 = _guard83 & _guard84;
wire _guard86 = fsm_out == 1'd0;
wire _guard87 = _guard85 & _guard86;
wire _guard88 = _guard82 | _guard87;
wire _guard89 = early_reset_static_par0_go_out;
wire _guard90 = _guard88 & _guard89;
wire _guard91 = cond_wire57_out;
wire _guard92 = early_reset_static_par0_go_out;
wire _guard93 = _guard91 & _guard92;
wire _guard94 = cond_wire57_out;
wire _guard95 = early_reset_static_par0_go_out;
wire _guard96 = _guard94 & _guard95;
wire _guard97 = cond_wire86_out;
wire _guard98 = early_reset_static_par0_go_out;
wire _guard99 = _guard97 & _guard98;
wire _guard100 = cond_wire86_out;
wire _guard101 = early_reset_static_par0_go_out;
wire _guard102 = _guard100 & _guard101;
wire _guard103 = cond_wire94_out;
wire _guard104 = early_reset_static_par0_go_out;
wire _guard105 = _guard103 & _guard104;
wire _guard106 = cond_wire94_out;
wire _guard107 = early_reset_static_par0_go_out;
wire _guard108 = _guard106 & _guard107;
wire _guard109 = cond_wire98_out;
wire _guard110 = early_reset_static_par0_go_out;
wire _guard111 = _guard109 & _guard110;
wire _guard112 = cond_wire98_out;
wire _guard113 = early_reset_static_par0_go_out;
wire _guard114 = _guard112 & _guard113;
wire _guard115 = cond_wire138_out;
wire _guard116 = early_reset_static_par0_go_out;
wire _guard117 = _guard115 & _guard116;
wire _guard118 = cond_wire138_out;
wire _guard119 = early_reset_static_par0_go_out;
wire _guard120 = _guard118 & _guard119;
wire _guard121 = cond_wire123_out;
wire _guard122 = early_reset_static_par0_go_out;
wire _guard123 = _guard121 & _guard122;
wire _guard124 = cond_wire123_out;
wire _guard125 = early_reset_static_par0_go_out;
wire _guard126 = _guard124 & _guard125;
wire _guard127 = cond_wire182_out;
wire _guard128 = early_reset_static_par0_go_out;
wire _guard129 = _guard127 & _guard128;
wire _guard130 = cond_wire180_out;
wire _guard131 = early_reset_static_par0_go_out;
wire _guard132 = _guard130 & _guard131;
wire _guard133 = fsm_out == 1'd0;
wire _guard134 = cond_wire180_out;
wire _guard135 = _guard133 & _guard134;
wire _guard136 = fsm_out == 1'd0;
wire _guard137 = _guard135 & _guard136;
wire _guard138 = fsm_out == 1'd0;
wire _guard139 = cond_wire182_out;
wire _guard140 = _guard138 & _guard139;
wire _guard141 = fsm_out == 1'd0;
wire _guard142 = _guard140 & _guard141;
wire _guard143 = _guard137 | _guard142;
wire _guard144 = early_reset_static_par0_go_out;
wire _guard145 = _guard143 & _guard144;
wire _guard146 = fsm_out == 1'd0;
wire _guard147 = cond_wire180_out;
wire _guard148 = _guard146 & _guard147;
wire _guard149 = fsm_out == 1'd0;
wire _guard150 = _guard148 & _guard149;
wire _guard151 = fsm_out == 1'd0;
wire _guard152 = cond_wire182_out;
wire _guard153 = _guard151 & _guard152;
wire _guard154 = fsm_out == 1'd0;
wire _guard155 = _guard153 & _guard154;
wire _guard156 = _guard150 | _guard155;
wire _guard157 = early_reset_static_par0_go_out;
wire _guard158 = _guard156 & _guard157;
wire _guard159 = fsm_out == 1'd0;
wire _guard160 = cond_wire180_out;
wire _guard161 = _guard159 & _guard160;
wire _guard162 = fsm_out == 1'd0;
wire _guard163 = _guard161 & _guard162;
wire _guard164 = fsm_out == 1'd0;
wire _guard165 = cond_wire182_out;
wire _guard166 = _guard164 & _guard165;
wire _guard167 = fsm_out == 1'd0;
wire _guard168 = _guard166 & _guard167;
wire _guard169 = _guard163 | _guard168;
wire _guard170 = early_reset_static_par0_go_out;
wire _guard171 = _guard169 & _guard170;
wire _guard172 = cond_wire177_out;
wire _guard173 = early_reset_static_par0_go_out;
wire _guard174 = _guard172 & _guard173;
wire _guard175 = cond_wire177_out;
wire _guard176 = early_reset_static_par0_go_out;
wire _guard177 = _guard175 & _guard176;
wire _guard178 = cond_wire210_out;
wire _guard179 = early_reset_static_par0_go_out;
wire _guard180 = _guard178 & _guard179;
wire _guard181 = cond_wire210_out;
wire _guard182 = early_reset_static_par0_go_out;
wire _guard183 = _guard181 & _guard182;
wire _guard184 = cond_wire185_out;
wire _guard185 = early_reset_static_par0_go_out;
wire _guard186 = _guard184 & _guard185;
wire _guard187 = cond_wire185_out;
wire _guard188 = early_reset_static_par0_go_out;
wire _guard189 = _guard187 & _guard188;
wire _guard190 = cond_wire218_out;
wire _guard191 = early_reset_static_par0_go_out;
wire _guard192 = _guard190 & _guard191;
wire _guard193 = cond_wire218_out;
wire _guard194 = early_reset_static_par0_go_out;
wire _guard195 = _guard193 & _guard194;
wire _guard196 = cond_wire206_out;
wire _guard197 = early_reset_static_par0_go_out;
wire _guard198 = _guard196 & _guard197;
wire _guard199 = cond_wire206_out;
wire _guard200 = early_reset_static_par0_go_out;
wire _guard201 = _guard199 & _guard200;
wire _guard202 = cond_wire14_out;
wire _guard203 = early_reset_static_par0_go_out;
wire _guard204 = _guard202 & _guard203;
wire _guard205 = cond_wire14_out;
wire _guard206 = early_reset_static_par0_go_out;
wire _guard207 = _guard205 & _guard206;
wire _guard208 = cond_wire39_out;
wire _guard209 = early_reset_static_par0_go_out;
wire _guard210 = _guard208 & _guard209;
wire _guard211 = cond_wire39_out;
wire _guard212 = early_reset_static_par0_go_out;
wire _guard213 = _guard211 & _guard212;
wire _guard214 = early_reset_static_par0_go_out;
wire _guard215 = early_reset_static_par0_go_out;
wire _guard216 = fsm0_out == 5'd0;
wire _guard217 = early_reset_static_seq_go_out;
wire _guard218 = _guard216 & _guard217;
wire _guard219 = early_reset_static_par0_go_out;
wire _guard220 = _guard218 | _guard219;
wire _guard221 = early_reset_static_par0_go_out;
wire _guard222 = fsm0_out == 5'd0;
wire _guard223 = early_reset_static_seq_go_out;
wire _guard224 = _guard222 & _guard223;
wire _guard225 = early_reset_static_par0_go_out;
wire _guard226 = early_reset_static_par0_go_out;
wire _guard227 = early_reset_static_par0_go_out;
wire _guard228 = early_reset_static_par0_go_out;
wire _guard229 = fsm0_out == 5'd0;
wire _guard230 = early_reset_static_seq_go_out;
wire _guard231 = _guard229 & _guard230;
wire _guard232 = early_reset_static_par0_go_out;
wire _guard233 = _guard231 | _guard232;
wire _guard234 = fsm0_out == 5'd0;
wire _guard235 = early_reset_static_seq_go_out;
wire _guard236 = _guard234 & _guard235;
wire _guard237 = early_reset_static_par0_go_out;
wire _guard238 = early_reset_static_par0_go_out;
wire _guard239 = early_reset_static_par0_go_out;
wire _guard240 = fsm0_out == 5'd0;
wire _guard241 = early_reset_static_seq_go_out;
wire _guard242 = _guard240 & _guard241;
wire _guard243 = early_reset_static_par0_go_out;
wire _guard244 = _guard242 | _guard243;
wire _guard245 = early_reset_static_par0_go_out;
wire _guard246 = fsm0_out == 5'd0;
wire _guard247 = early_reset_static_seq_go_out;
wire _guard248 = _guard246 & _guard247;
wire _guard249 = early_reset_static_par0_go_out;
wire _guard250 = early_reset_static_par0_go_out;
wire _guard251 = early_reset_static_par0_go_out;
wire _guard252 = early_reset_static_par0_go_out;
wire _guard253 = early_reset_static_par0_go_out;
wire _guard254 = ~_guard0;
wire _guard255 = early_reset_static_par0_go_out;
wire _guard256 = _guard254 & _guard255;
wire _guard257 = ~_guard0;
wire _guard258 = early_reset_static_par0_go_out;
wire _guard259 = _guard257 & _guard258;
wire _guard260 = early_reset_static_par0_go_out;
wire _guard261 = early_reset_static_par0_go_out;
wire _guard262 = ~_guard0;
wire _guard263 = early_reset_static_par0_go_out;
wire _guard264 = _guard262 & _guard263;
wire _guard265 = ~_guard0;
wire _guard266 = early_reset_static_par0_go_out;
wire _guard267 = _guard265 & _guard266;
wire _guard268 = early_reset_static_par0_go_out;
wire _guard269 = early_reset_static_par0_go_out;
wire _guard270 = ~_guard0;
wire _guard271 = early_reset_static_par0_go_out;
wire _guard272 = _guard270 & _guard271;
wire _guard273 = early_reset_static_par0_go_out;
wire _guard274 = early_reset_static_par0_go_out;
wire _guard275 = ~_guard0;
wire _guard276 = early_reset_static_par0_go_out;
wire _guard277 = _guard275 & _guard276;
wire _guard278 = early_reset_static_par0_go_out;
wire _guard279 = early_reset_static_par0_go_out;
wire _guard280 = early_reset_static_par0_go_out;
wire _guard281 = early_reset_static_par0_go_out;
wire _guard282 = early_reset_static_par0_go_out;
wire _guard283 = early_reset_static_par0_go_out;
wire _guard284 = early_reset_static_par0_go_out;
wire _guard285 = early_reset_static_par0_go_out;
wire _guard286 = ~_guard0;
wire _guard287 = early_reset_static_par0_go_out;
wire _guard288 = _guard286 & _guard287;
wire _guard289 = early_reset_static_par0_go_out;
wire _guard290 = ~_guard0;
wire _guard291 = early_reset_static_par0_go_out;
wire _guard292 = _guard290 & _guard291;
wire _guard293 = ~_guard0;
wire _guard294 = early_reset_static_par0_go_out;
wire _guard295 = _guard293 & _guard294;
wire _guard296 = early_reset_static_par0_go_out;
wire _guard297 = ~_guard0;
wire _guard298 = early_reset_static_par0_go_out;
wire _guard299 = _guard297 & _guard298;
wire _guard300 = early_reset_static_par0_go_out;
wire _guard301 = early_reset_static_par0_go_out;
wire _guard302 = ~_guard0;
wire _guard303 = early_reset_static_par0_go_out;
wire _guard304 = _guard302 & _guard303;
wire _guard305 = early_reset_static_par0_go_out;
wire _guard306 = early_reset_static_par0_go_out;
wire _guard307 = early_reset_static_par0_go_out;
wire _guard308 = early_reset_static_par0_go_out;
wire _guard309 = ~_guard0;
wire _guard310 = early_reset_static_par0_go_out;
wire _guard311 = _guard309 & _guard310;
wire _guard312 = early_reset_static_par0_go_out;
wire _guard313 = early_reset_static_par0_go_out;
wire _guard314 = ~_guard0;
wire _guard315 = early_reset_static_par0_go_out;
wire _guard316 = _guard314 & _guard315;
wire _guard317 = early_reset_static_par0_go_out;
wire _guard318 = early_reset_static_par0_go_out;
wire _guard319 = early_reset_static_par0_go_out;
wire _guard320 = ~_guard0;
wire _guard321 = early_reset_static_par0_go_out;
wire _guard322 = _guard320 & _guard321;
wire _guard323 = early_reset_static_par0_go_out;
wire _guard324 = ~_guard0;
wire _guard325 = early_reset_static_par0_go_out;
wire _guard326 = _guard324 & _guard325;
wire _guard327 = early_reset_static_par0_go_out;
wire _guard328 = early_reset_static_par0_go_out;
wire _guard329 = early_reset_static_par0_go_out;
wire _guard330 = early_reset_static_par0_go_out;
wire _guard331 = early_reset_static_par0_go_out;
wire _guard332 = ~_guard0;
wire _guard333 = early_reset_static_par0_go_out;
wire _guard334 = _guard332 & _guard333;
wire _guard335 = early_reset_static_par0_go_out;
wire _guard336 = early_reset_static_par0_go_out;
wire _guard337 = ~_guard0;
wire _guard338 = early_reset_static_par0_go_out;
wire _guard339 = _guard337 & _guard338;
wire _guard340 = early_reset_static_par0_go_out;
wire _guard341 = early_reset_static_par0_go_out;
wire _guard342 = early_reset_static_par0_go_out;
wire _guard343 = cond_wire11_out;
wire _guard344 = early_reset_static_par0_go_out;
wire _guard345 = _guard343 & _guard344;
wire _guard346 = cond_wire11_out;
wire _guard347 = early_reset_static_par0_go_out;
wire _guard348 = _guard346 & _guard347;
wire _guard349 = cond_wire16_out;
wire _guard350 = early_reset_static_par0_go_out;
wire _guard351 = _guard349 & _guard350;
wire _guard352 = cond_wire16_out;
wire _guard353 = early_reset_static_par0_go_out;
wire _guard354 = _guard352 & _guard353;
wire _guard355 = cond_wire1_out;
wire _guard356 = early_reset_static_par0_go_out;
wire _guard357 = _guard355 & _guard356;
wire _guard358 = cond_wire1_out;
wire _guard359 = early_reset_static_par0_go_out;
wire _guard360 = _guard358 & _guard359;
wire _guard361 = cond_wire50_out;
wire _guard362 = early_reset_static_par0_go_out;
wire _guard363 = _guard361 & _guard362;
wire _guard364 = cond_wire48_out;
wire _guard365 = early_reset_static_par0_go_out;
wire _guard366 = _guard364 & _guard365;
wire _guard367 = fsm_out == 1'd0;
wire _guard368 = cond_wire48_out;
wire _guard369 = _guard367 & _guard368;
wire _guard370 = fsm_out == 1'd0;
wire _guard371 = _guard369 & _guard370;
wire _guard372 = fsm_out == 1'd0;
wire _guard373 = cond_wire50_out;
wire _guard374 = _guard372 & _guard373;
wire _guard375 = fsm_out == 1'd0;
wire _guard376 = _guard374 & _guard375;
wire _guard377 = _guard371 | _guard376;
wire _guard378 = early_reset_static_par0_go_out;
wire _guard379 = _guard377 & _guard378;
wire _guard380 = fsm_out == 1'd0;
wire _guard381 = cond_wire48_out;
wire _guard382 = _guard380 & _guard381;
wire _guard383 = fsm_out == 1'd0;
wire _guard384 = _guard382 & _guard383;
wire _guard385 = fsm_out == 1'd0;
wire _guard386 = cond_wire50_out;
wire _guard387 = _guard385 & _guard386;
wire _guard388 = fsm_out == 1'd0;
wire _guard389 = _guard387 & _guard388;
wire _guard390 = _guard384 | _guard389;
wire _guard391 = early_reset_static_par0_go_out;
wire _guard392 = _guard390 & _guard391;
wire _guard393 = fsm_out == 1'd0;
wire _guard394 = cond_wire48_out;
wire _guard395 = _guard393 & _guard394;
wire _guard396 = fsm_out == 1'd0;
wire _guard397 = _guard395 & _guard396;
wire _guard398 = fsm_out == 1'd0;
wire _guard399 = cond_wire50_out;
wire _guard400 = _guard398 & _guard399;
wire _guard401 = fsm_out == 1'd0;
wire _guard402 = _guard400 & _guard401;
wire _guard403 = _guard397 | _guard402;
wire _guard404 = early_reset_static_par0_go_out;
wire _guard405 = _guard403 & _guard404;
wire _guard406 = cond_wire54_out;
wire _guard407 = early_reset_static_par0_go_out;
wire _guard408 = _guard406 & _guard407;
wire _guard409 = cond_wire52_out;
wire _guard410 = early_reset_static_par0_go_out;
wire _guard411 = _guard409 & _guard410;
wire _guard412 = fsm_out == 1'd0;
wire _guard413 = cond_wire52_out;
wire _guard414 = _guard412 & _guard413;
wire _guard415 = fsm_out == 1'd0;
wire _guard416 = _guard414 & _guard415;
wire _guard417 = fsm_out == 1'd0;
wire _guard418 = cond_wire54_out;
wire _guard419 = _guard417 & _guard418;
wire _guard420 = fsm_out == 1'd0;
wire _guard421 = _guard419 & _guard420;
wire _guard422 = _guard416 | _guard421;
wire _guard423 = early_reset_static_par0_go_out;
wire _guard424 = _guard422 & _guard423;
wire _guard425 = fsm_out == 1'd0;
wire _guard426 = cond_wire52_out;
wire _guard427 = _guard425 & _guard426;
wire _guard428 = fsm_out == 1'd0;
wire _guard429 = _guard427 & _guard428;
wire _guard430 = fsm_out == 1'd0;
wire _guard431 = cond_wire54_out;
wire _guard432 = _guard430 & _guard431;
wire _guard433 = fsm_out == 1'd0;
wire _guard434 = _guard432 & _guard433;
wire _guard435 = _guard429 | _guard434;
wire _guard436 = early_reset_static_par0_go_out;
wire _guard437 = _guard435 & _guard436;
wire _guard438 = fsm_out == 1'd0;
wire _guard439 = cond_wire52_out;
wire _guard440 = _guard438 & _guard439;
wire _guard441 = fsm_out == 1'd0;
wire _guard442 = _guard440 & _guard441;
wire _guard443 = fsm_out == 1'd0;
wire _guard444 = cond_wire54_out;
wire _guard445 = _guard443 & _guard444;
wire _guard446 = fsm_out == 1'd0;
wire _guard447 = _guard445 & _guard446;
wire _guard448 = _guard442 | _guard447;
wire _guard449 = early_reset_static_par0_go_out;
wire _guard450 = _guard448 & _guard449;
wire _guard451 = cond_wire49_out;
wire _guard452 = early_reset_static_par0_go_out;
wire _guard453 = _guard451 & _guard452;
wire _guard454 = cond_wire49_out;
wire _guard455 = early_reset_static_par0_go_out;
wire _guard456 = _guard454 & _guard455;
wire _guard457 = cond_wire94_out;
wire _guard458 = early_reset_static_par0_go_out;
wire _guard459 = _guard457 & _guard458;
wire _guard460 = cond_wire94_out;
wire _guard461 = early_reset_static_par0_go_out;
wire _guard462 = _guard460 & _guard461;
wire _guard463 = cond_wire135_out;
wire _guard464 = early_reset_static_par0_go_out;
wire _guard465 = _guard463 & _guard464;
wire _guard466 = cond_wire135_out;
wire _guard467 = early_reset_static_par0_go_out;
wire _guard468 = _guard466 & _guard467;
wire _guard469 = cond_wire173_out;
wire _guard470 = early_reset_static_par0_go_out;
wire _guard471 = _guard469 & _guard470;
wire _guard472 = cond_wire173_out;
wire _guard473 = early_reset_static_par0_go_out;
wire _guard474 = _guard472 & _guard473;
wire _guard475 = cond_wire181_out;
wire _guard476 = early_reset_static_par0_go_out;
wire _guard477 = _guard475 & _guard476;
wire _guard478 = cond_wire181_out;
wire _guard479 = early_reset_static_par0_go_out;
wire _guard480 = _guard478 & _guard479;
wire _guard481 = cond_wire223_out;
wire _guard482 = early_reset_static_par0_go_out;
wire _guard483 = _guard481 & _guard482;
wire _guard484 = cond_wire221_out;
wire _guard485 = early_reset_static_par0_go_out;
wire _guard486 = _guard484 & _guard485;
wire _guard487 = fsm_out == 1'd0;
wire _guard488 = cond_wire221_out;
wire _guard489 = _guard487 & _guard488;
wire _guard490 = fsm_out == 1'd0;
wire _guard491 = _guard489 & _guard490;
wire _guard492 = fsm_out == 1'd0;
wire _guard493 = cond_wire223_out;
wire _guard494 = _guard492 & _guard493;
wire _guard495 = fsm_out == 1'd0;
wire _guard496 = _guard494 & _guard495;
wire _guard497 = _guard491 | _guard496;
wire _guard498 = early_reset_static_par0_go_out;
wire _guard499 = _guard497 & _guard498;
wire _guard500 = fsm_out == 1'd0;
wire _guard501 = cond_wire221_out;
wire _guard502 = _guard500 & _guard501;
wire _guard503 = fsm_out == 1'd0;
wire _guard504 = _guard502 & _guard503;
wire _guard505 = fsm_out == 1'd0;
wire _guard506 = cond_wire223_out;
wire _guard507 = _guard505 & _guard506;
wire _guard508 = fsm_out == 1'd0;
wire _guard509 = _guard507 & _guard508;
wire _guard510 = _guard504 | _guard509;
wire _guard511 = early_reset_static_par0_go_out;
wire _guard512 = _guard510 & _guard511;
wire _guard513 = fsm_out == 1'd0;
wire _guard514 = cond_wire221_out;
wire _guard515 = _guard513 & _guard514;
wire _guard516 = fsm_out == 1'd0;
wire _guard517 = _guard515 & _guard516;
wire _guard518 = fsm_out == 1'd0;
wire _guard519 = cond_wire223_out;
wire _guard520 = _guard518 & _guard519;
wire _guard521 = fsm_out == 1'd0;
wire _guard522 = _guard520 & _guard521;
wire _guard523 = _guard517 | _guard522;
wire _guard524 = early_reset_static_par0_go_out;
wire _guard525 = _guard523 & _guard524;
wire _guard526 = cond_wire201_out;
wire _guard527 = early_reset_static_par0_go_out;
wire _guard528 = _guard526 & _guard527;
wire _guard529 = cond_wire201_out;
wire _guard530 = early_reset_static_par0_go_out;
wire _guard531 = _guard529 & _guard530;
wire _guard532 = cond_wire252_out;
wire _guard533 = early_reset_static_par0_go_out;
wire _guard534 = _guard532 & _guard533;
wire _guard535 = cond_wire250_out;
wire _guard536 = early_reset_static_par0_go_out;
wire _guard537 = _guard535 & _guard536;
wire _guard538 = fsm_out == 1'd0;
wire _guard539 = cond_wire250_out;
wire _guard540 = _guard538 & _guard539;
wire _guard541 = fsm_out == 1'd0;
wire _guard542 = _guard540 & _guard541;
wire _guard543 = fsm_out == 1'd0;
wire _guard544 = cond_wire252_out;
wire _guard545 = _guard543 & _guard544;
wire _guard546 = fsm_out == 1'd0;
wire _guard547 = _guard545 & _guard546;
wire _guard548 = _guard542 | _guard547;
wire _guard549 = early_reset_static_par0_go_out;
wire _guard550 = _guard548 & _guard549;
wire _guard551 = fsm_out == 1'd0;
wire _guard552 = cond_wire250_out;
wire _guard553 = _guard551 & _guard552;
wire _guard554 = fsm_out == 1'd0;
wire _guard555 = _guard553 & _guard554;
wire _guard556 = fsm_out == 1'd0;
wire _guard557 = cond_wire252_out;
wire _guard558 = _guard556 & _guard557;
wire _guard559 = fsm_out == 1'd0;
wire _guard560 = _guard558 & _guard559;
wire _guard561 = _guard555 | _guard560;
wire _guard562 = early_reset_static_par0_go_out;
wire _guard563 = _guard561 & _guard562;
wire _guard564 = fsm_out == 1'd0;
wire _guard565 = cond_wire250_out;
wire _guard566 = _guard564 & _guard565;
wire _guard567 = fsm_out == 1'd0;
wire _guard568 = _guard566 & _guard567;
wire _guard569 = fsm_out == 1'd0;
wire _guard570 = cond_wire252_out;
wire _guard571 = _guard569 & _guard570;
wire _guard572 = fsm_out == 1'd0;
wire _guard573 = _guard571 & _guard572;
wire _guard574 = _guard568 | _guard573;
wire _guard575 = early_reset_static_par0_go_out;
wire _guard576 = _guard574 & _guard575;
wire _guard577 = cond_wire251_out;
wire _guard578 = early_reset_static_par0_go_out;
wire _guard579 = _guard577 & _guard578;
wire _guard580 = cond_wire251_out;
wire _guard581 = early_reset_static_par0_go_out;
wire _guard582 = _guard580 & _guard581;
wire _guard583 = cond_wire259_out;
wire _guard584 = early_reset_static_par0_go_out;
wire _guard585 = _guard583 & _guard584;
wire _guard586 = cond_wire259_out;
wire _guard587 = early_reset_static_par0_go_out;
wire _guard588 = _guard586 & _guard587;
wire _guard589 = cond_wire234_out;
wire _guard590 = early_reset_static_par0_go_out;
wire _guard591 = _guard589 & _guard590;
wire _guard592 = cond_wire234_out;
wire _guard593 = early_reset_static_par0_go_out;
wire _guard594 = _guard592 & _guard593;
wire _guard595 = fsm0_out == 5'd0;
wire _guard596 = early_reset_static_seq_go_out;
wire _guard597 = _guard595 & _guard596;
wire _guard598 = cond_wire105_out;
wire _guard599 = early_reset_static_par0_go_out;
wire _guard600 = _guard598 & _guard599;
wire _guard601 = _guard597 | _guard600;
wire _guard602 = cond_wire105_out;
wire _guard603 = early_reset_static_par0_go_out;
wire _guard604 = _guard602 & _guard603;
wire _guard605 = fsm0_out == 5'd0;
wire _guard606 = early_reset_static_seq_go_out;
wire _guard607 = _guard605 & _guard606;
wire _guard608 = fsm0_out == 5'd0;
wire _guard609 = early_reset_static_seq_go_out;
wire _guard610 = _guard608 & _guard609;
wire _guard611 = cond_wire237_out;
wire _guard612 = early_reset_static_par0_go_out;
wire _guard613 = _guard611 & _guard612;
wire _guard614 = _guard610 | _guard613;
wire _guard615 = fsm0_out == 5'd0;
wire _guard616 = early_reset_static_seq_go_out;
wire _guard617 = _guard615 & _guard616;
wire _guard618 = cond_wire237_out;
wire _guard619 = early_reset_static_par0_go_out;
wire _guard620 = _guard618 & _guard619;
wire _guard621 = fsm0_out == 5'd0;
wire _guard622 = early_reset_static_seq_go_out;
wire _guard623 = _guard621 & _guard622;
wire _guard624 = early_reset_static_par0_go_out;
wire _guard625 = _guard623 | _guard624;
wire _guard626 = early_reset_static_par0_go_out;
wire _guard627 = fsm0_out == 5'd0;
wire _guard628 = early_reset_static_seq_go_out;
wire _guard629 = _guard627 & _guard628;
wire _guard630 = early_reset_static_par0_go_out;
wire _guard631 = early_reset_static_par0_go_out;
wire _guard632 = early_reset_static_par0_go_out;
wire _guard633 = early_reset_static_par0_go_out;
wire _guard634 = early_reset_static_par0_go_out;
wire _guard635 = early_reset_static_par0_go_out;
wire _guard636 = early_reset_static_par0_go_out;
wire _guard637 = early_reset_static_par0_go_out;
wire _guard638 = fsm0_out == 5'd0;
wire _guard639 = early_reset_static_seq_go_out;
wire _guard640 = _guard638 & _guard639;
wire _guard641 = early_reset_static_par0_go_out;
wire _guard642 = _guard640 | _guard641;
wire _guard643 = fsm0_out == 5'd0;
wire _guard644 = early_reset_static_seq_go_out;
wire _guard645 = _guard643 & _guard644;
wire _guard646 = early_reset_static_par0_go_out;
wire _guard647 = fsm0_out == 5'd0;
wire _guard648 = early_reset_static_seq_go_out;
wire _guard649 = _guard647 & _guard648;
wire _guard650 = early_reset_static_par0_go_out;
wire _guard651 = _guard649 | _guard650;
wire _guard652 = early_reset_static_par0_go_out;
wire _guard653 = fsm0_out == 5'd0;
wire _guard654 = early_reset_static_seq_go_out;
wire _guard655 = _guard653 & _guard654;
wire _guard656 = fsm0_out == 5'd0;
wire _guard657 = early_reset_static_seq_go_out;
wire _guard658 = _guard656 & _guard657;
wire _guard659 = early_reset_static_par0_go_out;
wire _guard660 = _guard658 | _guard659;
wire _guard661 = early_reset_static_par0_go_out;
wire _guard662 = fsm0_out == 5'd0;
wire _guard663 = early_reset_static_seq_go_out;
wire _guard664 = _guard662 & _guard663;
wire _guard665 = fsm0_out == 5'd0;
wire _guard666 = early_reset_static_seq_go_out;
wire _guard667 = _guard665 & _guard666;
wire _guard668 = early_reset_static_par0_go_out;
wire _guard669 = _guard667 | _guard668;
wire _guard670 = fsm0_out == 5'd0;
wire _guard671 = early_reset_static_seq_go_out;
wire _guard672 = _guard670 & _guard671;
wire _guard673 = early_reset_static_par0_go_out;
wire _guard674 = wrapper_early_reset_static_seq_done_out;
wire _guard675 = cond_wire9_out;
wire _guard676 = early_reset_static_par0_go_out;
wire _guard677 = _guard675 & _guard676;
wire _guard678 = cond_wire142_out;
wire _guard679 = early_reset_static_par0_go_out;
wire _guard680 = _guard678 & _guard679;
wire _guard681 = cond_wire162_out;
wire _guard682 = early_reset_static_par0_go_out;
wire _guard683 = _guard681 & _guard682;
wire _guard684 = cond_wire166_out;
wire _guard685 = early_reset_static_par0_go_out;
wire _guard686 = _guard684 & _guard685;
wire _guard687 = cond_wire150_out;
wire _guard688 = early_reset_static_par0_go_out;
wire _guard689 = _guard687 & _guard688;
wire _guard690 = cond_wire158_out;
wire _guard691 = early_reset_static_par0_go_out;
wire _guard692 = _guard690 & _guard691;
wire _guard693 = cond_wire170_out;
wire _guard694 = early_reset_static_par0_go_out;
wire _guard695 = _guard693 & _guard694;
wire _guard696 = cond_wire154_out;
wire _guard697 = early_reset_static_par0_go_out;
wire _guard698 = _guard696 & _guard697;
wire _guard699 = cond_wire146_out;
wire _guard700 = early_reset_static_par0_go_out;
wire _guard701 = _guard699 & _guard700;
wire _guard702 = cond_wire171_out;
wire _guard703 = early_reset_static_par0_go_out;
wire _guard704 = _guard702 & _guard703;
wire _guard705 = cond_wire_out;
wire _guard706 = early_reset_static_par0_go_out;
wire _guard707 = _guard705 & _guard706;
wire _guard708 = cond_wire55_out;
wire _guard709 = early_reset_static_par0_go_out;
wire _guard710 = _guard708 & _guard709;
wire _guard711 = cond_wire63_out;
wire _guard712 = early_reset_static_par0_go_out;
wire _guard713 = _guard711 & _guard712;
wire _guard714 = cond_wire59_out;
wire _guard715 = early_reset_static_par0_go_out;
wire _guard716 = _guard714 & _guard715;
wire _guard717 = cond_wire43_out;
wire _guard718 = early_reset_static_par0_go_out;
wire _guard719 = _guard717 & _guard718;
wire _guard720 = cond_wire71_out;
wire _guard721 = early_reset_static_par0_go_out;
wire _guard722 = _guard720 & _guard721;
wire _guard723 = cond_wire51_out;
wire _guard724 = early_reset_static_par0_go_out;
wire _guard725 = _guard723 & _guard724;
wire _guard726 = cond_wire67_out;
wire _guard727 = early_reset_static_par0_go_out;
wire _guard728 = _guard726 & _guard727;
wire _guard729 = cond_wire47_out;
wire _guard730 = early_reset_static_par0_go_out;
wire _guard731 = _guard729 & _guard730;
wire _guard732 = cond_wire187_out;
wire _guard733 = early_reset_static_par0_go_out;
wire _guard734 = _guard732 & _guard733;
wire _guard735 = cond_wire195_out;
wire _guard736 = early_reset_static_par0_go_out;
wire _guard737 = _guard735 & _guard736;
wire _guard738 = cond_wire191_out;
wire _guard739 = early_reset_static_par0_go_out;
wire _guard740 = _guard738 & _guard739;
wire _guard741 = cond_wire175_out;
wire _guard742 = early_reset_static_par0_go_out;
wire _guard743 = _guard741 & _guard742;
wire _guard744 = cond_wire203_out;
wire _guard745 = early_reset_static_par0_go_out;
wire _guard746 = _guard744 & _guard745;
wire _guard747 = cond_wire183_out;
wire _guard748 = early_reset_static_par0_go_out;
wire _guard749 = _guard747 & _guard748;
wire _guard750 = cond_wire199_out;
wire _guard751 = early_reset_static_par0_go_out;
wire _guard752 = _guard750 & _guard751;
wire _guard753 = cond_wire179_out;
wire _guard754 = early_reset_static_par0_go_out;
wire _guard755 = _guard753 & _guard754;
wire _guard756 = cond_wire183_out;
wire _guard757 = early_reset_static_par0_go_out;
wire _guard758 = _guard756 & _guard757;
wire _guard759 = cond_wire175_out;
wire _guard760 = early_reset_static_par0_go_out;
wire _guard761 = _guard759 & _guard760;
wire _guard762 = cond_wire191_out;
wire _guard763 = early_reset_static_par0_go_out;
wire _guard764 = _guard762 & _guard763;
wire _guard765 = cond_wire179_out;
wire _guard766 = early_reset_static_par0_go_out;
wire _guard767 = _guard765 & _guard766;
wire _guard768 = cond_wire203_out;
wire _guard769 = early_reset_static_par0_go_out;
wire _guard770 = _guard768 & _guard769;
wire _guard771 = cond_wire187_out;
wire _guard772 = early_reset_static_par0_go_out;
wire _guard773 = _guard771 & _guard772;
wire _guard774 = cond_wire195_out;
wire _guard775 = early_reset_static_par0_go_out;
wire _guard776 = _guard774 & _guard775;
wire _guard777 = cond_wire199_out;
wire _guard778 = early_reset_static_par0_go_out;
wire _guard779 = _guard777 & _guard778;
wire _guard780 = cond_wire204_out;
wire _guard781 = early_reset_static_par0_go_out;
wire _guard782 = _guard780 & _guard781;
wire _guard783 = cond_wire8_out;
wire _guard784 = early_reset_static_par0_go_out;
wire _guard785 = _guard783 & _guard784;
wire _guard786 = cond_wire38_out;
wire _guard787 = early_reset_static_par0_go_out;
wire _guard788 = _guard786 & _guard787;
wire _guard789 = cond_wire18_out;
wire _guard790 = early_reset_static_par0_go_out;
wire _guard791 = _guard789 & _guard790;
wire _guard792 = cond_wire28_out;
wire _guard793 = early_reset_static_par0_go_out;
wire _guard794 = _guard792 & _guard793;
wire _guard795 = cond_wire13_out;
wire _guard796 = early_reset_static_par0_go_out;
wire _guard797 = _guard795 & _guard796;
wire _guard798 = cond_wire23_out;
wire _guard799 = early_reset_static_par0_go_out;
wire _guard800 = _guard798 & _guard799;
wire _guard801 = cond_wire3_out;
wire _guard802 = early_reset_static_par0_go_out;
wire _guard803 = _guard801 & _guard802;
wire _guard804 = cond_wire33_out;
wire _guard805 = early_reset_static_par0_go_out;
wire _guard806 = _guard804 & _guard805;
wire _guard807 = cond_wire220_out;
wire _guard808 = early_reset_static_par0_go_out;
wire _guard809 = _guard807 & _guard808;
wire _guard810 = cond_wire228_out;
wire _guard811 = early_reset_static_par0_go_out;
wire _guard812 = _guard810 & _guard811;
wire _guard813 = cond_wire224_out;
wire _guard814 = early_reset_static_par0_go_out;
wire _guard815 = _guard813 & _guard814;
wire _guard816 = cond_wire208_out;
wire _guard817 = early_reset_static_par0_go_out;
wire _guard818 = _guard816 & _guard817;
wire _guard819 = cond_wire236_out;
wire _guard820 = early_reset_static_par0_go_out;
wire _guard821 = _guard819 & _guard820;
wire _guard822 = cond_wire216_out;
wire _guard823 = early_reset_static_par0_go_out;
wire _guard824 = _guard822 & _guard823;
wire _guard825 = cond_wire232_out;
wire _guard826 = early_reset_static_par0_go_out;
wire _guard827 = _guard825 & _guard826;
wire _guard828 = cond_wire212_out;
wire _guard829 = early_reset_static_par0_go_out;
wire _guard830 = _guard828 & _guard829;
wire _guard831 = cond_wire125_out;
wire _guard832 = early_reset_static_par0_go_out;
wire _guard833 = _guard831 & _guard832;
wire _guard834 = cond_wire137_out;
wire _guard835 = early_reset_static_par0_go_out;
wire _guard836 = _guard834 & _guard835;
wire _guard837 = cond_wire117_out;
wire _guard838 = early_reset_static_par0_go_out;
wire _guard839 = _guard837 & _guard838;
wire _guard840 = cond_wire129_out;
wire _guard841 = early_reset_static_par0_go_out;
wire _guard842 = _guard840 & _guard841;
wire _guard843 = cond_wire133_out;
wire _guard844 = early_reset_static_par0_go_out;
wire _guard845 = _guard843 & _guard844;
wire _guard846 = cond_wire109_out;
wire _guard847 = early_reset_static_par0_go_out;
wire _guard848 = _guard846 & _guard847;
wire _guard849 = cond_wire113_out;
wire _guard850 = early_reset_static_par0_go_out;
wire _guard851 = _guard849 & _guard850;
wire _guard852 = cond_wire121_out;
wire _guard853 = early_reset_static_par0_go_out;
wire _guard854 = _guard852 & _guard853;
wire _guard855 = cond_wire24_out;
wire _guard856 = early_reset_static_par0_go_out;
wire _guard857 = _guard855 & _guard856;
wire _guard858 = cond_wire39_out;
wire _guard859 = early_reset_static_par0_go_out;
wire _guard860 = _guard858 & _guard859;
wire _guard861 = fsm_out == 1'd0;
wire _guard862 = cond_wire175_out;
wire _guard863 = _guard861 & _guard862;
wire _guard864 = fsm_out == 1'd0;
wire _guard865 = _guard863 & _guard864;
wire _guard866 = fsm_out == 1'd0;
wire _guard867 = cond_wire179_out;
wire _guard868 = _guard866 & _guard867;
wire _guard869 = fsm_out == 1'd0;
wire _guard870 = _guard868 & _guard869;
wire _guard871 = _guard865 | _guard870;
wire _guard872 = fsm_out == 1'd0;
wire _guard873 = cond_wire183_out;
wire _guard874 = _guard872 & _guard873;
wire _guard875 = fsm_out == 1'd0;
wire _guard876 = _guard874 & _guard875;
wire _guard877 = _guard871 | _guard876;
wire _guard878 = fsm_out == 1'd0;
wire _guard879 = cond_wire187_out;
wire _guard880 = _guard878 & _guard879;
wire _guard881 = fsm_out == 1'd0;
wire _guard882 = _guard880 & _guard881;
wire _guard883 = _guard877 | _guard882;
wire _guard884 = fsm_out == 1'd0;
wire _guard885 = cond_wire191_out;
wire _guard886 = _guard884 & _guard885;
wire _guard887 = fsm_out == 1'd0;
wire _guard888 = _guard886 & _guard887;
wire _guard889 = _guard883 | _guard888;
wire _guard890 = fsm_out == 1'd0;
wire _guard891 = cond_wire195_out;
wire _guard892 = _guard890 & _guard891;
wire _guard893 = fsm_out == 1'd0;
wire _guard894 = _guard892 & _guard893;
wire _guard895 = _guard889 | _guard894;
wire _guard896 = fsm_out == 1'd0;
wire _guard897 = cond_wire199_out;
wire _guard898 = _guard896 & _guard897;
wire _guard899 = fsm_out == 1'd0;
wire _guard900 = _guard898 & _guard899;
wire _guard901 = _guard895 | _guard900;
wire _guard902 = fsm_out == 1'd0;
wire _guard903 = cond_wire203_out;
wire _guard904 = _guard902 & _guard903;
wire _guard905 = fsm_out == 1'd0;
wire _guard906 = _guard904 & _guard905;
wire _guard907 = _guard901 | _guard906;
wire _guard908 = early_reset_static_par0_go_out;
wire _guard909 = _guard907 & _guard908;
wire _guard910 = cond_wire253_out;
wire _guard911 = early_reset_static_par0_go_out;
wire _guard912 = _guard910 & _guard911;
wire _guard913 = cond_wire261_out;
wire _guard914 = early_reset_static_par0_go_out;
wire _guard915 = _guard913 & _guard914;
wire _guard916 = cond_wire257_out;
wire _guard917 = early_reset_static_par0_go_out;
wire _guard918 = _guard916 & _guard917;
wire _guard919 = cond_wire241_out;
wire _guard920 = early_reset_static_par0_go_out;
wire _guard921 = _guard919 & _guard920;
wire _guard922 = cond_wire268_out;
wire _guard923 = early_reset_static_par0_go_out;
wire _guard924 = _guard922 & _guard923;
wire _guard925 = cond_wire249_out;
wire _guard926 = early_reset_static_par0_go_out;
wire _guard927 = _guard925 & _guard926;
wire _guard928 = cond_wire265_out;
wire _guard929 = early_reset_static_par0_go_out;
wire _guard930 = _guard928 & _guard929;
wire _guard931 = cond_wire245_out;
wire _guard932 = early_reset_static_par0_go_out;
wire _guard933 = _guard931 & _guard932;
wire _guard934 = cond_wire19_out;
wire _guard935 = early_reset_static_par0_go_out;
wire _guard936 = _guard934 & _guard935;
wire _guard937 = cond_wire29_out;
wire _guard938 = early_reset_static_par0_go_out;
wire _guard939 = _guard937 & _guard938;
wire _guard940 = fsm_out == 1'd0;
wire _guard941 = cond_wire241_out;
wire _guard942 = _guard940 & _guard941;
wire _guard943 = fsm_out == 1'd0;
wire _guard944 = _guard942 & _guard943;
wire _guard945 = fsm_out == 1'd0;
wire _guard946 = cond_wire245_out;
wire _guard947 = _guard945 & _guard946;
wire _guard948 = fsm_out == 1'd0;
wire _guard949 = _guard947 & _guard948;
wire _guard950 = _guard944 | _guard949;
wire _guard951 = fsm_out == 1'd0;
wire _guard952 = cond_wire249_out;
wire _guard953 = _guard951 & _guard952;
wire _guard954 = fsm_out == 1'd0;
wire _guard955 = _guard953 & _guard954;
wire _guard956 = _guard950 | _guard955;
wire _guard957 = fsm_out == 1'd0;
wire _guard958 = cond_wire253_out;
wire _guard959 = _guard957 & _guard958;
wire _guard960 = fsm_out == 1'd0;
wire _guard961 = _guard959 & _guard960;
wire _guard962 = _guard956 | _guard961;
wire _guard963 = fsm_out == 1'd0;
wire _guard964 = cond_wire257_out;
wire _guard965 = _guard963 & _guard964;
wire _guard966 = fsm_out == 1'd0;
wire _guard967 = _guard965 & _guard966;
wire _guard968 = _guard962 | _guard967;
wire _guard969 = fsm_out == 1'd0;
wire _guard970 = cond_wire261_out;
wire _guard971 = _guard969 & _guard970;
wire _guard972 = fsm_out == 1'd0;
wire _guard973 = _guard971 & _guard972;
wire _guard974 = _guard968 | _guard973;
wire _guard975 = fsm_out == 1'd0;
wire _guard976 = cond_wire265_out;
wire _guard977 = _guard975 & _guard976;
wire _guard978 = fsm_out == 1'd0;
wire _guard979 = _guard977 & _guard978;
wire _guard980 = _guard974 | _guard979;
wire _guard981 = fsm_out == 1'd0;
wire _guard982 = cond_wire268_out;
wire _guard983 = _guard981 & _guard982;
wire _guard984 = fsm_out == 1'd0;
wire _guard985 = _guard983 & _guard984;
wire _guard986 = _guard980 | _guard985;
wire _guard987 = early_reset_static_par0_go_out;
wire _guard988 = _guard986 & _guard987;
wire _guard989 = cond_wire154_out;
wire _guard990 = early_reset_static_par0_go_out;
wire _guard991 = _guard989 & _guard990;
wire _guard992 = cond_wire162_out;
wire _guard993 = early_reset_static_par0_go_out;
wire _guard994 = _guard992 & _guard993;
wire _guard995 = cond_wire158_out;
wire _guard996 = early_reset_static_par0_go_out;
wire _guard997 = _guard995 & _guard996;
wire _guard998 = cond_wire142_out;
wire _guard999 = early_reset_static_par0_go_out;
wire _guard1000 = _guard998 & _guard999;
wire _guard1001 = cond_wire170_out;
wire _guard1002 = early_reset_static_par0_go_out;
wire _guard1003 = _guard1001 & _guard1002;
wire _guard1004 = cond_wire150_out;
wire _guard1005 = early_reset_static_par0_go_out;
wire _guard1006 = _guard1004 & _guard1005;
wire _guard1007 = cond_wire166_out;
wire _guard1008 = early_reset_static_par0_go_out;
wire _guard1009 = _guard1007 & _guard1008;
wire _guard1010 = cond_wire146_out;
wire _guard1011 = early_reset_static_par0_go_out;
wire _guard1012 = _guard1010 & _guard1011;
wire _guard1013 = cond_wire105_out;
wire _guard1014 = early_reset_static_par0_go_out;
wire _guard1015 = _guard1013 & _guard1014;
wire _guard1016 = cond_wire104_out;
wire _guard1017 = early_reset_static_par0_go_out;
wire _guard1018 = _guard1016 & _guard1017;
wire _guard1019 = cond_wire92_out;
wire _guard1020 = early_reset_static_par0_go_out;
wire _guard1021 = _guard1019 & _guard1020;
wire _guard1022 = cond_wire80_out;
wire _guard1023 = early_reset_static_par0_go_out;
wire _guard1024 = _guard1022 & _guard1023;
wire _guard1025 = cond_wire88_out;
wire _guard1026 = early_reset_static_par0_go_out;
wire _guard1027 = _guard1025 & _guard1026;
wire _guard1028 = cond_wire96_out;
wire _guard1029 = early_reset_static_par0_go_out;
wire _guard1030 = _guard1028 & _guard1029;
wire _guard1031 = cond_wire100_out;
wire _guard1032 = early_reset_static_par0_go_out;
wire _guard1033 = _guard1031 & _guard1032;
wire _guard1034 = cond_wire76_out;
wire _guard1035 = early_reset_static_par0_go_out;
wire _guard1036 = _guard1034 & _guard1035;
wire _guard1037 = cond_wire84_out;
wire _guard1038 = early_reset_static_par0_go_out;
wire _guard1039 = _guard1037 & _guard1038;
wire _guard1040 = cond_wire138_out;
wire _guard1041 = early_reset_static_par0_go_out;
wire _guard1042 = _guard1040 & _guard1041;
wire _guard1043 = cond_wire237_out;
wire _guard1044 = early_reset_static_par0_go_out;
wire _guard1045 = _guard1043 & _guard1044;
wire _guard1046 = cond_wire59_out;
wire _guard1047 = early_reset_static_par0_go_out;
wire _guard1048 = _guard1046 & _guard1047;
wire _guard1049 = cond_wire71_out;
wire _guard1050 = early_reset_static_par0_go_out;
wire _guard1051 = _guard1049 & _guard1050;
wire _guard1052 = cond_wire51_out;
wire _guard1053 = early_reset_static_par0_go_out;
wire _guard1054 = _guard1052 & _guard1053;
wire _guard1055 = cond_wire55_out;
wire _guard1056 = early_reset_static_par0_go_out;
wire _guard1057 = _guard1055 & _guard1056;
wire _guard1058 = cond_wire43_out;
wire _guard1059 = early_reset_static_par0_go_out;
wire _guard1060 = _guard1058 & _guard1059;
wire _guard1061 = cond_wire67_out;
wire _guard1062 = early_reset_static_par0_go_out;
wire _guard1063 = _guard1061 & _guard1062;
wire _guard1064 = cond_wire63_out;
wire _guard1065 = early_reset_static_par0_go_out;
wire _guard1066 = _guard1064 & _guard1065;
wire _guard1067 = cond_wire47_out;
wire _guard1068 = early_reset_static_par0_go_out;
wire _guard1069 = _guard1067 & _guard1068;
wire _guard1070 = fsm_out == 1'd0;
wire _guard1071 = cond_wire43_out;
wire _guard1072 = _guard1070 & _guard1071;
wire _guard1073 = fsm_out == 1'd0;
wire _guard1074 = _guard1072 & _guard1073;
wire _guard1075 = fsm_out == 1'd0;
wire _guard1076 = cond_wire47_out;
wire _guard1077 = _guard1075 & _guard1076;
wire _guard1078 = fsm_out == 1'd0;
wire _guard1079 = _guard1077 & _guard1078;
wire _guard1080 = _guard1074 | _guard1079;
wire _guard1081 = fsm_out == 1'd0;
wire _guard1082 = cond_wire51_out;
wire _guard1083 = _guard1081 & _guard1082;
wire _guard1084 = fsm_out == 1'd0;
wire _guard1085 = _guard1083 & _guard1084;
wire _guard1086 = _guard1080 | _guard1085;
wire _guard1087 = fsm_out == 1'd0;
wire _guard1088 = cond_wire55_out;
wire _guard1089 = _guard1087 & _guard1088;
wire _guard1090 = fsm_out == 1'd0;
wire _guard1091 = _guard1089 & _guard1090;
wire _guard1092 = _guard1086 | _guard1091;
wire _guard1093 = fsm_out == 1'd0;
wire _guard1094 = cond_wire59_out;
wire _guard1095 = _guard1093 & _guard1094;
wire _guard1096 = fsm_out == 1'd0;
wire _guard1097 = _guard1095 & _guard1096;
wire _guard1098 = _guard1092 | _guard1097;
wire _guard1099 = fsm_out == 1'd0;
wire _guard1100 = cond_wire63_out;
wire _guard1101 = _guard1099 & _guard1100;
wire _guard1102 = fsm_out == 1'd0;
wire _guard1103 = _guard1101 & _guard1102;
wire _guard1104 = _guard1098 | _guard1103;
wire _guard1105 = fsm_out == 1'd0;
wire _guard1106 = cond_wire67_out;
wire _guard1107 = _guard1105 & _guard1106;
wire _guard1108 = fsm_out == 1'd0;
wire _guard1109 = _guard1107 & _guard1108;
wire _guard1110 = _guard1104 | _guard1109;
wire _guard1111 = fsm_out == 1'd0;
wire _guard1112 = cond_wire71_out;
wire _guard1113 = _guard1111 & _guard1112;
wire _guard1114 = fsm_out == 1'd0;
wire _guard1115 = _guard1113 & _guard1114;
wire _guard1116 = _guard1110 | _guard1115;
wire _guard1117 = early_reset_static_par0_go_out;
wire _guard1118 = _guard1116 & _guard1117;
wire _guard1119 = fsm_out == 1'd0;
wire _guard1120 = cond_wire142_out;
wire _guard1121 = _guard1119 & _guard1120;
wire _guard1122 = fsm_out == 1'd0;
wire _guard1123 = _guard1121 & _guard1122;
wire _guard1124 = fsm_out == 1'd0;
wire _guard1125 = cond_wire146_out;
wire _guard1126 = _guard1124 & _guard1125;
wire _guard1127 = fsm_out == 1'd0;
wire _guard1128 = _guard1126 & _guard1127;
wire _guard1129 = _guard1123 | _guard1128;
wire _guard1130 = fsm_out == 1'd0;
wire _guard1131 = cond_wire150_out;
wire _guard1132 = _guard1130 & _guard1131;
wire _guard1133 = fsm_out == 1'd0;
wire _guard1134 = _guard1132 & _guard1133;
wire _guard1135 = _guard1129 | _guard1134;
wire _guard1136 = fsm_out == 1'd0;
wire _guard1137 = cond_wire154_out;
wire _guard1138 = _guard1136 & _guard1137;
wire _guard1139 = fsm_out == 1'd0;
wire _guard1140 = _guard1138 & _guard1139;
wire _guard1141 = _guard1135 | _guard1140;
wire _guard1142 = fsm_out == 1'd0;
wire _guard1143 = cond_wire158_out;
wire _guard1144 = _guard1142 & _guard1143;
wire _guard1145 = fsm_out == 1'd0;
wire _guard1146 = _guard1144 & _guard1145;
wire _guard1147 = _guard1141 | _guard1146;
wire _guard1148 = fsm_out == 1'd0;
wire _guard1149 = cond_wire162_out;
wire _guard1150 = _guard1148 & _guard1149;
wire _guard1151 = fsm_out == 1'd0;
wire _guard1152 = _guard1150 & _guard1151;
wire _guard1153 = _guard1147 | _guard1152;
wire _guard1154 = fsm_out == 1'd0;
wire _guard1155 = cond_wire166_out;
wire _guard1156 = _guard1154 & _guard1155;
wire _guard1157 = fsm_out == 1'd0;
wire _guard1158 = _guard1156 & _guard1157;
wire _guard1159 = _guard1153 | _guard1158;
wire _guard1160 = fsm_out == 1'd0;
wire _guard1161 = cond_wire170_out;
wire _guard1162 = _guard1160 & _guard1161;
wire _guard1163 = fsm_out == 1'd0;
wire _guard1164 = _guard1162 & _guard1163;
wire _guard1165 = _guard1159 | _guard1164;
wire _guard1166 = early_reset_static_par0_go_out;
wire _guard1167 = _guard1165 & _guard1166;
wire _guard1168 = cond_wire_out;
wire _guard1169 = early_reset_static_par0_go_out;
wire _guard1170 = _guard1168 & _guard1169;
wire _guard1171 = cond_wire4_out;
wire _guard1172 = early_reset_static_par0_go_out;
wire _guard1173 = _guard1171 & _guard1172;
wire _guard1174 = fsm_out == 1'd0;
wire _guard1175 = cond_wire3_out;
wire _guard1176 = _guard1174 & _guard1175;
wire _guard1177 = fsm_out == 1'd0;
wire _guard1178 = _guard1176 & _guard1177;
wire _guard1179 = fsm_out == 1'd0;
wire _guard1180 = cond_wire8_out;
wire _guard1181 = _guard1179 & _guard1180;
wire _guard1182 = fsm_out == 1'd0;
wire _guard1183 = _guard1181 & _guard1182;
wire _guard1184 = _guard1178 | _guard1183;
wire _guard1185 = fsm_out == 1'd0;
wire _guard1186 = cond_wire13_out;
wire _guard1187 = _guard1185 & _guard1186;
wire _guard1188 = fsm_out == 1'd0;
wire _guard1189 = _guard1187 & _guard1188;
wire _guard1190 = _guard1184 | _guard1189;
wire _guard1191 = fsm_out == 1'd0;
wire _guard1192 = cond_wire18_out;
wire _guard1193 = _guard1191 & _guard1192;
wire _guard1194 = fsm_out == 1'd0;
wire _guard1195 = _guard1193 & _guard1194;
wire _guard1196 = _guard1190 | _guard1195;
wire _guard1197 = fsm_out == 1'd0;
wire _guard1198 = cond_wire23_out;
wire _guard1199 = _guard1197 & _guard1198;
wire _guard1200 = fsm_out == 1'd0;
wire _guard1201 = _guard1199 & _guard1200;
wire _guard1202 = _guard1196 | _guard1201;
wire _guard1203 = fsm_out == 1'd0;
wire _guard1204 = cond_wire28_out;
wire _guard1205 = _guard1203 & _guard1204;
wire _guard1206 = fsm_out == 1'd0;
wire _guard1207 = _guard1205 & _guard1206;
wire _guard1208 = _guard1202 | _guard1207;
wire _guard1209 = fsm_out == 1'd0;
wire _guard1210 = cond_wire33_out;
wire _guard1211 = _guard1209 & _guard1210;
wire _guard1212 = fsm_out == 1'd0;
wire _guard1213 = _guard1211 & _guard1212;
wire _guard1214 = _guard1208 | _guard1213;
wire _guard1215 = fsm_out == 1'd0;
wire _guard1216 = cond_wire38_out;
wire _guard1217 = _guard1215 & _guard1216;
wire _guard1218 = fsm_out == 1'd0;
wire _guard1219 = _guard1217 & _guard1218;
wire _guard1220 = _guard1214 | _guard1219;
wire _guard1221 = early_reset_static_par0_go_out;
wire _guard1222 = _guard1220 & _guard1221;
wire _guard1223 = fsm_out == 1'd0;
wire _guard1224 = cond_wire76_out;
wire _guard1225 = _guard1223 & _guard1224;
wire _guard1226 = fsm_out == 1'd0;
wire _guard1227 = _guard1225 & _guard1226;
wire _guard1228 = fsm_out == 1'd0;
wire _guard1229 = cond_wire80_out;
wire _guard1230 = _guard1228 & _guard1229;
wire _guard1231 = fsm_out == 1'd0;
wire _guard1232 = _guard1230 & _guard1231;
wire _guard1233 = _guard1227 | _guard1232;
wire _guard1234 = fsm_out == 1'd0;
wire _guard1235 = cond_wire84_out;
wire _guard1236 = _guard1234 & _guard1235;
wire _guard1237 = fsm_out == 1'd0;
wire _guard1238 = _guard1236 & _guard1237;
wire _guard1239 = _guard1233 | _guard1238;
wire _guard1240 = fsm_out == 1'd0;
wire _guard1241 = cond_wire88_out;
wire _guard1242 = _guard1240 & _guard1241;
wire _guard1243 = fsm_out == 1'd0;
wire _guard1244 = _guard1242 & _guard1243;
wire _guard1245 = _guard1239 | _guard1244;
wire _guard1246 = fsm_out == 1'd0;
wire _guard1247 = cond_wire92_out;
wire _guard1248 = _guard1246 & _guard1247;
wire _guard1249 = fsm_out == 1'd0;
wire _guard1250 = _guard1248 & _guard1249;
wire _guard1251 = _guard1245 | _guard1250;
wire _guard1252 = fsm_out == 1'd0;
wire _guard1253 = cond_wire96_out;
wire _guard1254 = _guard1252 & _guard1253;
wire _guard1255 = fsm_out == 1'd0;
wire _guard1256 = _guard1254 & _guard1255;
wire _guard1257 = _guard1251 | _guard1256;
wire _guard1258 = fsm_out == 1'd0;
wire _guard1259 = cond_wire100_out;
wire _guard1260 = _guard1258 & _guard1259;
wire _guard1261 = fsm_out == 1'd0;
wire _guard1262 = _guard1260 & _guard1261;
wire _guard1263 = _guard1257 | _guard1262;
wire _guard1264 = fsm_out == 1'd0;
wire _guard1265 = cond_wire104_out;
wire _guard1266 = _guard1264 & _guard1265;
wire _guard1267 = fsm_out == 1'd0;
wire _guard1268 = _guard1266 & _guard1267;
wire _guard1269 = _guard1263 | _guard1268;
wire _guard1270 = early_reset_static_par0_go_out;
wire _guard1271 = _guard1269 & _guard1270;
wire _guard1272 = fsm_out == 1'd0;
wire _guard1273 = cond_wire109_out;
wire _guard1274 = _guard1272 & _guard1273;
wire _guard1275 = fsm_out == 1'd0;
wire _guard1276 = _guard1274 & _guard1275;
wire _guard1277 = fsm_out == 1'd0;
wire _guard1278 = cond_wire113_out;
wire _guard1279 = _guard1277 & _guard1278;
wire _guard1280 = fsm_out == 1'd0;
wire _guard1281 = _guard1279 & _guard1280;
wire _guard1282 = _guard1276 | _guard1281;
wire _guard1283 = fsm_out == 1'd0;
wire _guard1284 = cond_wire117_out;
wire _guard1285 = _guard1283 & _guard1284;
wire _guard1286 = fsm_out == 1'd0;
wire _guard1287 = _guard1285 & _guard1286;
wire _guard1288 = _guard1282 | _guard1287;
wire _guard1289 = fsm_out == 1'd0;
wire _guard1290 = cond_wire121_out;
wire _guard1291 = _guard1289 & _guard1290;
wire _guard1292 = fsm_out == 1'd0;
wire _guard1293 = _guard1291 & _guard1292;
wire _guard1294 = _guard1288 | _guard1293;
wire _guard1295 = fsm_out == 1'd0;
wire _guard1296 = cond_wire125_out;
wire _guard1297 = _guard1295 & _guard1296;
wire _guard1298 = fsm_out == 1'd0;
wire _guard1299 = _guard1297 & _guard1298;
wire _guard1300 = _guard1294 | _guard1299;
wire _guard1301 = fsm_out == 1'd0;
wire _guard1302 = cond_wire129_out;
wire _guard1303 = _guard1301 & _guard1302;
wire _guard1304 = fsm_out == 1'd0;
wire _guard1305 = _guard1303 & _guard1304;
wire _guard1306 = _guard1300 | _guard1305;
wire _guard1307 = fsm_out == 1'd0;
wire _guard1308 = cond_wire133_out;
wire _guard1309 = _guard1307 & _guard1308;
wire _guard1310 = fsm_out == 1'd0;
wire _guard1311 = _guard1309 & _guard1310;
wire _guard1312 = _guard1306 | _guard1311;
wire _guard1313 = fsm_out == 1'd0;
wire _guard1314 = cond_wire137_out;
wire _guard1315 = _guard1313 & _guard1314;
wire _guard1316 = fsm_out == 1'd0;
wire _guard1317 = _guard1315 & _guard1316;
wire _guard1318 = _guard1312 | _guard1317;
wire _guard1319 = early_reset_static_par0_go_out;
wire _guard1320 = _guard1318 & _guard1319;
wire _guard1321 = cond_wire224_out;
wire _guard1322 = early_reset_static_par0_go_out;
wire _guard1323 = _guard1321 & _guard1322;
wire _guard1324 = cond_wire208_out;
wire _guard1325 = early_reset_static_par0_go_out;
wire _guard1326 = _guard1324 & _guard1325;
wire _guard1327 = cond_wire212_out;
wire _guard1328 = early_reset_static_par0_go_out;
wire _guard1329 = _guard1327 & _guard1328;
wire _guard1330 = cond_wire228_out;
wire _guard1331 = early_reset_static_par0_go_out;
wire _guard1332 = _guard1330 & _guard1331;
wire _guard1333 = cond_wire216_out;
wire _guard1334 = early_reset_static_par0_go_out;
wire _guard1335 = _guard1333 & _guard1334;
wire _guard1336 = cond_wire220_out;
wire _guard1337 = early_reset_static_par0_go_out;
wire _guard1338 = _guard1336 & _guard1337;
wire _guard1339 = cond_wire236_out;
wire _guard1340 = early_reset_static_par0_go_out;
wire _guard1341 = _guard1339 & _guard1340;
wire _guard1342 = cond_wire232_out;
wire _guard1343 = early_reset_static_par0_go_out;
wire _guard1344 = _guard1342 & _guard1343;
wire _guard1345 = fsm_out == 1'd0;
wire _guard1346 = cond_wire208_out;
wire _guard1347 = _guard1345 & _guard1346;
wire _guard1348 = fsm_out == 1'd0;
wire _guard1349 = _guard1347 & _guard1348;
wire _guard1350 = fsm_out == 1'd0;
wire _guard1351 = cond_wire212_out;
wire _guard1352 = _guard1350 & _guard1351;
wire _guard1353 = fsm_out == 1'd0;
wire _guard1354 = _guard1352 & _guard1353;
wire _guard1355 = _guard1349 | _guard1354;
wire _guard1356 = fsm_out == 1'd0;
wire _guard1357 = cond_wire216_out;
wire _guard1358 = _guard1356 & _guard1357;
wire _guard1359 = fsm_out == 1'd0;
wire _guard1360 = _guard1358 & _guard1359;
wire _guard1361 = _guard1355 | _guard1360;
wire _guard1362 = fsm_out == 1'd0;
wire _guard1363 = cond_wire220_out;
wire _guard1364 = _guard1362 & _guard1363;
wire _guard1365 = fsm_out == 1'd0;
wire _guard1366 = _guard1364 & _guard1365;
wire _guard1367 = _guard1361 | _guard1366;
wire _guard1368 = fsm_out == 1'd0;
wire _guard1369 = cond_wire224_out;
wire _guard1370 = _guard1368 & _guard1369;
wire _guard1371 = fsm_out == 1'd0;
wire _guard1372 = _guard1370 & _guard1371;
wire _guard1373 = _guard1367 | _guard1372;
wire _guard1374 = fsm_out == 1'd0;
wire _guard1375 = cond_wire228_out;
wire _guard1376 = _guard1374 & _guard1375;
wire _guard1377 = fsm_out == 1'd0;
wire _guard1378 = _guard1376 & _guard1377;
wire _guard1379 = _guard1373 | _guard1378;
wire _guard1380 = fsm_out == 1'd0;
wire _guard1381 = cond_wire232_out;
wire _guard1382 = _guard1380 & _guard1381;
wire _guard1383 = fsm_out == 1'd0;
wire _guard1384 = _guard1382 & _guard1383;
wire _guard1385 = _guard1379 | _guard1384;
wire _guard1386 = fsm_out == 1'd0;
wire _guard1387 = cond_wire236_out;
wire _guard1388 = _guard1386 & _guard1387;
wire _guard1389 = fsm_out == 1'd0;
wire _guard1390 = _guard1388 & _guard1389;
wire _guard1391 = _guard1385 | _guard1390;
wire _guard1392 = early_reset_static_par0_go_out;
wire _guard1393 = _guard1391 & _guard1392;
wire _guard1394 = cond_wire253_out;
wire _guard1395 = early_reset_static_par0_go_out;
wire _guard1396 = _guard1394 & _guard1395;
wire _guard1397 = cond_wire257_out;
wire _guard1398 = early_reset_static_par0_go_out;
wire _guard1399 = _guard1397 & _guard1398;
wire _guard1400 = cond_wire241_out;
wire _guard1401 = early_reset_static_par0_go_out;
wire _guard1402 = _guard1400 & _guard1401;
wire _guard1403 = cond_wire261_out;
wire _guard1404 = early_reset_static_par0_go_out;
wire _guard1405 = _guard1403 & _guard1404;
wire _guard1406 = cond_wire265_out;
wire _guard1407 = early_reset_static_par0_go_out;
wire _guard1408 = _guard1406 & _guard1407;
wire _guard1409 = cond_wire245_out;
wire _guard1410 = early_reset_static_par0_go_out;
wire _guard1411 = _guard1409 & _guard1410;
wire _guard1412 = cond_wire249_out;
wire _guard1413 = early_reset_static_par0_go_out;
wire _guard1414 = _guard1412 & _guard1413;
wire _guard1415 = cond_wire268_out;
wire _guard1416 = early_reset_static_par0_go_out;
wire _guard1417 = _guard1415 & _guard1416;
wire _guard1418 = cond_wire72_out;
wire _guard1419 = early_reset_static_par0_go_out;
wire _guard1420 = _guard1418 & _guard1419;
wire _guard1421 = cond_wire18_out;
wire _guard1422 = early_reset_static_par0_go_out;
wire _guard1423 = _guard1421 & _guard1422;
wire _guard1424 = cond_wire28_out;
wire _guard1425 = early_reset_static_par0_go_out;
wire _guard1426 = _guard1424 & _guard1425;
wire _guard1427 = cond_wire23_out;
wire _guard1428 = early_reset_static_par0_go_out;
wire _guard1429 = _guard1427 & _guard1428;
wire _guard1430 = cond_wire3_out;
wire _guard1431 = early_reset_static_par0_go_out;
wire _guard1432 = _guard1430 & _guard1431;
wire _guard1433 = cond_wire38_out;
wire _guard1434 = early_reset_static_par0_go_out;
wire _guard1435 = _guard1433 & _guard1434;
wire _guard1436 = cond_wire13_out;
wire _guard1437 = early_reset_static_par0_go_out;
wire _guard1438 = _guard1436 & _guard1437;
wire _guard1439 = cond_wire33_out;
wire _guard1440 = early_reset_static_par0_go_out;
wire _guard1441 = _guard1439 & _guard1440;
wire _guard1442 = cond_wire8_out;
wire _guard1443 = early_reset_static_par0_go_out;
wire _guard1444 = _guard1442 & _guard1443;
wire _guard1445 = cond_wire121_out;
wire _guard1446 = early_reset_static_par0_go_out;
wire _guard1447 = _guard1445 & _guard1446;
wire _guard1448 = cond_wire129_out;
wire _guard1449 = early_reset_static_par0_go_out;
wire _guard1450 = _guard1448 & _guard1449;
wire _guard1451 = cond_wire125_out;
wire _guard1452 = early_reset_static_par0_go_out;
wire _guard1453 = _guard1451 & _guard1452;
wire _guard1454 = cond_wire109_out;
wire _guard1455 = early_reset_static_par0_go_out;
wire _guard1456 = _guard1454 & _guard1455;
wire _guard1457 = cond_wire137_out;
wire _guard1458 = early_reset_static_par0_go_out;
wire _guard1459 = _guard1457 & _guard1458;
wire _guard1460 = cond_wire117_out;
wire _guard1461 = early_reset_static_par0_go_out;
wire _guard1462 = _guard1460 & _guard1461;
wire _guard1463 = cond_wire133_out;
wire _guard1464 = early_reset_static_par0_go_out;
wire _guard1465 = _guard1463 & _guard1464;
wire _guard1466 = cond_wire113_out;
wire _guard1467 = early_reset_static_par0_go_out;
wire _guard1468 = _guard1466 & _guard1467;
wire _guard1469 = cond_wire14_out;
wire _guard1470 = early_reset_static_par0_go_out;
wire _guard1471 = _guard1469 & _guard1470;
wire _guard1472 = cond_wire34_out;
wire _guard1473 = early_reset_static_par0_go_out;
wire _guard1474 = _guard1472 & _guard1473;
wire _guard1475 = cond_wire88_out;
wire _guard1476 = early_reset_static_par0_go_out;
wire _guard1477 = _guard1475 & _guard1476;
wire _guard1478 = cond_wire96_out;
wire _guard1479 = early_reset_static_par0_go_out;
wire _guard1480 = _guard1478 & _guard1479;
wire _guard1481 = cond_wire92_out;
wire _guard1482 = early_reset_static_par0_go_out;
wire _guard1483 = _guard1481 & _guard1482;
wire _guard1484 = cond_wire76_out;
wire _guard1485 = early_reset_static_par0_go_out;
wire _guard1486 = _guard1484 & _guard1485;
wire _guard1487 = cond_wire104_out;
wire _guard1488 = early_reset_static_par0_go_out;
wire _guard1489 = _guard1487 & _guard1488;
wire _guard1490 = cond_wire84_out;
wire _guard1491 = early_reset_static_par0_go_out;
wire _guard1492 = _guard1490 & _guard1491;
wire _guard1493 = cond_wire100_out;
wire _guard1494 = early_reset_static_par0_go_out;
wire _guard1495 = _guard1493 & _guard1494;
wire _guard1496 = cond_wire80_out;
wire _guard1497 = early_reset_static_par0_go_out;
wire _guard1498 = _guard1496 & _guard1497;
wire _guard1499 = early_reset_static_par0_go_out;
wire _guard1500 = ~_guard0;
wire _guard1501 = early_reset_static_par0_go_out;
wire _guard1502 = _guard1500 & _guard1501;
wire _guard1503 = ~_guard0;
wire _guard1504 = early_reset_static_par0_go_out;
wire _guard1505 = _guard1503 & _guard1504;
wire _guard1506 = early_reset_static_par0_go_out;
wire _guard1507 = early_reset_static_par0_go_out;
wire _guard1508 = early_reset_static_par0_go_out;
wire _guard1509 = early_reset_static_par0_go_out;
wire _guard1510 = ~_guard0;
wire _guard1511 = early_reset_static_par0_go_out;
wire _guard1512 = _guard1510 & _guard1511;
wire _guard1513 = early_reset_static_par0_go_out;
wire _guard1514 = ~_guard0;
wire _guard1515 = early_reset_static_par0_go_out;
wire _guard1516 = _guard1514 & _guard1515;
wire _guard1517 = early_reset_static_par0_go_out;
wire _guard1518 = early_reset_static_par0_go_out;
wire _guard1519 = early_reset_static_par0_go_out;
wire _guard1520 = ~_guard0;
wire _guard1521 = early_reset_static_par0_go_out;
wire _guard1522 = _guard1520 & _guard1521;
wire _guard1523 = ~_guard0;
wire _guard1524 = early_reset_static_par0_go_out;
wire _guard1525 = _guard1523 & _guard1524;
wire _guard1526 = early_reset_static_par0_go_out;
wire _guard1527 = early_reset_static_par0_go_out;
wire _guard1528 = early_reset_static_par0_go_out;
wire _guard1529 = early_reset_static_par0_go_out;
wire _guard1530 = early_reset_static_par0_go_out;
wire _guard1531 = early_reset_static_par0_go_out;
wire _guard1532 = ~_guard0;
wire _guard1533 = early_reset_static_par0_go_out;
wire _guard1534 = _guard1532 & _guard1533;
wire _guard1535 = early_reset_static_par0_go_out;
wire _guard1536 = early_reset_static_par0_go_out;
wire _guard1537 = early_reset_static_par0_go_out;
wire _guard1538 = early_reset_static_par0_go_out;
wire _guard1539 = early_reset_static_par0_go_out;
wire _guard1540 = early_reset_static_par0_go_out;
wire _guard1541 = ~_guard0;
wire _guard1542 = early_reset_static_par0_go_out;
wire _guard1543 = _guard1541 & _guard1542;
wire _guard1544 = early_reset_static_par0_go_out;
wire _guard1545 = early_reset_static_par0_go_out;
wire _guard1546 = early_reset_static_par0_go_out;
wire _guard1547 = ~_guard0;
wire _guard1548 = early_reset_static_par0_go_out;
wire _guard1549 = _guard1547 & _guard1548;
wire _guard1550 = early_reset_static_par0_go_out;
wire _guard1551 = early_reset_static_par0_go_out;
wire _guard1552 = early_reset_static_par0_go_out;
wire _guard1553 = ~_guard0;
wire _guard1554 = early_reset_static_par0_go_out;
wire _guard1555 = _guard1553 & _guard1554;
wire _guard1556 = early_reset_static_par0_go_out;
wire _guard1557 = ~_guard0;
wire _guard1558 = early_reset_static_par0_go_out;
wire _guard1559 = _guard1557 & _guard1558;
wire _guard1560 = early_reset_static_par0_go_out;
wire _guard1561 = early_reset_static_par0_go_out;
wire _guard1562 = ~_guard0;
wire _guard1563 = early_reset_static_par0_go_out;
wire _guard1564 = _guard1562 & _guard1563;
wire _guard1565 = early_reset_static_par0_go_out;
wire _guard1566 = early_reset_static_par0_go_out;
wire _guard1567 = early_reset_static_par0_go_out;
wire _guard1568 = early_reset_static_par0_go_out;
wire _guard1569 = early_reset_static_par0_go_out;
wire _guard1570 = ~_guard0;
wire _guard1571 = early_reset_static_par0_go_out;
wire _guard1572 = _guard1570 & _guard1571;
wire _guard1573 = early_reset_static_par0_go_out;
wire _guard1574 = early_reset_static_par0_go_out;
wire _guard1575 = early_reset_static_par0_go_out;
wire _guard1576 = early_reset_static_par0_go_out;
wire _guard1577 = early_reset_static_par0_go_out;
wire _guard1578 = early_reset_static_par0_go_out;
wire _guard1579 = early_reset_static_par0_go_out;
wire _guard1580 = ~_guard0;
wire _guard1581 = early_reset_static_par0_go_out;
wire _guard1582 = _guard1580 & _guard1581;
wire _guard1583 = early_reset_static_par0_go_out;
wire _guard1584 = early_reset_static_par0_go_out;
wire _guard1585 = ~_guard0;
wire _guard1586 = early_reset_static_par0_go_out;
wire _guard1587 = _guard1585 & _guard1586;
wire _guard1588 = early_reset_static_par0_go_out;
wire _guard1589 = early_reset_static_par0_go_out;
wire _guard1590 = early_reset_static_par0_go_out;
wire _guard1591 = ~_guard0;
wire _guard1592 = early_reset_static_par0_go_out;
wire _guard1593 = _guard1591 & _guard1592;
wire _guard1594 = early_reset_static_par0_go_out;
wire _guard1595 = early_reset_static_par0_go_out;
wire _guard1596 = early_reset_static_par0_go_out;
wire _guard1597 = early_reset_static_par0_go_out;
wire _guard1598 = early_reset_static_par0_go_out;
wire _guard1599 = early_reset_static_par0_go_out;
wire _guard1600 = ~_guard0;
wire _guard1601 = early_reset_static_par0_go_out;
wire _guard1602 = _guard1600 & _guard1601;
wire _guard1603 = early_reset_static_par0_go_out;
wire _guard1604 = fsm_out == 1'd0;
wire _guard1605 = early_reset_static_par0_go_out;
wire _guard1606 = _guard1604 & _guard1605;
wire _guard1607 = fsm_out != 1'd0;
wire _guard1608 = early_reset_static_par0_go_out;
wire _guard1609 = _guard1607 & _guard1608;
wire _guard1610 = early_reset_static_seq_go_out;
wire _guard1611 = early_reset_static_seq_go_out;
wire _guard1612 = fsm0_out >= 5'd1;
wire _guard1613 = fsm0_out < 5'd29;
wire _guard1614 = _guard1612 & _guard1613;
wire _guard1615 = early_reset_static_seq_go_out;
wire _guard1616 = _guard1614 & _guard1615;
wire _guard1617 = cond_wire29_out;
wire _guard1618 = early_reset_static_par0_go_out;
wire _guard1619 = _guard1617 & _guard1618;
wire _guard1620 = cond_wire29_out;
wire _guard1621 = early_reset_static_par0_go_out;
wire _guard1622 = _guard1620 & _guard1621;
wire _guard1623 = cond_wire53_out;
wire _guard1624 = early_reset_static_par0_go_out;
wire _guard1625 = _guard1623 & _guard1624;
wire _guard1626 = cond_wire53_out;
wire _guard1627 = early_reset_static_par0_go_out;
wire _guard1628 = _guard1626 & _guard1627;
wire _guard1629 = cond_wire26_out;
wire _guard1630 = early_reset_static_par0_go_out;
wire _guard1631 = _guard1629 & _guard1630;
wire _guard1632 = cond_wire26_out;
wire _guard1633 = early_reset_static_par0_go_out;
wire _guard1634 = _guard1632 & _guard1633;
wire _guard1635 = cond_wire57_out;
wire _guard1636 = early_reset_static_par0_go_out;
wire _guard1637 = _guard1635 & _guard1636;
wire _guard1638 = cond_wire57_out;
wire _guard1639 = early_reset_static_par0_go_out;
wire _guard1640 = _guard1638 & _guard1639;
wire _guard1641 = cond_wire124_out;
wire _guard1642 = early_reset_static_par0_go_out;
wire _guard1643 = _guard1641 & _guard1642;
wire _guard1644 = cond_wire122_out;
wire _guard1645 = early_reset_static_par0_go_out;
wire _guard1646 = _guard1644 & _guard1645;
wire _guard1647 = fsm_out == 1'd0;
wire _guard1648 = cond_wire122_out;
wire _guard1649 = _guard1647 & _guard1648;
wire _guard1650 = fsm_out == 1'd0;
wire _guard1651 = _guard1649 & _guard1650;
wire _guard1652 = fsm_out == 1'd0;
wire _guard1653 = cond_wire124_out;
wire _guard1654 = _guard1652 & _guard1653;
wire _guard1655 = fsm_out == 1'd0;
wire _guard1656 = _guard1654 & _guard1655;
wire _guard1657 = _guard1651 | _guard1656;
wire _guard1658 = early_reset_static_par0_go_out;
wire _guard1659 = _guard1657 & _guard1658;
wire _guard1660 = fsm_out == 1'd0;
wire _guard1661 = cond_wire122_out;
wire _guard1662 = _guard1660 & _guard1661;
wire _guard1663 = fsm_out == 1'd0;
wire _guard1664 = _guard1662 & _guard1663;
wire _guard1665 = fsm_out == 1'd0;
wire _guard1666 = cond_wire124_out;
wire _guard1667 = _guard1665 & _guard1666;
wire _guard1668 = fsm_out == 1'd0;
wire _guard1669 = _guard1667 & _guard1668;
wire _guard1670 = _guard1664 | _guard1669;
wire _guard1671 = early_reset_static_par0_go_out;
wire _guard1672 = _guard1670 & _guard1671;
wire _guard1673 = fsm_out == 1'd0;
wire _guard1674 = cond_wire122_out;
wire _guard1675 = _guard1673 & _guard1674;
wire _guard1676 = fsm_out == 1'd0;
wire _guard1677 = _guard1675 & _guard1676;
wire _guard1678 = fsm_out == 1'd0;
wire _guard1679 = cond_wire124_out;
wire _guard1680 = _guard1678 & _guard1679;
wire _guard1681 = fsm_out == 1'd0;
wire _guard1682 = _guard1680 & _guard1681;
wire _guard1683 = _guard1677 | _guard1682;
wire _guard1684 = early_reset_static_par0_go_out;
wire _guard1685 = _guard1683 & _guard1684;
wire _guard1686 = cond_wire136_out;
wire _guard1687 = early_reset_static_par0_go_out;
wire _guard1688 = _guard1686 & _guard1687;
wire _guard1689 = cond_wire134_out;
wire _guard1690 = early_reset_static_par0_go_out;
wire _guard1691 = _guard1689 & _guard1690;
wire _guard1692 = fsm_out == 1'd0;
wire _guard1693 = cond_wire134_out;
wire _guard1694 = _guard1692 & _guard1693;
wire _guard1695 = fsm_out == 1'd0;
wire _guard1696 = _guard1694 & _guard1695;
wire _guard1697 = fsm_out == 1'd0;
wire _guard1698 = cond_wire136_out;
wire _guard1699 = _guard1697 & _guard1698;
wire _guard1700 = fsm_out == 1'd0;
wire _guard1701 = _guard1699 & _guard1700;
wire _guard1702 = _guard1696 | _guard1701;
wire _guard1703 = early_reset_static_par0_go_out;
wire _guard1704 = _guard1702 & _guard1703;
wire _guard1705 = fsm_out == 1'd0;
wire _guard1706 = cond_wire134_out;
wire _guard1707 = _guard1705 & _guard1706;
wire _guard1708 = fsm_out == 1'd0;
wire _guard1709 = _guard1707 & _guard1708;
wire _guard1710 = fsm_out == 1'd0;
wire _guard1711 = cond_wire136_out;
wire _guard1712 = _guard1710 & _guard1711;
wire _guard1713 = fsm_out == 1'd0;
wire _guard1714 = _guard1712 & _guard1713;
wire _guard1715 = _guard1709 | _guard1714;
wire _guard1716 = early_reset_static_par0_go_out;
wire _guard1717 = _guard1715 & _guard1716;
wire _guard1718 = fsm_out == 1'd0;
wire _guard1719 = cond_wire134_out;
wire _guard1720 = _guard1718 & _guard1719;
wire _guard1721 = fsm_out == 1'd0;
wire _guard1722 = _guard1720 & _guard1721;
wire _guard1723 = fsm_out == 1'd0;
wire _guard1724 = cond_wire136_out;
wire _guard1725 = _guard1723 & _guard1724;
wire _guard1726 = fsm_out == 1'd0;
wire _guard1727 = _guard1725 & _guard1726;
wire _guard1728 = _guard1722 | _guard1727;
wire _guard1729 = early_reset_static_par0_go_out;
wire _guard1730 = _guard1728 & _guard1729;
wire _guard1731 = cond_wire141_out;
wire _guard1732 = early_reset_static_par0_go_out;
wire _guard1733 = _guard1731 & _guard1732;
wire _guard1734 = cond_wire139_out;
wire _guard1735 = early_reset_static_par0_go_out;
wire _guard1736 = _guard1734 & _guard1735;
wire _guard1737 = fsm_out == 1'd0;
wire _guard1738 = cond_wire139_out;
wire _guard1739 = _guard1737 & _guard1738;
wire _guard1740 = fsm_out == 1'd0;
wire _guard1741 = _guard1739 & _guard1740;
wire _guard1742 = fsm_out == 1'd0;
wire _guard1743 = cond_wire141_out;
wire _guard1744 = _guard1742 & _guard1743;
wire _guard1745 = fsm_out == 1'd0;
wire _guard1746 = _guard1744 & _guard1745;
wire _guard1747 = _guard1741 | _guard1746;
wire _guard1748 = early_reset_static_par0_go_out;
wire _guard1749 = _guard1747 & _guard1748;
wire _guard1750 = fsm_out == 1'd0;
wire _guard1751 = cond_wire139_out;
wire _guard1752 = _guard1750 & _guard1751;
wire _guard1753 = fsm_out == 1'd0;
wire _guard1754 = _guard1752 & _guard1753;
wire _guard1755 = fsm_out == 1'd0;
wire _guard1756 = cond_wire141_out;
wire _guard1757 = _guard1755 & _guard1756;
wire _guard1758 = fsm_out == 1'd0;
wire _guard1759 = _guard1757 & _guard1758;
wire _guard1760 = _guard1754 | _guard1759;
wire _guard1761 = early_reset_static_par0_go_out;
wire _guard1762 = _guard1760 & _guard1761;
wire _guard1763 = fsm_out == 1'd0;
wire _guard1764 = cond_wire139_out;
wire _guard1765 = _guard1763 & _guard1764;
wire _guard1766 = fsm_out == 1'd0;
wire _guard1767 = _guard1765 & _guard1766;
wire _guard1768 = fsm_out == 1'd0;
wire _guard1769 = cond_wire141_out;
wire _guard1770 = _guard1768 & _guard1769;
wire _guard1771 = fsm_out == 1'd0;
wire _guard1772 = _guard1770 & _guard1771;
wire _guard1773 = _guard1767 | _guard1772;
wire _guard1774 = early_reset_static_par0_go_out;
wire _guard1775 = _guard1773 & _guard1774;
wire _guard1776 = cond_wire144_out;
wire _guard1777 = early_reset_static_par0_go_out;
wire _guard1778 = _guard1776 & _guard1777;
wire _guard1779 = cond_wire144_out;
wire _guard1780 = early_reset_static_par0_go_out;
wire _guard1781 = _guard1779 & _guard1780;
wire _guard1782 = cond_wire174_out;
wire _guard1783 = early_reset_static_par0_go_out;
wire _guard1784 = _guard1782 & _guard1783;
wire _guard1785 = cond_wire172_out;
wire _guard1786 = early_reset_static_par0_go_out;
wire _guard1787 = _guard1785 & _guard1786;
wire _guard1788 = fsm_out == 1'd0;
wire _guard1789 = cond_wire172_out;
wire _guard1790 = _guard1788 & _guard1789;
wire _guard1791 = fsm_out == 1'd0;
wire _guard1792 = _guard1790 & _guard1791;
wire _guard1793 = fsm_out == 1'd0;
wire _guard1794 = cond_wire174_out;
wire _guard1795 = _guard1793 & _guard1794;
wire _guard1796 = fsm_out == 1'd0;
wire _guard1797 = _guard1795 & _guard1796;
wire _guard1798 = _guard1792 | _guard1797;
wire _guard1799 = early_reset_static_par0_go_out;
wire _guard1800 = _guard1798 & _guard1799;
wire _guard1801 = fsm_out == 1'd0;
wire _guard1802 = cond_wire172_out;
wire _guard1803 = _guard1801 & _guard1802;
wire _guard1804 = fsm_out == 1'd0;
wire _guard1805 = _guard1803 & _guard1804;
wire _guard1806 = fsm_out == 1'd0;
wire _guard1807 = cond_wire174_out;
wire _guard1808 = _guard1806 & _guard1807;
wire _guard1809 = fsm_out == 1'd0;
wire _guard1810 = _guard1808 & _guard1809;
wire _guard1811 = _guard1805 | _guard1810;
wire _guard1812 = early_reset_static_par0_go_out;
wire _guard1813 = _guard1811 & _guard1812;
wire _guard1814 = fsm_out == 1'd0;
wire _guard1815 = cond_wire172_out;
wire _guard1816 = _guard1814 & _guard1815;
wire _guard1817 = fsm_out == 1'd0;
wire _guard1818 = _guard1816 & _guard1817;
wire _guard1819 = fsm_out == 1'd0;
wire _guard1820 = cond_wire174_out;
wire _guard1821 = _guard1819 & _guard1820;
wire _guard1822 = fsm_out == 1'd0;
wire _guard1823 = _guard1821 & _guard1822;
wire _guard1824 = _guard1818 | _guard1823;
wire _guard1825 = early_reset_static_par0_go_out;
wire _guard1826 = _guard1824 & _guard1825;
wire _guard1827 = cond_wire193_out;
wire _guard1828 = early_reset_static_par0_go_out;
wire _guard1829 = _guard1827 & _guard1828;
wire _guard1830 = cond_wire193_out;
wire _guard1831 = early_reset_static_par0_go_out;
wire _guard1832 = _guard1830 & _guard1831;
wire _guard1833 = cond_wire222_out;
wire _guard1834 = early_reset_static_par0_go_out;
wire _guard1835 = _guard1833 & _guard1834;
wire _guard1836 = cond_wire222_out;
wire _guard1837 = early_reset_static_par0_go_out;
wire _guard1838 = _guard1836 & _guard1837;
wire _guard1839 = cond_wire197_out;
wire _guard1840 = early_reset_static_par0_go_out;
wire _guard1841 = _guard1839 & _guard1840;
wire _guard1842 = cond_wire197_out;
wire _guard1843 = early_reset_static_par0_go_out;
wire _guard1844 = _guard1842 & _guard1843;
wire _guard1845 = fsm0_out == 5'd0;
wire _guard1846 = early_reset_static_seq_go_out;
wire _guard1847 = _guard1845 & _guard1846;
wire _guard1848 = cond_wire_out;
wire _guard1849 = early_reset_static_par0_go_out;
wire _guard1850 = _guard1848 & _guard1849;
wire _guard1851 = _guard1847 | _guard1850;
wire _guard1852 = fsm0_out == 5'd0;
wire _guard1853 = early_reset_static_seq_go_out;
wire _guard1854 = _guard1852 & _guard1853;
wire _guard1855 = cond_wire_out;
wire _guard1856 = early_reset_static_par0_go_out;
wire _guard1857 = _guard1855 & _guard1856;
wire _guard1858 = fsm0_out == 5'd0;
wire _guard1859 = early_reset_static_seq_go_out;
wire _guard1860 = _guard1858 & _guard1859;
wire _guard1861 = early_reset_static_par0_go_out;
wire _guard1862 = _guard1860 | _guard1861;
wire _guard1863 = fsm0_out == 5'd0;
wire _guard1864 = early_reset_static_seq_go_out;
wire _guard1865 = _guard1863 & _guard1864;
wire _guard1866 = early_reset_static_par0_go_out;
wire _guard1867 = early_reset_static_par0_go_out;
wire _guard1868 = early_reset_static_par0_go_out;
wire _guard1869 = fsm0_out == 5'd0;
wire _guard1870 = early_reset_static_seq_go_out;
wire _guard1871 = _guard1869 & _guard1870;
wire _guard1872 = early_reset_static_par0_go_out;
wire _guard1873 = _guard1871 | _guard1872;
wire _guard1874 = early_reset_static_par0_go_out;
wire _guard1875 = fsm0_out == 5'd0;
wire _guard1876 = early_reset_static_seq_go_out;
wire _guard1877 = _guard1875 & _guard1876;
wire _guard1878 = early_reset_static_par0_go_out;
wire _guard1879 = early_reset_static_par0_go_out;
wire _guard1880 = fsm0_out == 5'd0;
wire _guard1881 = early_reset_static_seq_go_out;
wire _guard1882 = _guard1880 & _guard1881;
wire _guard1883 = early_reset_static_par0_go_out;
wire _guard1884 = _guard1882 | _guard1883;
wire _guard1885 = early_reset_static_par0_go_out;
wire _guard1886 = fsm0_out == 5'd0;
wire _guard1887 = early_reset_static_seq_go_out;
wire _guard1888 = _guard1886 & _guard1887;
wire _guard1889 = early_reset_static_par0_go_out;
wire _guard1890 = early_reset_static_par0_go_out;
wire _guard1891 = fsm0_out == 5'd0;
wire _guard1892 = early_reset_static_seq_go_out;
wire _guard1893 = _guard1891 & _guard1892;
wire _guard1894 = early_reset_static_par0_go_out;
wire _guard1895 = _guard1893 | _guard1894;
wire _guard1896 = early_reset_static_par0_go_out;
wire _guard1897 = fsm0_out == 5'd0;
wire _guard1898 = early_reset_static_seq_go_out;
wire _guard1899 = _guard1897 & _guard1898;
wire _guard1900 = early_reset_static_par0_go_out;
wire _guard1901 = early_reset_static_par0_go_out;
wire _guard1902 = early_reset_static_par0_go_out;
wire _guard1903 = early_reset_static_par0_go_out;
wire _guard1904 = early_reset_static_par0_go_out;
wire _guard1905 = early_reset_static_par0_go_out;
wire _guard1906 = fsm0_out == 5'd0;
wire _guard1907 = early_reset_static_seq_go_out;
wire _guard1908 = _guard1906 & _guard1907;
wire _guard1909 = early_reset_static_par0_go_out;
wire _guard1910 = _guard1908 | _guard1909;
wire _guard1911 = fsm0_out == 5'd0;
wire _guard1912 = early_reset_static_seq_go_out;
wire _guard1913 = _guard1911 & _guard1912;
wire _guard1914 = early_reset_static_par0_go_out;
wire _guard1915 = early_reset_static_par0_go_out;
wire _guard1916 = early_reset_static_par0_go_out;
wire _guard1917 = early_reset_static_par0_go_out;
wire _guard1918 = early_reset_static_par0_go_out;
wire _guard1919 = early_reset_static_par0_go_out;
wire _guard1920 = ~_guard0;
wire _guard1921 = early_reset_static_par0_go_out;
wire _guard1922 = _guard1920 & _guard1921;
wire _guard1923 = early_reset_static_par0_go_out;
wire _guard1924 = early_reset_static_par0_go_out;
wire _guard1925 = ~_guard0;
wire _guard1926 = early_reset_static_par0_go_out;
wire _guard1927 = _guard1925 & _guard1926;
wire _guard1928 = early_reset_static_par0_go_out;
wire _guard1929 = early_reset_static_par0_go_out;
wire _guard1930 = ~_guard0;
wire _guard1931 = early_reset_static_par0_go_out;
wire _guard1932 = _guard1930 & _guard1931;
wire _guard1933 = early_reset_static_par0_go_out;
wire _guard1934 = early_reset_static_par0_go_out;
wire _guard1935 = early_reset_static_par0_go_out;
wire _guard1936 = ~_guard0;
wire _guard1937 = early_reset_static_par0_go_out;
wire _guard1938 = _guard1936 & _guard1937;
wire _guard1939 = early_reset_static_par0_go_out;
wire _guard1940 = ~_guard0;
wire _guard1941 = early_reset_static_par0_go_out;
wire _guard1942 = _guard1940 & _guard1941;
wire _guard1943 = early_reset_static_par0_go_out;
wire _guard1944 = early_reset_static_par0_go_out;
wire _guard1945 = early_reset_static_par0_go_out;
wire _guard1946 = ~_guard0;
wire _guard1947 = early_reset_static_par0_go_out;
wire _guard1948 = _guard1946 & _guard1947;
wire _guard1949 = early_reset_static_par0_go_out;
wire _guard1950 = early_reset_static_par0_go_out;
wire _guard1951 = early_reset_static_par0_go_out;
wire _guard1952 = early_reset_static_par0_go_out;
wire _guard1953 = early_reset_static_par0_go_out;
wire _guard1954 = early_reset_static_par0_go_out;
wire _guard1955 = early_reset_static_par0_go_out;
wire _guard1956 = early_reset_static_par0_go_out;
wire _guard1957 = early_reset_static_par0_go_out;
wire _guard1958 = early_reset_static_par0_go_out;
wire _guard1959 = early_reset_static_par0_go_out;
wire _guard1960 = ~_guard0;
wire _guard1961 = early_reset_static_par0_go_out;
wire _guard1962 = _guard1960 & _guard1961;
wire _guard1963 = early_reset_static_par0_go_out;
wire _guard1964 = ~_guard0;
wire _guard1965 = early_reset_static_par0_go_out;
wire _guard1966 = _guard1964 & _guard1965;
wire _guard1967 = early_reset_static_par0_go_out;
wire _guard1968 = ~_guard0;
wire _guard1969 = early_reset_static_par0_go_out;
wire _guard1970 = _guard1968 & _guard1969;
wire _guard1971 = early_reset_static_par0_go_out;
wire _guard1972 = early_reset_static_par0_go_out;
wire _guard1973 = early_reset_static_par0_go_out;
wire _guard1974 = early_reset_static_par0_go_out;
wire _guard1975 = early_reset_static_par0_go_out;
wire _guard1976 = ~_guard0;
wire _guard1977 = early_reset_static_par0_go_out;
wire _guard1978 = _guard1976 & _guard1977;
wire _guard1979 = early_reset_static_par0_go_out;
wire _guard1980 = ~_guard0;
wire _guard1981 = early_reset_static_par0_go_out;
wire _guard1982 = _guard1980 & _guard1981;
wire _guard1983 = early_reset_static_par0_go_out;
wire _guard1984 = early_reset_static_par0_go_out;
wire _guard1985 = early_reset_static_par0_go_out;
wire _guard1986 = early_reset_static_par0_go_out;
wire _guard1987 = early_reset_static_par0_go_out;
wire _guard1988 = early_reset_static_par0_go_out;
wire _guard1989 = early_reset_static_par0_go_out;
wire _guard1990 = ~_guard0;
wire _guard1991 = early_reset_static_par0_go_out;
wire _guard1992 = _guard1990 & _guard1991;
wire _guard1993 = cond_wire7_out;
wire _guard1994 = early_reset_static_par0_go_out;
wire _guard1995 = _guard1993 & _guard1994;
wire _guard1996 = cond_wire5_out;
wire _guard1997 = early_reset_static_par0_go_out;
wire _guard1998 = _guard1996 & _guard1997;
wire _guard1999 = fsm_out == 1'd0;
wire _guard2000 = cond_wire5_out;
wire _guard2001 = _guard1999 & _guard2000;
wire _guard2002 = fsm_out == 1'd0;
wire _guard2003 = _guard2001 & _guard2002;
wire _guard2004 = fsm_out == 1'd0;
wire _guard2005 = cond_wire7_out;
wire _guard2006 = _guard2004 & _guard2005;
wire _guard2007 = fsm_out == 1'd0;
wire _guard2008 = _guard2006 & _guard2007;
wire _guard2009 = _guard2003 | _guard2008;
wire _guard2010 = early_reset_static_par0_go_out;
wire _guard2011 = _guard2009 & _guard2010;
wire _guard2012 = fsm_out == 1'd0;
wire _guard2013 = cond_wire5_out;
wire _guard2014 = _guard2012 & _guard2013;
wire _guard2015 = fsm_out == 1'd0;
wire _guard2016 = _guard2014 & _guard2015;
wire _guard2017 = fsm_out == 1'd0;
wire _guard2018 = cond_wire7_out;
wire _guard2019 = _guard2017 & _guard2018;
wire _guard2020 = fsm_out == 1'd0;
wire _guard2021 = _guard2019 & _guard2020;
wire _guard2022 = _guard2016 | _guard2021;
wire _guard2023 = early_reset_static_par0_go_out;
wire _guard2024 = _guard2022 & _guard2023;
wire _guard2025 = fsm_out == 1'd0;
wire _guard2026 = cond_wire5_out;
wire _guard2027 = _guard2025 & _guard2026;
wire _guard2028 = fsm_out == 1'd0;
wire _guard2029 = _guard2027 & _guard2028;
wire _guard2030 = fsm_out == 1'd0;
wire _guard2031 = cond_wire7_out;
wire _guard2032 = _guard2030 & _guard2031;
wire _guard2033 = fsm_out == 1'd0;
wire _guard2034 = _guard2032 & _guard2033;
wire _guard2035 = _guard2029 | _guard2034;
wire _guard2036 = early_reset_static_par0_go_out;
wire _guard2037 = _guard2035 & _guard2036;
wire _guard2038 = cond_wire26_out;
wire _guard2039 = early_reset_static_par0_go_out;
wire _guard2040 = _guard2038 & _guard2039;
wire _guard2041 = cond_wire26_out;
wire _guard2042 = early_reset_static_par0_go_out;
wire _guard2043 = _guard2041 & _guard2042;
wire _guard2044 = cond_wire37_out;
wire _guard2045 = early_reset_static_par0_go_out;
wire _guard2046 = _guard2044 & _guard2045;
wire _guard2047 = cond_wire35_out;
wire _guard2048 = early_reset_static_par0_go_out;
wire _guard2049 = _guard2047 & _guard2048;
wire _guard2050 = fsm_out == 1'd0;
wire _guard2051 = cond_wire35_out;
wire _guard2052 = _guard2050 & _guard2051;
wire _guard2053 = fsm_out == 1'd0;
wire _guard2054 = _guard2052 & _guard2053;
wire _guard2055 = fsm_out == 1'd0;
wire _guard2056 = cond_wire37_out;
wire _guard2057 = _guard2055 & _guard2056;
wire _guard2058 = fsm_out == 1'd0;
wire _guard2059 = _guard2057 & _guard2058;
wire _guard2060 = _guard2054 | _guard2059;
wire _guard2061 = early_reset_static_par0_go_out;
wire _guard2062 = _guard2060 & _guard2061;
wire _guard2063 = fsm_out == 1'd0;
wire _guard2064 = cond_wire35_out;
wire _guard2065 = _guard2063 & _guard2064;
wire _guard2066 = fsm_out == 1'd0;
wire _guard2067 = _guard2065 & _guard2066;
wire _guard2068 = fsm_out == 1'd0;
wire _guard2069 = cond_wire37_out;
wire _guard2070 = _guard2068 & _guard2069;
wire _guard2071 = fsm_out == 1'd0;
wire _guard2072 = _guard2070 & _guard2071;
wire _guard2073 = _guard2067 | _guard2072;
wire _guard2074 = early_reset_static_par0_go_out;
wire _guard2075 = _guard2073 & _guard2074;
wire _guard2076 = fsm_out == 1'd0;
wire _guard2077 = cond_wire35_out;
wire _guard2078 = _guard2076 & _guard2077;
wire _guard2079 = fsm_out == 1'd0;
wire _guard2080 = _guard2078 & _guard2079;
wire _guard2081 = fsm_out == 1'd0;
wire _guard2082 = cond_wire37_out;
wire _guard2083 = _guard2081 & _guard2082;
wire _guard2084 = fsm_out == 1'd0;
wire _guard2085 = _guard2083 & _guard2084;
wire _guard2086 = _guard2080 | _guard2085;
wire _guard2087 = early_reset_static_par0_go_out;
wire _guard2088 = _guard2086 & _guard2087;
wire _guard2089 = cond_wire45_out;
wire _guard2090 = early_reset_static_par0_go_out;
wire _guard2091 = _guard2089 & _guard2090;
wire _guard2092 = cond_wire45_out;
wire _guard2093 = early_reset_static_par0_go_out;
wire _guard2094 = _guard2092 & _guard2093;
wire _guard2095 = cond_wire78_out;
wire _guard2096 = early_reset_static_par0_go_out;
wire _guard2097 = _guard2095 & _guard2096;
wire _guard2098 = cond_wire78_out;
wire _guard2099 = early_reset_static_par0_go_out;
wire _guard2100 = _guard2098 & _guard2099;
wire _guard2101 = cond_wire61_out;
wire _guard2102 = early_reset_static_par0_go_out;
wire _guard2103 = _guard2101 & _guard2102;
wire _guard2104 = cond_wire61_out;
wire _guard2105 = early_reset_static_par0_go_out;
wire _guard2106 = _guard2104 & _guard2105;
wire _guard2107 = cond_wire103_out;
wire _guard2108 = early_reset_static_par0_go_out;
wire _guard2109 = _guard2107 & _guard2108;
wire _guard2110 = cond_wire101_out;
wire _guard2111 = early_reset_static_par0_go_out;
wire _guard2112 = _guard2110 & _guard2111;
wire _guard2113 = fsm_out == 1'd0;
wire _guard2114 = cond_wire101_out;
wire _guard2115 = _guard2113 & _guard2114;
wire _guard2116 = fsm_out == 1'd0;
wire _guard2117 = _guard2115 & _guard2116;
wire _guard2118 = fsm_out == 1'd0;
wire _guard2119 = cond_wire103_out;
wire _guard2120 = _guard2118 & _guard2119;
wire _guard2121 = fsm_out == 1'd0;
wire _guard2122 = _guard2120 & _guard2121;
wire _guard2123 = _guard2117 | _guard2122;
wire _guard2124 = early_reset_static_par0_go_out;
wire _guard2125 = _guard2123 & _guard2124;
wire _guard2126 = fsm_out == 1'd0;
wire _guard2127 = cond_wire101_out;
wire _guard2128 = _guard2126 & _guard2127;
wire _guard2129 = fsm_out == 1'd0;
wire _guard2130 = _guard2128 & _guard2129;
wire _guard2131 = fsm_out == 1'd0;
wire _guard2132 = cond_wire103_out;
wire _guard2133 = _guard2131 & _guard2132;
wire _guard2134 = fsm_out == 1'd0;
wire _guard2135 = _guard2133 & _guard2134;
wire _guard2136 = _guard2130 | _guard2135;
wire _guard2137 = early_reset_static_par0_go_out;
wire _guard2138 = _guard2136 & _guard2137;
wire _guard2139 = fsm_out == 1'd0;
wire _guard2140 = cond_wire101_out;
wire _guard2141 = _guard2139 & _guard2140;
wire _guard2142 = fsm_out == 1'd0;
wire _guard2143 = _guard2141 & _guard2142;
wire _guard2144 = fsm_out == 1'd0;
wire _guard2145 = cond_wire103_out;
wire _guard2146 = _guard2144 & _guard2145;
wire _guard2147 = fsm_out == 1'd0;
wire _guard2148 = _guard2146 & _guard2147;
wire _guard2149 = _guard2143 | _guard2148;
wire _guard2150 = early_reset_static_par0_go_out;
wire _guard2151 = _guard2149 & _guard2150;
wire _guard2152 = cond_wire98_out;
wire _guard2153 = early_reset_static_par0_go_out;
wire _guard2154 = _guard2152 & _guard2153;
wire _guard2155 = cond_wire98_out;
wire _guard2156 = early_reset_static_par0_go_out;
wire _guard2157 = _guard2155 & _guard2156;
wire _guard2158 = cond_wire161_out;
wire _guard2159 = early_reset_static_par0_go_out;
wire _guard2160 = _guard2158 & _guard2159;
wire _guard2161 = cond_wire159_out;
wire _guard2162 = early_reset_static_par0_go_out;
wire _guard2163 = _guard2161 & _guard2162;
wire _guard2164 = fsm_out == 1'd0;
wire _guard2165 = cond_wire159_out;
wire _guard2166 = _guard2164 & _guard2165;
wire _guard2167 = fsm_out == 1'd0;
wire _guard2168 = _guard2166 & _guard2167;
wire _guard2169 = fsm_out == 1'd0;
wire _guard2170 = cond_wire161_out;
wire _guard2171 = _guard2169 & _guard2170;
wire _guard2172 = fsm_out == 1'd0;
wire _guard2173 = _guard2171 & _guard2172;
wire _guard2174 = _guard2168 | _guard2173;
wire _guard2175 = early_reset_static_par0_go_out;
wire _guard2176 = _guard2174 & _guard2175;
wire _guard2177 = fsm_out == 1'd0;
wire _guard2178 = cond_wire159_out;
wire _guard2179 = _guard2177 & _guard2178;
wire _guard2180 = fsm_out == 1'd0;
wire _guard2181 = _guard2179 & _guard2180;
wire _guard2182 = fsm_out == 1'd0;
wire _guard2183 = cond_wire161_out;
wire _guard2184 = _guard2182 & _guard2183;
wire _guard2185 = fsm_out == 1'd0;
wire _guard2186 = _guard2184 & _guard2185;
wire _guard2187 = _guard2181 | _guard2186;
wire _guard2188 = early_reset_static_par0_go_out;
wire _guard2189 = _guard2187 & _guard2188;
wire _guard2190 = fsm_out == 1'd0;
wire _guard2191 = cond_wire159_out;
wire _guard2192 = _guard2190 & _guard2191;
wire _guard2193 = fsm_out == 1'd0;
wire _guard2194 = _guard2192 & _guard2193;
wire _guard2195 = fsm_out == 1'd0;
wire _guard2196 = cond_wire161_out;
wire _guard2197 = _guard2195 & _guard2196;
wire _guard2198 = fsm_out == 1'd0;
wire _guard2199 = _guard2197 & _guard2198;
wire _guard2200 = _guard2194 | _guard2199;
wire _guard2201 = early_reset_static_par0_go_out;
wire _guard2202 = _guard2200 & _guard2201;
wire _guard2203 = cond_wire156_out;
wire _guard2204 = early_reset_static_par0_go_out;
wire _guard2205 = _guard2203 & _guard2204;
wire _guard2206 = cond_wire156_out;
wire _guard2207 = early_reset_static_par0_go_out;
wire _guard2208 = _guard2206 & _guard2207;
wire _guard2209 = cond_wire140_out;
wire _guard2210 = early_reset_static_par0_go_out;
wire _guard2211 = _guard2209 & _guard2210;
wire _guard2212 = cond_wire140_out;
wire _guard2213 = early_reset_static_par0_go_out;
wire _guard2214 = _guard2212 & _guard2213;
wire _guard2215 = cond_wire152_out;
wire _guard2216 = early_reset_static_par0_go_out;
wire _guard2217 = _guard2215 & _guard2216;
wire _guard2218 = cond_wire152_out;
wire _guard2219 = early_reset_static_par0_go_out;
wire _guard2220 = _guard2218 & _guard2219;
wire _guard2221 = cond_wire105_out;
wire _guard2222 = early_reset_static_par0_go_out;
wire _guard2223 = _guard2221 & _guard2222;
wire _guard2224 = cond_wire105_out;
wire _guard2225 = early_reset_static_par0_go_out;
wire _guard2226 = _guard2224 & _guard2225;
wire _guard2227 = early_reset_static_par0_go_out;
wire _guard2228 = early_reset_static_par0_go_out;
wire _guard2229 = early_reset_static_par0_go_out;
wire _guard2230 = early_reset_static_par0_go_out;
wire _guard2231 = fsm0_out == 5'd0;
wire _guard2232 = early_reset_static_seq_go_out;
wire _guard2233 = _guard2231 & _guard2232;
wire _guard2234 = early_reset_static_par0_go_out;
wire _guard2235 = _guard2233 | _guard2234;
wire _guard2236 = fsm0_out == 5'd0;
wire _guard2237 = early_reset_static_seq_go_out;
wire _guard2238 = _guard2236 & _guard2237;
wire _guard2239 = early_reset_static_par0_go_out;
wire _guard2240 = early_reset_static_par0_go_out;
wire _guard2241 = early_reset_static_par0_go_out;
wire _guard2242 = fsm0_out == 5'd0;
wire _guard2243 = early_reset_static_seq_go_out;
wire _guard2244 = _guard2242 & _guard2243;
wire _guard2245 = early_reset_static_par0_go_out;
wire _guard2246 = _guard2244 | _guard2245;
wire _guard2247 = fsm0_out == 5'd0;
wire _guard2248 = early_reset_static_seq_go_out;
wire _guard2249 = _guard2247 & _guard2248;
wire _guard2250 = early_reset_static_par0_go_out;
wire _guard2251 = early_reset_static_par0_go_out;
wire _guard2252 = early_reset_static_par0_go_out;
wire _guard2253 = early_reset_static_par0_go_out;
wire _guard2254 = early_reset_static_par0_go_out;
wire _guard2255 = early_reset_static_par0_go_out;
wire _guard2256 = early_reset_static_par0_go_out;
wire _guard2257 = early_reset_static_par0_go_out;
wire _guard2258 = early_reset_static_par0_go_out;
wire _guard2259 = early_reset_static_par0_go_out;
wire _guard2260 = early_reset_static_par0_go_out;
wire _guard2261 = early_reset_static_par0_go_out;
wire _guard2262 = early_reset_static_par0_go_out;
wire _guard2263 = early_reset_static_par0_go_out;
wire _guard2264 = early_reset_static_par0_go_out;
wire _guard2265 = early_reset_static_par0_go_out;
wire _guard2266 = ~_guard0;
wire _guard2267 = early_reset_static_par0_go_out;
wire _guard2268 = _guard2266 & _guard2267;
wire _guard2269 = early_reset_static_par0_go_out;
wire _guard2270 = early_reset_static_par0_go_out;
wire _guard2271 = ~_guard0;
wire _guard2272 = early_reset_static_par0_go_out;
wire _guard2273 = _guard2271 & _guard2272;
wire _guard2274 = early_reset_static_par0_go_out;
wire _guard2275 = ~_guard0;
wire _guard2276 = early_reset_static_par0_go_out;
wire _guard2277 = _guard2275 & _guard2276;
wire _guard2278 = early_reset_static_par0_go_out;
wire _guard2279 = early_reset_static_par0_go_out;
wire _guard2280 = ~_guard0;
wire _guard2281 = early_reset_static_par0_go_out;
wire _guard2282 = _guard2280 & _guard2281;
wire _guard2283 = early_reset_static_par0_go_out;
wire _guard2284 = early_reset_static_par0_go_out;
wire _guard2285 = early_reset_static_par0_go_out;
wire _guard2286 = early_reset_static_par0_go_out;
wire _guard2287 = early_reset_static_par0_go_out;
wire _guard2288 = early_reset_static_par0_go_out;
wire _guard2289 = early_reset_static_par0_go_out;
wire _guard2290 = early_reset_static_par0_go_out;
wire _guard2291 = early_reset_static_par0_go_out;
wire _guard2292 = ~_guard0;
wire _guard2293 = early_reset_static_par0_go_out;
wire _guard2294 = _guard2292 & _guard2293;
wire _guard2295 = early_reset_static_par0_go_out;
wire _guard2296 = early_reset_static_par0_go_out;
wire _guard2297 = early_reset_static_par0_go_out;
wire _guard2298 = ~_guard0;
wire _guard2299 = early_reset_static_par0_go_out;
wire _guard2300 = _guard2298 & _guard2299;
wire _guard2301 = early_reset_static_par0_go_out;
wire _guard2302 = ~_guard0;
wire _guard2303 = early_reset_static_par0_go_out;
wire _guard2304 = _guard2302 & _guard2303;
wire _guard2305 = ~_guard0;
wire _guard2306 = early_reset_static_par0_go_out;
wire _guard2307 = _guard2305 & _guard2306;
wire _guard2308 = early_reset_static_par0_go_out;
wire _guard2309 = early_reset_static_par0_go_out;
wire _guard2310 = ~_guard0;
wire _guard2311 = early_reset_static_par0_go_out;
wire _guard2312 = _guard2310 & _guard2311;
wire _guard2313 = early_reset_static_par0_go_out;
wire _guard2314 = early_reset_static_par0_go_out;
wire _guard2315 = ~_guard0;
wire _guard2316 = early_reset_static_par0_go_out;
wire _guard2317 = _guard2315 & _guard2316;
wire _guard2318 = early_reset_static_par0_go_out;
wire _guard2319 = early_reset_static_par0_go_out;
wire _guard2320 = ~_guard0;
wire _guard2321 = early_reset_static_par0_go_out;
wire _guard2322 = _guard2320 & _guard2321;
wire _guard2323 = early_reset_static_par0_go_out;
wire _guard2324 = ~_guard0;
wire _guard2325 = early_reset_static_par0_go_out;
wire _guard2326 = _guard2324 & _guard2325;
wire _guard2327 = early_reset_static_par0_go_out;
wire _guard2328 = early_reset_static_par0_go_out;
wire _guard2329 = early_reset_static_par0_go_out;
wire _guard2330 = early_reset_static_par0_go_out;
wire _guard2331 = early_reset_static_par0_go_out;
wire _guard2332 = early_reset_static_par0_go_out;
wire _guard2333 = ~_guard0;
wire _guard2334 = early_reset_static_par0_go_out;
wire _guard2335 = _guard2333 & _guard2334;
wire _guard2336 = early_reset_static_par0_go_out;
wire _guard2337 = ~_guard0;
wire _guard2338 = early_reset_static_par0_go_out;
wire _guard2339 = _guard2337 & _guard2338;
wire _guard2340 = early_reset_static_par0_go_out;
wire _guard2341 = early_reset_static_par0_go_out;
wire _guard2342 = early_reset_static_par0_go_out;
wire _guard2343 = early_reset_static_par0_go_out;
wire _guard2344 = early_reset_static_par0_go_out;
wire _guard2345 = ~_guard0;
wire _guard2346 = early_reset_static_par0_go_out;
wire _guard2347 = _guard2345 & _guard2346;
wire _guard2348 = early_reset_static_par0_go_out;
wire _guard2349 = early_reset_static_par0_go_out;
wire _guard2350 = early_reset_static_par0_go_out;
wire _guard2351 = cond_wire42_out;
wire _guard2352 = early_reset_static_par0_go_out;
wire _guard2353 = _guard2351 & _guard2352;
wire _guard2354 = cond_wire40_out;
wire _guard2355 = early_reset_static_par0_go_out;
wire _guard2356 = _guard2354 & _guard2355;
wire _guard2357 = fsm_out == 1'd0;
wire _guard2358 = cond_wire40_out;
wire _guard2359 = _guard2357 & _guard2358;
wire _guard2360 = fsm_out == 1'd0;
wire _guard2361 = _guard2359 & _guard2360;
wire _guard2362 = fsm_out == 1'd0;
wire _guard2363 = cond_wire42_out;
wire _guard2364 = _guard2362 & _guard2363;
wire _guard2365 = fsm_out == 1'd0;
wire _guard2366 = _guard2364 & _guard2365;
wire _guard2367 = _guard2361 | _guard2366;
wire _guard2368 = early_reset_static_par0_go_out;
wire _guard2369 = _guard2367 & _guard2368;
wire _guard2370 = fsm_out == 1'd0;
wire _guard2371 = cond_wire40_out;
wire _guard2372 = _guard2370 & _guard2371;
wire _guard2373 = fsm_out == 1'd0;
wire _guard2374 = _guard2372 & _guard2373;
wire _guard2375 = fsm_out == 1'd0;
wire _guard2376 = cond_wire42_out;
wire _guard2377 = _guard2375 & _guard2376;
wire _guard2378 = fsm_out == 1'd0;
wire _guard2379 = _guard2377 & _guard2378;
wire _guard2380 = _guard2374 | _guard2379;
wire _guard2381 = early_reset_static_par0_go_out;
wire _guard2382 = _guard2380 & _guard2381;
wire _guard2383 = fsm_out == 1'd0;
wire _guard2384 = cond_wire40_out;
wire _guard2385 = _guard2383 & _guard2384;
wire _guard2386 = fsm_out == 1'd0;
wire _guard2387 = _guard2385 & _guard2386;
wire _guard2388 = fsm_out == 1'd0;
wire _guard2389 = cond_wire42_out;
wire _guard2390 = _guard2388 & _guard2389;
wire _guard2391 = fsm_out == 1'd0;
wire _guard2392 = _guard2390 & _guard2391;
wire _guard2393 = _guard2387 | _guard2392;
wire _guard2394 = early_reset_static_par0_go_out;
wire _guard2395 = _guard2393 & _guard2394;
wire _guard2396 = cond_wire39_out;
wire _guard2397 = early_reset_static_par0_go_out;
wire _guard2398 = _guard2396 & _guard2397;
wire _guard2399 = cond_wire39_out;
wire _guard2400 = early_reset_static_par0_go_out;
wire _guard2401 = _guard2399 & _guard2400;
wire _guard2402 = cond_wire41_out;
wire _guard2403 = early_reset_static_par0_go_out;
wire _guard2404 = _guard2402 & _guard2403;
wire _guard2405 = cond_wire41_out;
wire _guard2406 = early_reset_static_par0_go_out;
wire _guard2407 = _guard2405 & _guard2406;
wire _guard2408 = cond_wire11_out;
wire _guard2409 = early_reset_static_par0_go_out;
wire _guard2410 = _guard2408 & _guard2409;
wire _guard2411 = cond_wire11_out;
wire _guard2412 = early_reset_static_par0_go_out;
wire _guard2413 = _guard2411 & _guard2412;
wire _guard2414 = cond_wire72_out;
wire _guard2415 = early_reset_static_par0_go_out;
wire _guard2416 = _guard2414 & _guard2415;
wire _guard2417 = cond_wire72_out;
wire _guard2418 = early_reset_static_par0_go_out;
wire _guard2419 = _guard2417 & _guard2418;
wire _guard2420 = cond_wire107_out;
wire _guard2421 = early_reset_static_par0_go_out;
wire _guard2422 = _guard2420 & _guard2421;
wire _guard2423 = cond_wire107_out;
wire _guard2424 = early_reset_static_par0_go_out;
wire _guard2425 = _guard2423 & _guard2424;
wire _guard2426 = cond_wire116_out;
wire _guard2427 = early_reset_static_par0_go_out;
wire _guard2428 = _guard2426 & _guard2427;
wire _guard2429 = cond_wire114_out;
wire _guard2430 = early_reset_static_par0_go_out;
wire _guard2431 = _guard2429 & _guard2430;
wire _guard2432 = fsm_out == 1'd0;
wire _guard2433 = cond_wire114_out;
wire _guard2434 = _guard2432 & _guard2433;
wire _guard2435 = fsm_out == 1'd0;
wire _guard2436 = _guard2434 & _guard2435;
wire _guard2437 = fsm_out == 1'd0;
wire _guard2438 = cond_wire116_out;
wire _guard2439 = _guard2437 & _guard2438;
wire _guard2440 = fsm_out == 1'd0;
wire _guard2441 = _guard2439 & _guard2440;
wire _guard2442 = _guard2436 | _guard2441;
wire _guard2443 = early_reset_static_par0_go_out;
wire _guard2444 = _guard2442 & _guard2443;
wire _guard2445 = fsm_out == 1'd0;
wire _guard2446 = cond_wire114_out;
wire _guard2447 = _guard2445 & _guard2446;
wire _guard2448 = fsm_out == 1'd0;
wire _guard2449 = _guard2447 & _guard2448;
wire _guard2450 = fsm_out == 1'd0;
wire _guard2451 = cond_wire116_out;
wire _guard2452 = _guard2450 & _guard2451;
wire _guard2453 = fsm_out == 1'd0;
wire _guard2454 = _guard2452 & _guard2453;
wire _guard2455 = _guard2449 | _guard2454;
wire _guard2456 = early_reset_static_par0_go_out;
wire _guard2457 = _guard2455 & _guard2456;
wire _guard2458 = fsm_out == 1'd0;
wire _guard2459 = cond_wire114_out;
wire _guard2460 = _guard2458 & _guard2459;
wire _guard2461 = fsm_out == 1'd0;
wire _guard2462 = _guard2460 & _guard2461;
wire _guard2463 = fsm_out == 1'd0;
wire _guard2464 = cond_wire116_out;
wire _guard2465 = _guard2463 & _guard2464;
wire _guard2466 = fsm_out == 1'd0;
wire _guard2467 = _guard2465 & _guard2466;
wire _guard2468 = _guard2462 | _guard2467;
wire _guard2469 = early_reset_static_par0_go_out;
wire _guard2470 = _guard2468 & _guard2469;
wire _guard2471 = cond_wire128_out;
wire _guard2472 = early_reset_static_par0_go_out;
wire _guard2473 = _guard2471 & _guard2472;
wire _guard2474 = cond_wire126_out;
wire _guard2475 = early_reset_static_par0_go_out;
wire _guard2476 = _guard2474 & _guard2475;
wire _guard2477 = fsm_out == 1'd0;
wire _guard2478 = cond_wire126_out;
wire _guard2479 = _guard2477 & _guard2478;
wire _guard2480 = fsm_out == 1'd0;
wire _guard2481 = _guard2479 & _guard2480;
wire _guard2482 = fsm_out == 1'd0;
wire _guard2483 = cond_wire128_out;
wire _guard2484 = _guard2482 & _guard2483;
wire _guard2485 = fsm_out == 1'd0;
wire _guard2486 = _guard2484 & _guard2485;
wire _guard2487 = _guard2481 | _guard2486;
wire _guard2488 = early_reset_static_par0_go_out;
wire _guard2489 = _guard2487 & _guard2488;
wire _guard2490 = fsm_out == 1'd0;
wire _guard2491 = cond_wire126_out;
wire _guard2492 = _guard2490 & _guard2491;
wire _guard2493 = fsm_out == 1'd0;
wire _guard2494 = _guard2492 & _guard2493;
wire _guard2495 = fsm_out == 1'd0;
wire _guard2496 = cond_wire128_out;
wire _guard2497 = _guard2495 & _guard2496;
wire _guard2498 = fsm_out == 1'd0;
wire _guard2499 = _guard2497 & _guard2498;
wire _guard2500 = _guard2494 | _guard2499;
wire _guard2501 = early_reset_static_par0_go_out;
wire _guard2502 = _guard2500 & _guard2501;
wire _guard2503 = fsm_out == 1'd0;
wire _guard2504 = cond_wire126_out;
wire _guard2505 = _guard2503 & _guard2504;
wire _guard2506 = fsm_out == 1'd0;
wire _guard2507 = _guard2505 & _guard2506;
wire _guard2508 = fsm_out == 1'd0;
wire _guard2509 = cond_wire128_out;
wire _guard2510 = _guard2508 & _guard2509;
wire _guard2511 = fsm_out == 1'd0;
wire _guard2512 = _guard2510 & _guard2511;
wire _guard2513 = _guard2507 | _guard2512;
wire _guard2514 = early_reset_static_par0_go_out;
wire _guard2515 = _guard2513 & _guard2514;
wire _guard2516 = cond_wire132_out;
wire _guard2517 = early_reset_static_par0_go_out;
wire _guard2518 = _guard2516 & _guard2517;
wire _guard2519 = cond_wire130_out;
wire _guard2520 = early_reset_static_par0_go_out;
wire _guard2521 = _guard2519 & _guard2520;
wire _guard2522 = fsm_out == 1'd0;
wire _guard2523 = cond_wire130_out;
wire _guard2524 = _guard2522 & _guard2523;
wire _guard2525 = fsm_out == 1'd0;
wire _guard2526 = _guard2524 & _guard2525;
wire _guard2527 = fsm_out == 1'd0;
wire _guard2528 = cond_wire132_out;
wire _guard2529 = _guard2527 & _guard2528;
wire _guard2530 = fsm_out == 1'd0;
wire _guard2531 = _guard2529 & _guard2530;
wire _guard2532 = _guard2526 | _guard2531;
wire _guard2533 = early_reset_static_par0_go_out;
wire _guard2534 = _guard2532 & _guard2533;
wire _guard2535 = fsm_out == 1'd0;
wire _guard2536 = cond_wire130_out;
wire _guard2537 = _guard2535 & _guard2536;
wire _guard2538 = fsm_out == 1'd0;
wire _guard2539 = _guard2537 & _guard2538;
wire _guard2540 = fsm_out == 1'd0;
wire _guard2541 = cond_wire132_out;
wire _guard2542 = _guard2540 & _guard2541;
wire _guard2543 = fsm_out == 1'd0;
wire _guard2544 = _guard2542 & _guard2543;
wire _guard2545 = _guard2539 | _guard2544;
wire _guard2546 = early_reset_static_par0_go_out;
wire _guard2547 = _guard2545 & _guard2546;
wire _guard2548 = fsm_out == 1'd0;
wire _guard2549 = cond_wire130_out;
wire _guard2550 = _guard2548 & _guard2549;
wire _guard2551 = fsm_out == 1'd0;
wire _guard2552 = _guard2550 & _guard2551;
wire _guard2553 = fsm_out == 1'd0;
wire _guard2554 = cond_wire132_out;
wire _guard2555 = _guard2553 & _guard2554;
wire _guard2556 = fsm_out == 1'd0;
wire _guard2557 = _guard2555 & _guard2556;
wire _guard2558 = _guard2552 | _guard2557;
wire _guard2559 = early_reset_static_par0_go_out;
wire _guard2560 = _guard2558 & _guard2559;
wire _guard2561 = cond_wire131_out;
wire _guard2562 = early_reset_static_par0_go_out;
wire _guard2563 = _guard2561 & _guard2562;
wire _guard2564 = cond_wire131_out;
wire _guard2565 = early_reset_static_par0_go_out;
wire _guard2566 = _guard2564 & _guard2565;
wire _guard2567 = cond_wire127_out;
wire _guard2568 = early_reset_static_par0_go_out;
wire _guard2569 = _guard2567 & _guard2568;
wire _guard2570 = cond_wire127_out;
wire _guard2571 = early_reset_static_par0_go_out;
wire _guard2572 = _guard2570 & _guard2571;
wire _guard2573 = cond_wire190_out;
wire _guard2574 = early_reset_static_par0_go_out;
wire _guard2575 = _guard2573 & _guard2574;
wire _guard2576 = cond_wire188_out;
wire _guard2577 = early_reset_static_par0_go_out;
wire _guard2578 = _guard2576 & _guard2577;
wire _guard2579 = fsm_out == 1'd0;
wire _guard2580 = cond_wire188_out;
wire _guard2581 = _guard2579 & _guard2580;
wire _guard2582 = fsm_out == 1'd0;
wire _guard2583 = _guard2581 & _guard2582;
wire _guard2584 = fsm_out == 1'd0;
wire _guard2585 = cond_wire190_out;
wire _guard2586 = _guard2584 & _guard2585;
wire _guard2587 = fsm_out == 1'd0;
wire _guard2588 = _guard2586 & _guard2587;
wire _guard2589 = _guard2583 | _guard2588;
wire _guard2590 = early_reset_static_par0_go_out;
wire _guard2591 = _guard2589 & _guard2590;
wire _guard2592 = fsm_out == 1'd0;
wire _guard2593 = cond_wire188_out;
wire _guard2594 = _guard2592 & _guard2593;
wire _guard2595 = fsm_out == 1'd0;
wire _guard2596 = _guard2594 & _guard2595;
wire _guard2597 = fsm_out == 1'd0;
wire _guard2598 = cond_wire190_out;
wire _guard2599 = _guard2597 & _guard2598;
wire _guard2600 = fsm_out == 1'd0;
wire _guard2601 = _guard2599 & _guard2600;
wire _guard2602 = _guard2596 | _guard2601;
wire _guard2603 = early_reset_static_par0_go_out;
wire _guard2604 = _guard2602 & _guard2603;
wire _guard2605 = fsm_out == 1'd0;
wire _guard2606 = cond_wire188_out;
wire _guard2607 = _guard2605 & _guard2606;
wire _guard2608 = fsm_out == 1'd0;
wire _guard2609 = _guard2607 & _guard2608;
wire _guard2610 = fsm_out == 1'd0;
wire _guard2611 = cond_wire190_out;
wire _guard2612 = _guard2610 & _guard2611;
wire _guard2613 = fsm_out == 1'd0;
wire _guard2614 = _guard2612 & _guard2613;
wire _guard2615 = _guard2609 | _guard2614;
wire _guard2616 = early_reset_static_par0_go_out;
wire _guard2617 = _guard2615 & _guard2616;
wire _guard2618 = cond_wire214_out;
wire _guard2619 = early_reset_static_par0_go_out;
wire _guard2620 = _guard2618 & _guard2619;
wire _guard2621 = cond_wire214_out;
wire _guard2622 = early_reset_static_par0_go_out;
wire _guard2623 = _guard2621 & _guard2622;
wire _guard2624 = cond_wire256_out;
wire _guard2625 = early_reset_static_par0_go_out;
wire _guard2626 = _guard2624 & _guard2625;
wire _guard2627 = cond_wire254_out;
wire _guard2628 = early_reset_static_par0_go_out;
wire _guard2629 = _guard2627 & _guard2628;
wire _guard2630 = fsm_out == 1'd0;
wire _guard2631 = cond_wire254_out;
wire _guard2632 = _guard2630 & _guard2631;
wire _guard2633 = fsm_out == 1'd0;
wire _guard2634 = _guard2632 & _guard2633;
wire _guard2635 = fsm_out == 1'd0;
wire _guard2636 = cond_wire256_out;
wire _guard2637 = _guard2635 & _guard2636;
wire _guard2638 = fsm_out == 1'd0;
wire _guard2639 = _guard2637 & _guard2638;
wire _guard2640 = _guard2634 | _guard2639;
wire _guard2641 = early_reset_static_par0_go_out;
wire _guard2642 = _guard2640 & _guard2641;
wire _guard2643 = fsm_out == 1'd0;
wire _guard2644 = cond_wire254_out;
wire _guard2645 = _guard2643 & _guard2644;
wire _guard2646 = fsm_out == 1'd0;
wire _guard2647 = _guard2645 & _guard2646;
wire _guard2648 = fsm_out == 1'd0;
wire _guard2649 = cond_wire256_out;
wire _guard2650 = _guard2648 & _guard2649;
wire _guard2651 = fsm_out == 1'd0;
wire _guard2652 = _guard2650 & _guard2651;
wire _guard2653 = _guard2647 | _guard2652;
wire _guard2654 = early_reset_static_par0_go_out;
wire _guard2655 = _guard2653 & _guard2654;
wire _guard2656 = fsm_out == 1'd0;
wire _guard2657 = cond_wire254_out;
wire _guard2658 = _guard2656 & _guard2657;
wire _guard2659 = fsm_out == 1'd0;
wire _guard2660 = _guard2658 & _guard2659;
wire _guard2661 = fsm_out == 1'd0;
wire _guard2662 = cond_wire256_out;
wire _guard2663 = _guard2661 & _guard2662;
wire _guard2664 = fsm_out == 1'd0;
wire _guard2665 = _guard2663 & _guard2664;
wire _guard2666 = _guard2660 | _guard2665;
wire _guard2667 = early_reset_static_par0_go_out;
wire _guard2668 = _guard2666 & _guard2667;
wire _guard2669 = fsm0_out == 5'd0;
wire _guard2670 = early_reset_static_seq_go_out;
wire _guard2671 = _guard2669 & _guard2670;
wire _guard2672 = cond_wire4_out;
wire _guard2673 = early_reset_static_par0_go_out;
wire _guard2674 = _guard2672 & _guard2673;
wire _guard2675 = _guard2671 | _guard2674;
wire _guard2676 = fsm0_out == 5'd0;
wire _guard2677 = early_reset_static_seq_go_out;
wire _guard2678 = _guard2676 & _guard2677;
wire _guard2679 = cond_wire4_out;
wire _guard2680 = early_reset_static_par0_go_out;
wire _guard2681 = _guard2679 & _guard2680;
wire _guard2682 = fsm0_out == 5'd0;
wire _guard2683 = early_reset_static_seq_go_out;
wire _guard2684 = _guard2682 & _guard2683;
wire _guard2685 = cond_wire34_out;
wire _guard2686 = early_reset_static_par0_go_out;
wire _guard2687 = _guard2685 & _guard2686;
wire _guard2688 = _guard2684 | _guard2687;
wire _guard2689 = fsm0_out == 5'd0;
wire _guard2690 = early_reset_static_seq_go_out;
wire _guard2691 = _guard2689 & _guard2690;
wire _guard2692 = cond_wire34_out;
wire _guard2693 = early_reset_static_par0_go_out;
wire _guard2694 = _guard2692 & _guard2693;
wire _guard2695 = early_reset_static_par0_go_out;
wire _guard2696 = early_reset_static_par0_go_out;
wire _guard2697 = early_reset_static_par0_go_out;
wire _guard2698 = early_reset_static_par0_go_out;
wire _guard2699 = fsm0_out == 5'd0;
wire _guard2700 = early_reset_static_seq_go_out;
wire _guard2701 = _guard2699 & _guard2700;
wire _guard2702 = early_reset_static_par0_go_out;
wire _guard2703 = _guard2701 | _guard2702;
wire _guard2704 = fsm0_out == 5'd0;
wire _guard2705 = early_reset_static_seq_go_out;
wire _guard2706 = _guard2704 & _guard2705;
wire _guard2707 = early_reset_static_par0_go_out;
wire _guard2708 = fsm0_out == 5'd0;
wire _guard2709 = early_reset_static_seq_go_out;
wire _guard2710 = _guard2708 & _guard2709;
wire _guard2711 = early_reset_static_par0_go_out;
wire _guard2712 = _guard2710 | _guard2711;
wire _guard2713 = early_reset_static_par0_go_out;
wire _guard2714 = fsm0_out == 5'd0;
wire _guard2715 = early_reset_static_seq_go_out;
wire _guard2716 = _guard2714 & _guard2715;
wire _guard2717 = early_reset_static_par0_go_out;
wire _guard2718 = early_reset_static_par0_go_out;
wire _guard2719 = early_reset_static_par0_go_out;
wire _guard2720 = early_reset_static_par0_go_out;
wire _guard2721 = early_reset_static_par0_go_out;
wire _guard2722 = early_reset_static_par0_go_out;
wire _guard2723 = early_reset_static_par0_go_out;
wire _guard2724 = ~_guard0;
wire _guard2725 = early_reset_static_par0_go_out;
wire _guard2726 = _guard2724 & _guard2725;
wire _guard2727 = early_reset_static_par0_go_out;
wire _guard2728 = ~_guard0;
wire _guard2729 = early_reset_static_par0_go_out;
wire _guard2730 = _guard2728 & _guard2729;
wire _guard2731 = early_reset_static_par0_go_out;
wire _guard2732 = ~_guard0;
wire _guard2733 = early_reset_static_par0_go_out;
wire _guard2734 = _guard2732 & _guard2733;
wire _guard2735 = early_reset_static_par0_go_out;
wire _guard2736 = ~_guard0;
wire _guard2737 = early_reset_static_par0_go_out;
wire _guard2738 = _guard2736 & _guard2737;
wire _guard2739 = ~_guard0;
wire _guard2740 = early_reset_static_par0_go_out;
wire _guard2741 = _guard2739 & _guard2740;
wire _guard2742 = early_reset_static_par0_go_out;
wire _guard2743 = early_reset_static_par0_go_out;
wire _guard2744 = ~_guard0;
wire _guard2745 = early_reset_static_par0_go_out;
wire _guard2746 = _guard2744 & _guard2745;
wire _guard2747 = ~_guard0;
wire _guard2748 = early_reset_static_par0_go_out;
wire _guard2749 = _guard2747 & _guard2748;
wire _guard2750 = early_reset_static_par0_go_out;
wire _guard2751 = early_reset_static_par0_go_out;
wire _guard2752 = early_reset_static_par0_go_out;
wire _guard2753 = ~_guard0;
wire _guard2754 = early_reset_static_par0_go_out;
wire _guard2755 = _guard2753 & _guard2754;
wire _guard2756 = early_reset_static_par0_go_out;
wire _guard2757 = early_reset_static_par0_go_out;
wire _guard2758 = early_reset_static_par0_go_out;
wire _guard2759 = ~_guard0;
wire _guard2760 = early_reset_static_par0_go_out;
wire _guard2761 = _guard2759 & _guard2760;
wire _guard2762 = early_reset_static_par0_go_out;
wire _guard2763 = early_reset_static_par0_go_out;
wire _guard2764 = early_reset_static_par0_go_out;
wire _guard2765 = early_reset_static_par0_go_out;
wire _guard2766 = ~_guard0;
wire _guard2767 = early_reset_static_par0_go_out;
wire _guard2768 = _guard2766 & _guard2767;
wire _guard2769 = ~_guard0;
wire _guard2770 = early_reset_static_par0_go_out;
wire _guard2771 = _guard2769 & _guard2770;
wire _guard2772 = early_reset_static_par0_go_out;
wire _guard2773 = early_reset_static_par0_go_out;
wire _guard2774 = ~_guard0;
wire _guard2775 = early_reset_static_par0_go_out;
wire _guard2776 = _guard2774 & _guard2775;
wire _guard2777 = early_reset_static_par0_go_out;
wire _guard2778 = early_reset_static_par0_go_out;
wire _guard2779 = early_reset_static_par0_go_out;
wire _guard2780 = early_reset_static_par0_go_out;
wire _guard2781 = early_reset_static_par0_go_out;
wire _guard2782 = ~_guard0;
wire _guard2783 = early_reset_static_par0_go_out;
wire _guard2784 = _guard2782 & _guard2783;
wire _guard2785 = ~_guard0;
wire _guard2786 = early_reset_static_par0_go_out;
wire _guard2787 = _guard2785 & _guard2786;
wire _guard2788 = early_reset_static_par0_go_out;
wire _guard2789 = early_reset_static_par0_go_out;
wire _guard2790 = early_reset_static_par0_go_out;
wire _guard2791 = early_reset_static_par0_go_out;
wire _guard2792 = early_reset_static_par0_go_out;
wire _guard2793 = ~_guard0;
wire _guard2794 = early_reset_static_par0_go_out;
wire _guard2795 = _guard2793 & _guard2794;
wire _guard2796 = early_reset_static_par0_go_out;
wire _guard2797 = ~_guard0;
wire _guard2798 = early_reset_static_par0_go_out;
wire _guard2799 = _guard2797 & _guard2798;
wire _guard2800 = early_reset_static_par0_go_out;
wire _guard2801 = early_reset_static_par0_go_out;
wire _guard2802 = early_reset_static_par0_go_out;
wire _guard2803 = ~_guard0;
wire _guard2804 = early_reset_static_par0_go_out;
wire _guard2805 = _guard2803 & _guard2804;
wire _guard2806 = early_reset_static_par0_go_out;
wire _guard2807 = early_reset_static_par0_go_out;
wire _guard2808 = early_reset_static_par0_go_out;
wire _guard2809 = cond_wire_out;
wire _guard2810 = early_reset_static_par0_go_out;
wire _guard2811 = _guard2809 & _guard2810;
wire _guard2812 = cond_wire_out;
wire _guard2813 = early_reset_static_par0_go_out;
wire _guard2814 = _guard2812 & _guard2813;
wire _guard2815 = cond_wire17_out;
wire _guard2816 = early_reset_static_par0_go_out;
wire _guard2817 = _guard2815 & _guard2816;
wire _guard2818 = cond_wire15_out;
wire _guard2819 = early_reset_static_par0_go_out;
wire _guard2820 = _guard2818 & _guard2819;
wire _guard2821 = fsm_out == 1'd0;
wire _guard2822 = cond_wire15_out;
wire _guard2823 = _guard2821 & _guard2822;
wire _guard2824 = fsm_out == 1'd0;
wire _guard2825 = _guard2823 & _guard2824;
wire _guard2826 = fsm_out == 1'd0;
wire _guard2827 = cond_wire17_out;
wire _guard2828 = _guard2826 & _guard2827;
wire _guard2829 = fsm_out == 1'd0;
wire _guard2830 = _guard2828 & _guard2829;
wire _guard2831 = _guard2825 | _guard2830;
wire _guard2832 = early_reset_static_par0_go_out;
wire _guard2833 = _guard2831 & _guard2832;
wire _guard2834 = fsm_out == 1'd0;
wire _guard2835 = cond_wire15_out;
wire _guard2836 = _guard2834 & _guard2835;
wire _guard2837 = fsm_out == 1'd0;
wire _guard2838 = _guard2836 & _guard2837;
wire _guard2839 = fsm_out == 1'd0;
wire _guard2840 = cond_wire17_out;
wire _guard2841 = _guard2839 & _guard2840;
wire _guard2842 = fsm_out == 1'd0;
wire _guard2843 = _guard2841 & _guard2842;
wire _guard2844 = _guard2838 | _guard2843;
wire _guard2845 = early_reset_static_par0_go_out;
wire _guard2846 = _guard2844 & _guard2845;
wire _guard2847 = fsm_out == 1'd0;
wire _guard2848 = cond_wire15_out;
wire _guard2849 = _guard2847 & _guard2848;
wire _guard2850 = fsm_out == 1'd0;
wire _guard2851 = _guard2849 & _guard2850;
wire _guard2852 = fsm_out == 1'd0;
wire _guard2853 = cond_wire17_out;
wire _guard2854 = _guard2852 & _guard2853;
wire _guard2855 = fsm_out == 1'd0;
wire _guard2856 = _guard2854 & _guard2855;
wire _guard2857 = _guard2851 | _guard2856;
wire _guard2858 = early_reset_static_par0_go_out;
wire _guard2859 = _guard2857 & _guard2858;
wire _guard2860 = cond_wire27_out;
wire _guard2861 = early_reset_static_par0_go_out;
wire _guard2862 = _guard2860 & _guard2861;
wire _guard2863 = cond_wire25_out;
wire _guard2864 = early_reset_static_par0_go_out;
wire _guard2865 = _guard2863 & _guard2864;
wire _guard2866 = fsm_out == 1'd0;
wire _guard2867 = cond_wire25_out;
wire _guard2868 = _guard2866 & _guard2867;
wire _guard2869 = fsm_out == 1'd0;
wire _guard2870 = _guard2868 & _guard2869;
wire _guard2871 = fsm_out == 1'd0;
wire _guard2872 = cond_wire27_out;
wire _guard2873 = _guard2871 & _guard2872;
wire _guard2874 = fsm_out == 1'd0;
wire _guard2875 = _guard2873 & _guard2874;
wire _guard2876 = _guard2870 | _guard2875;
wire _guard2877 = early_reset_static_par0_go_out;
wire _guard2878 = _guard2876 & _guard2877;
wire _guard2879 = fsm_out == 1'd0;
wire _guard2880 = cond_wire25_out;
wire _guard2881 = _guard2879 & _guard2880;
wire _guard2882 = fsm_out == 1'd0;
wire _guard2883 = _guard2881 & _guard2882;
wire _guard2884 = fsm_out == 1'd0;
wire _guard2885 = cond_wire27_out;
wire _guard2886 = _guard2884 & _guard2885;
wire _guard2887 = fsm_out == 1'd0;
wire _guard2888 = _guard2886 & _guard2887;
wire _guard2889 = _guard2883 | _guard2888;
wire _guard2890 = early_reset_static_par0_go_out;
wire _guard2891 = _guard2889 & _guard2890;
wire _guard2892 = fsm_out == 1'd0;
wire _guard2893 = cond_wire25_out;
wire _guard2894 = _guard2892 & _guard2893;
wire _guard2895 = fsm_out == 1'd0;
wire _guard2896 = _guard2894 & _guard2895;
wire _guard2897 = fsm_out == 1'd0;
wire _guard2898 = cond_wire27_out;
wire _guard2899 = _guard2897 & _guard2898;
wire _guard2900 = fsm_out == 1'd0;
wire _guard2901 = _guard2899 & _guard2900;
wire _guard2902 = _guard2896 | _guard2901;
wire _guard2903 = early_reset_static_par0_go_out;
wire _guard2904 = _guard2902 & _guard2903;
wire _guard2905 = cond_wire16_out;
wire _guard2906 = early_reset_static_par0_go_out;
wire _guard2907 = _guard2905 & _guard2906;
wire _guard2908 = cond_wire16_out;
wire _guard2909 = early_reset_static_par0_go_out;
wire _guard2910 = _guard2908 & _guard2909;
wire _guard2911 = cond_wire21_out;
wire _guard2912 = early_reset_static_par0_go_out;
wire _guard2913 = _guard2911 & _guard2912;
wire _guard2914 = cond_wire21_out;
wire _guard2915 = early_reset_static_par0_go_out;
wire _guard2916 = _guard2914 & _guard2915;
wire _guard2917 = cond_wire82_out;
wire _guard2918 = early_reset_static_par0_go_out;
wire _guard2919 = _guard2917 & _guard2918;
wire _guard2920 = cond_wire82_out;
wire _guard2921 = early_reset_static_par0_go_out;
wire _guard2922 = _guard2920 & _guard2921;
wire _guard2923 = cond_wire91_out;
wire _guard2924 = early_reset_static_par0_go_out;
wire _guard2925 = _guard2923 & _guard2924;
wire _guard2926 = cond_wire89_out;
wire _guard2927 = early_reset_static_par0_go_out;
wire _guard2928 = _guard2926 & _guard2927;
wire _guard2929 = fsm_out == 1'd0;
wire _guard2930 = cond_wire89_out;
wire _guard2931 = _guard2929 & _guard2930;
wire _guard2932 = fsm_out == 1'd0;
wire _guard2933 = _guard2931 & _guard2932;
wire _guard2934 = fsm_out == 1'd0;
wire _guard2935 = cond_wire91_out;
wire _guard2936 = _guard2934 & _guard2935;
wire _guard2937 = fsm_out == 1'd0;
wire _guard2938 = _guard2936 & _guard2937;
wire _guard2939 = _guard2933 | _guard2938;
wire _guard2940 = early_reset_static_par0_go_out;
wire _guard2941 = _guard2939 & _guard2940;
wire _guard2942 = fsm_out == 1'd0;
wire _guard2943 = cond_wire89_out;
wire _guard2944 = _guard2942 & _guard2943;
wire _guard2945 = fsm_out == 1'd0;
wire _guard2946 = _guard2944 & _guard2945;
wire _guard2947 = fsm_out == 1'd0;
wire _guard2948 = cond_wire91_out;
wire _guard2949 = _guard2947 & _guard2948;
wire _guard2950 = fsm_out == 1'd0;
wire _guard2951 = _guard2949 & _guard2950;
wire _guard2952 = _guard2946 | _guard2951;
wire _guard2953 = early_reset_static_par0_go_out;
wire _guard2954 = _guard2952 & _guard2953;
wire _guard2955 = fsm_out == 1'd0;
wire _guard2956 = cond_wire89_out;
wire _guard2957 = _guard2955 & _guard2956;
wire _guard2958 = fsm_out == 1'd0;
wire _guard2959 = _guard2957 & _guard2958;
wire _guard2960 = fsm_out == 1'd0;
wire _guard2961 = cond_wire91_out;
wire _guard2962 = _guard2960 & _guard2961;
wire _guard2963 = fsm_out == 1'd0;
wire _guard2964 = _guard2962 & _guard2963;
wire _guard2965 = _guard2959 | _guard2964;
wire _guard2966 = early_reset_static_par0_go_out;
wire _guard2967 = _guard2965 & _guard2966;
wire _guard2968 = cond_wire65_out;
wire _guard2969 = early_reset_static_par0_go_out;
wire _guard2970 = _guard2968 & _guard2969;
wire _guard2971 = cond_wire65_out;
wire _guard2972 = early_reset_static_par0_go_out;
wire _guard2973 = _guard2971 & _guard2972;
wire _guard2974 = cond_wire108_out;
wire _guard2975 = early_reset_static_par0_go_out;
wire _guard2976 = _guard2974 & _guard2975;
wire _guard2977 = cond_wire106_out;
wire _guard2978 = early_reset_static_par0_go_out;
wire _guard2979 = _guard2977 & _guard2978;
wire _guard2980 = fsm_out == 1'd0;
wire _guard2981 = cond_wire106_out;
wire _guard2982 = _guard2980 & _guard2981;
wire _guard2983 = fsm_out == 1'd0;
wire _guard2984 = _guard2982 & _guard2983;
wire _guard2985 = fsm_out == 1'd0;
wire _guard2986 = cond_wire108_out;
wire _guard2987 = _guard2985 & _guard2986;
wire _guard2988 = fsm_out == 1'd0;
wire _guard2989 = _guard2987 & _guard2988;
wire _guard2990 = _guard2984 | _guard2989;
wire _guard2991 = early_reset_static_par0_go_out;
wire _guard2992 = _guard2990 & _guard2991;
wire _guard2993 = fsm_out == 1'd0;
wire _guard2994 = cond_wire106_out;
wire _guard2995 = _guard2993 & _guard2994;
wire _guard2996 = fsm_out == 1'd0;
wire _guard2997 = _guard2995 & _guard2996;
wire _guard2998 = fsm_out == 1'd0;
wire _guard2999 = cond_wire108_out;
wire _guard3000 = _guard2998 & _guard2999;
wire _guard3001 = fsm_out == 1'd0;
wire _guard3002 = _guard3000 & _guard3001;
wire _guard3003 = _guard2997 | _guard3002;
wire _guard3004 = early_reset_static_par0_go_out;
wire _guard3005 = _guard3003 & _guard3004;
wire _guard3006 = fsm_out == 1'd0;
wire _guard3007 = cond_wire106_out;
wire _guard3008 = _guard3006 & _guard3007;
wire _guard3009 = fsm_out == 1'd0;
wire _guard3010 = _guard3008 & _guard3009;
wire _guard3011 = fsm_out == 1'd0;
wire _guard3012 = cond_wire108_out;
wire _guard3013 = _guard3011 & _guard3012;
wire _guard3014 = fsm_out == 1'd0;
wire _guard3015 = _guard3013 & _guard3014;
wire _guard3016 = _guard3010 | _guard3015;
wire _guard3017 = early_reset_static_par0_go_out;
wire _guard3018 = _guard3016 & _guard3017;
wire _guard3019 = cond_wire82_out;
wire _guard3020 = early_reset_static_par0_go_out;
wire _guard3021 = _guard3019 & _guard3020;
wire _guard3022 = cond_wire82_out;
wire _guard3023 = early_reset_static_par0_go_out;
wire _guard3024 = _guard3022 & _guard3023;
wire _guard3025 = cond_wire107_out;
wire _guard3026 = early_reset_static_par0_go_out;
wire _guard3027 = _guard3025 & _guard3026;
wire _guard3028 = cond_wire107_out;
wire _guard3029 = early_reset_static_par0_go_out;
wire _guard3030 = _guard3028 & _guard3029;
wire _guard3031 = cond_wire160_out;
wire _guard3032 = early_reset_static_par0_go_out;
wire _guard3033 = _guard3031 & _guard3032;
wire _guard3034 = cond_wire160_out;
wire _guard3035 = early_reset_static_par0_go_out;
wire _guard3036 = _guard3034 & _guard3035;
wire _guard3037 = cond_wire164_out;
wire _guard3038 = early_reset_static_par0_go_out;
wire _guard3039 = _guard3037 & _guard3038;
wire _guard3040 = cond_wire164_out;
wire _guard3041 = early_reset_static_par0_go_out;
wire _guard3042 = _guard3040 & _guard3041;
wire _guard3043 = cond_wire178_out;
wire _guard3044 = early_reset_static_par0_go_out;
wire _guard3045 = _guard3043 & _guard3044;
wire _guard3046 = cond_wire176_out;
wire _guard3047 = early_reset_static_par0_go_out;
wire _guard3048 = _guard3046 & _guard3047;
wire _guard3049 = fsm_out == 1'd0;
wire _guard3050 = cond_wire176_out;
wire _guard3051 = _guard3049 & _guard3050;
wire _guard3052 = fsm_out == 1'd0;
wire _guard3053 = _guard3051 & _guard3052;
wire _guard3054 = fsm_out == 1'd0;
wire _guard3055 = cond_wire178_out;
wire _guard3056 = _guard3054 & _guard3055;
wire _guard3057 = fsm_out == 1'd0;
wire _guard3058 = _guard3056 & _guard3057;
wire _guard3059 = _guard3053 | _guard3058;
wire _guard3060 = early_reset_static_par0_go_out;
wire _guard3061 = _guard3059 & _guard3060;
wire _guard3062 = fsm_out == 1'd0;
wire _guard3063 = cond_wire176_out;
wire _guard3064 = _guard3062 & _guard3063;
wire _guard3065 = fsm_out == 1'd0;
wire _guard3066 = _guard3064 & _guard3065;
wire _guard3067 = fsm_out == 1'd0;
wire _guard3068 = cond_wire178_out;
wire _guard3069 = _guard3067 & _guard3068;
wire _guard3070 = fsm_out == 1'd0;
wire _guard3071 = _guard3069 & _guard3070;
wire _guard3072 = _guard3066 | _guard3071;
wire _guard3073 = early_reset_static_par0_go_out;
wire _guard3074 = _guard3072 & _guard3073;
wire _guard3075 = fsm_out == 1'd0;
wire _guard3076 = cond_wire176_out;
wire _guard3077 = _guard3075 & _guard3076;
wire _guard3078 = fsm_out == 1'd0;
wire _guard3079 = _guard3077 & _guard3078;
wire _guard3080 = fsm_out == 1'd0;
wire _guard3081 = cond_wire178_out;
wire _guard3082 = _guard3080 & _guard3081;
wire _guard3083 = fsm_out == 1'd0;
wire _guard3084 = _guard3082 & _guard3083;
wire _guard3085 = _guard3079 | _guard3084;
wire _guard3086 = early_reset_static_par0_go_out;
wire _guard3087 = _guard3085 & _guard3086;
wire _guard3088 = cond_wire202_out;
wire _guard3089 = early_reset_static_par0_go_out;
wire _guard3090 = _guard3088 & _guard3089;
wire _guard3091 = cond_wire200_out;
wire _guard3092 = early_reset_static_par0_go_out;
wire _guard3093 = _guard3091 & _guard3092;
wire _guard3094 = fsm_out == 1'd0;
wire _guard3095 = cond_wire200_out;
wire _guard3096 = _guard3094 & _guard3095;
wire _guard3097 = fsm_out == 1'd0;
wire _guard3098 = _guard3096 & _guard3097;
wire _guard3099 = fsm_out == 1'd0;
wire _guard3100 = cond_wire202_out;
wire _guard3101 = _guard3099 & _guard3100;
wire _guard3102 = fsm_out == 1'd0;
wire _guard3103 = _guard3101 & _guard3102;
wire _guard3104 = _guard3098 | _guard3103;
wire _guard3105 = early_reset_static_par0_go_out;
wire _guard3106 = _guard3104 & _guard3105;
wire _guard3107 = fsm_out == 1'd0;
wire _guard3108 = cond_wire200_out;
wire _guard3109 = _guard3107 & _guard3108;
wire _guard3110 = fsm_out == 1'd0;
wire _guard3111 = _guard3109 & _guard3110;
wire _guard3112 = fsm_out == 1'd0;
wire _guard3113 = cond_wire202_out;
wire _guard3114 = _guard3112 & _guard3113;
wire _guard3115 = fsm_out == 1'd0;
wire _guard3116 = _guard3114 & _guard3115;
wire _guard3117 = _guard3111 | _guard3116;
wire _guard3118 = early_reset_static_par0_go_out;
wire _guard3119 = _guard3117 & _guard3118;
wire _guard3120 = fsm_out == 1'd0;
wire _guard3121 = cond_wire200_out;
wire _guard3122 = _guard3120 & _guard3121;
wire _guard3123 = fsm_out == 1'd0;
wire _guard3124 = _guard3122 & _guard3123;
wire _guard3125 = fsm_out == 1'd0;
wire _guard3126 = cond_wire202_out;
wire _guard3127 = _guard3125 & _guard3126;
wire _guard3128 = fsm_out == 1'd0;
wire _guard3129 = _guard3127 & _guard3128;
wire _guard3130 = _guard3124 | _guard3129;
wire _guard3131 = early_reset_static_par0_go_out;
wire _guard3132 = _guard3130 & _guard3131;
wire _guard3133 = cond_wire207_out;
wire _guard3134 = early_reset_static_par0_go_out;
wire _guard3135 = _guard3133 & _guard3134;
wire _guard3136 = cond_wire205_out;
wire _guard3137 = early_reset_static_par0_go_out;
wire _guard3138 = _guard3136 & _guard3137;
wire _guard3139 = fsm_out == 1'd0;
wire _guard3140 = cond_wire205_out;
wire _guard3141 = _guard3139 & _guard3140;
wire _guard3142 = fsm_out == 1'd0;
wire _guard3143 = _guard3141 & _guard3142;
wire _guard3144 = fsm_out == 1'd0;
wire _guard3145 = cond_wire207_out;
wire _guard3146 = _guard3144 & _guard3145;
wire _guard3147 = fsm_out == 1'd0;
wire _guard3148 = _guard3146 & _guard3147;
wire _guard3149 = _guard3143 | _guard3148;
wire _guard3150 = early_reset_static_par0_go_out;
wire _guard3151 = _guard3149 & _guard3150;
wire _guard3152 = fsm_out == 1'd0;
wire _guard3153 = cond_wire205_out;
wire _guard3154 = _guard3152 & _guard3153;
wire _guard3155 = fsm_out == 1'd0;
wire _guard3156 = _guard3154 & _guard3155;
wire _guard3157 = fsm_out == 1'd0;
wire _guard3158 = cond_wire207_out;
wire _guard3159 = _guard3157 & _guard3158;
wire _guard3160 = fsm_out == 1'd0;
wire _guard3161 = _guard3159 & _guard3160;
wire _guard3162 = _guard3156 | _guard3161;
wire _guard3163 = early_reset_static_par0_go_out;
wire _guard3164 = _guard3162 & _guard3163;
wire _guard3165 = fsm_out == 1'd0;
wire _guard3166 = cond_wire205_out;
wire _guard3167 = _guard3165 & _guard3166;
wire _guard3168 = fsm_out == 1'd0;
wire _guard3169 = _guard3167 & _guard3168;
wire _guard3170 = fsm_out == 1'd0;
wire _guard3171 = cond_wire207_out;
wire _guard3172 = _guard3170 & _guard3171;
wire _guard3173 = fsm_out == 1'd0;
wire _guard3174 = _guard3172 & _guard3173;
wire _guard3175 = _guard3169 | _guard3174;
wire _guard3176 = early_reset_static_par0_go_out;
wire _guard3177 = _guard3175 & _guard3176;
wire _guard3178 = cond_wire173_out;
wire _guard3179 = early_reset_static_par0_go_out;
wire _guard3180 = _guard3178 & _guard3179;
wire _guard3181 = cond_wire173_out;
wire _guard3182 = early_reset_static_par0_go_out;
wire _guard3183 = _guard3181 & _guard3182;
wire _guard3184 = cond_wire211_out;
wire _guard3185 = early_reset_static_par0_go_out;
wire _guard3186 = _guard3184 & _guard3185;
wire _guard3187 = cond_wire209_out;
wire _guard3188 = early_reset_static_par0_go_out;
wire _guard3189 = _guard3187 & _guard3188;
wire _guard3190 = fsm_out == 1'd0;
wire _guard3191 = cond_wire209_out;
wire _guard3192 = _guard3190 & _guard3191;
wire _guard3193 = fsm_out == 1'd0;
wire _guard3194 = _guard3192 & _guard3193;
wire _guard3195 = fsm_out == 1'd0;
wire _guard3196 = cond_wire211_out;
wire _guard3197 = _guard3195 & _guard3196;
wire _guard3198 = fsm_out == 1'd0;
wire _guard3199 = _guard3197 & _guard3198;
wire _guard3200 = _guard3194 | _guard3199;
wire _guard3201 = early_reset_static_par0_go_out;
wire _guard3202 = _guard3200 & _guard3201;
wire _guard3203 = fsm_out == 1'd0;
wire _guard3204 = cond_wire209_out;
wire _guard3205 = _guard3203 & _guard3204;
wire _guard3206 = fsm_out == 1'd0;
wire _guard3207 = _guard3205 & _guard3206;
wire _guard3208 = fsm_out == 1'd0;
wire _guard3209 = cond_wire211_out;
wire _guard3210 = _guard3208 & _guard3209;
wire _guard3211 = fsm_out == 1'd0;
wire _guard3212 = _guard3210 & _guard3211;
wire _guard3213 = _guard3207 | _guard3212;
wire _guard3214 = early_reset_static_par0_go_out;
wire _guard3215 = _guard3213 & _guard3214;
wire _guard3216 = fsm_out == 1'd0;
wire _guard3217 = cond_wire209_out;
wire _guard3218 = _guard3216 & _guard3217;
wire _guard3219 = fsm_out == 1'd0;
wire _guard3220 = _guard3218 & _guard3219;
wire _guard3221 = fsm_out == 1'd0;
wire _guard3222 = cond_wire211_out;
wire _guard3223 = _guard3221 & _guard3222;
wire _guard3224 = fsm_out == 1'd0;
wire _guard3225 = _guard3223 & _guard3224;
wire _guard3226 = _guard3220 | _guard3225;
wire _guard3227 = early_reset_static_par0_go_out;
wire _guard3228 = _guard3226 & _guard3227;
wire _guard3229 = cond_wire255_out;
wire _guard3230 = early_reset_static_par0_go_out;
wire _guard3231 = _guard3229 & _guard3230;
wire _guard3232 = cond_wire255_out;
wire _guard3233 = early_reset_static_par0_go_out;
wire _guard3234 = _guard3232 & _guard3233;
wire _guard3235 = early_reset_static_par0_go_out;
wire _guard3236 = early_reset_static_par0_go_out;
wire _guard3237 = fsm0_out == 5'd0;
wire _guard3238 = early_reset_static_seq_go_out;
wire _guard3239 = _guard3237 & _guard3238;
wire _guard3240 = early_reset_static_par0_go_out;
wire _guard3241 = _guard3239 | _guard3240;
wire _guard3242 = early_reset_static_par0_go_out;
wire _guard3243 = fsm0_out == 5'd0;
wire _guard3244 = early_reset_static_seq_go_out;
wire _guard3245 = _guard3243 & _guard3244;
wire _guard3246 = fsm0_out == 5'd0;
wire _guard3247 = early_reset_static_seq_go_out;
wire _guard3248 = _guard3246 & _guard3247;
wire _guard3249 = early_reset_static_par0_go_out;
wire _guard3250 = _guard3248 | _guard3249;
wire _guard3251 = fsm0_out == 5'd0;
wire _guard3252 = early_reset_static_seq_go_out;
wire _guard3253 = _guard3251 & _guard3252;
wire _guard3254 = early_reset_static_par0_go_out;
wire _guard3255 = early_reset_static_par0_go_out;
wire _guard3256 = early_reset_static_par0_go_out;
wire _guard3257 = early_reset_static_par0_go_out;
wire _guard3258 = early_reset_static_par0_go_out;
wire _guard3259 = early_reset_static_par0_go_out;
wire _guard3260 = early_reset_static_par0_go_out;
wire _guard3261 = early_reset_static_par0_go_out;
wire _guard3262 = early_reset_static_par0_go_out;
wire _guard3263 = early_reset_static_par0_go_out;
wire _guard3264 = early_reset_static_par0_go_out;
wire _guard3265 = fsm0_out == 5'd0;
wire _guard3266 = early_reset_static_seq_go_out;
wire _guard3267 = _guard3265 & _guard3266;
wire _guard3268 = early_reset_static_par0_go_out;
wire _guard3269 = _guard3267 | _guard3268;
wire _guard3270 = early_reset_static_par0_go_out;
wire _guard3271 = fsm0_out == 5'd0;
wire _guard3272 = early_reset_static_seq_go_out;
wire _guard3273 = _guard3271 & _guard3272;
wire _guard3274 = early_reset_static_par0_go_out;
wire _guard3275 = early_reset_static_par0_go_out;
wire _guard3276 = fsm0_out == 5'd0;
wire _guard3277 = early_reset_static_seq_go_out;
wire _guard3278 = _guard3276 & _guard3277;
wire _guard3279 = early_reset_static_par0_go_out;
wire _guard3280 = _guard3278 | _guard3279;
wire _guard3281 = fsm0_out == 5'd0;
wire _guard3282 = early_reset_static_seq_go_out;
wire _guard3283 = _guard3281 & _guard3282;
wire _guard3284 = early_reset_static_par0_go_out;
wire _guard3285 = ~_guard0;
wire _guard3286 = early_reset_static_par0_go_out;
wire _guard3287 = _guard3285 & _guard3286;
wire _guard3288 = early_reset_static_par0_go_out;
wire _guard3289 = early_reset_static_par0_go_out;
wire _guard3290 = early_reset_static_par0_go_out;
wire _guard3291 = early_reset_static_par0_go_out;
wire _guard3292 = ~_guard0;
wire _guard3293 = early_reset_static_par0_go_out;
wire _guard3294 = _guard3292 & _guard3293;
wire _guard3295 = early_reset_static_par0_go_out;
wire _guard3296 = early_reset_static_par0_go_out;
wire _guard3297 = early_reset_static_par0_go_out;
wire _guard3298 = early_reset_static_par0_go_out;
wire _guard3299 = early_reset_static_par0_go_out;
wire _guard3300 = early_reset_static_par0_go_out;
wire _guard3301 = early_reset_static_par0_go_out;
wire _guard3302 = ~_guard0;
wire _guard3303 = early_reset_static_par0_go_out;
wire _guard3304 = _guard3302 & _guard3303;
wire _guard3305 = early_reset_static_par0_go_out;
wire _guard3306 = ~_guard0;
wire _guard3307 = early_reset_static_par0_go_out;
wire _guard3308 = _guard3306 & _guard3307;
wire _guard3309 = early_reset_static_par0_go_out;
wire _guard3310 = early_reset_static_par0_go_out;
wire _guard3311 = early_reset_static_par0_go_out;
wire _guard3312 = early_reset_static_par0_go_out;
wire _guard3313 = early_reset_static_par0_go_out;
wire _guard3314 = early_reset_static_par0_go_out;
wire _guard3315 = early_reset_static_par0_go_out;
wire _guard3316 = ~_guard0;
wire _guard3317 = early_reset_static_par0_go_out;
wire _guard3318 = _guard3316 & _guard3317;
wire _guard3319 = ~_guard0;
wire _guard3320 = early_reset_static_par0_go_out;
wire _guard3321 = _guard3319 & _guard3320;
wire _guard3322 = early_reset_static_par0_go_out;
wire _guard3323 = early_reset_static_par0_go_out;
wire _guard3324 = ~_guard0;
wire _guard3325 = early_reset_static_par0_go_out;
wire _guard3326 = _guard3324 & _guard3325;
wire _guard3327 = early_reset_static_par0_go_out;
wire _guard3328 = ~_guard0;
wire _guard3329 = early_reset_static_par0_go_out;
wire _guard3330 = _guard3328 & _guard3329;
wire _guard3331 = early_reset_static_par0_go_out;
wire _guard3332 = early_reset_static_par0_go_out;
wire _guard3333 = early_reset_static_par0_go_out;
wire _guard3334 = early_reset_static_par0_go_out;
wire _guard3335 = early_reset_static_par0_go_out;
wire _guard3336 = early_reset_static_par0_go_out;
wire _guard3337 = early_reset_static_par0_go_out;
wire _guard3338 = early_reset_static_par0_go_out;
wire _guard3339 = early_reset_static_par0_go_out;
wire _guard3340 = early_reset_static_par0_go_out;
wire _guard3341 = early_reset_static_par0_go_out;
wire _guard3342 = ~_guard0;
wire _guard3343 = early_reset_static_par0_go_out;
wire _guard3344 = _guard3342 & _guard3343;
wire _guard3345 = early_reset_static_par0_go_out;
wire _guard3346 = ~_guard0;
wire _guard3347 = early_reset_static_par0_go_out;
wire _guard3348 = _guard3346 & _guard3347;
wire _guard3349 = early_reset_static_par0_go_out;
wire _guard3350 = early_reset_static_par0_go_out;
wire _guard3351 = ~_guard0;
wire _guard3352 = early_reset_static_par0_go_out;
wire _guard3353 = _guard3351 & _guard3352;
wire _guard3354 = early_reset_static_par0_go_out;
wire _guard3355 = early_reset_static_par0_go_out;
wire _guard3356 = early_reset_static_par0_go_out;
wire _guard3357 = early_reset_static_par0_go_out;
wire _guard3358 = early_reset_static_par0_go_out;
wire _guard3359 = early_reset_static_par0_go_out;
wire _guard3360 = early_reset_static_par0_go_out;
wire _guard3361 = early_reset_static_par0_go_out;
wire _guard3362 = ~_guard0;
wire _guard3363 = early_reset_static_par0_go_out;
wire _guard3364 = _guard3362 & _guard3363;
wire _guard3365 = early_reset_static_par0_go_out;
wire _guard3366 = ~_guard0;
wire _guard3367 = early_reset_static_par0_go_out;
wire _guard3368 = _guard3366 & _guard3367;
wire _guard3369 = ~_guard0;
wire _guard3370 = early_reset_static_par0_go_out;
wire _guard3371 = _guard3369 & _guard3370;
wire _guard3372 = early_reset_static_par0_go_out;
wire _guard3373 = ~_guard0;
wire _guard3374 = early_reset_static_par0_go_out;
wire _guard3375 = _guard3373 & _guard3374;
wire _guard3376 = early_reset_static_par0_go_out;
wire _guard3377 = early_reset_static_par0_go_out;
wire _guard3378 = early_reset_static_par0_go_out;
wire _guard3379 = early_reset_static_par0_go_out;
wire _guard3380 = ~_guard0;
wire _guard3381 = early_reset_static_par0_go_out;
wire _guard3382 = _guard3380 & _guard3381;
wire _guard3383 = cond_wire12_out;
wire _guard3384 = early_reset_static_par0_go_out;
wire _guard3385 = _guard3383 & _guard3384;
wire _guard3386 = cond_wire10_out;
wire _guard3387 = early_reset_static_par0_go_out;
wire _guard3388 = _guard3386 & _guard3387;
wire _guard3389 = fsm_out == 1'd0;
wire _guard3390 = cond_wire10_out;
wire _guard3391 = _guard3389 & _guard3390;
wire _guard3392 = fsm_out == 1'd0;
wire _guard3393 = _guard3391 & _guard3392;
wire _guard3394 = fsm_out == 1'd0;
wire _guard3395 = cond_wire12_out;
wire _guard3396 = _guard3394 & _guard3395;
wire _guard3397 = fsm_out == 1'd0;
wire _guard3398 = _guard3396 & _guard3397;
wire _guard3399 = _guard3393 | _guard3398;
wire _guard3400 = early_reset_static_par0_go_out;
wire _guard3401 = _guard3399 & _guard3400;
wire _guard3402 = fsm_out == 1'd0;
wire _guard3403 = cond_wire10_out;
wire _guard3404 = _guard3402 & _guard3403;
wire _guard3405 = fsm_out == 1'd0;
wire _guard3406 = _guard3404 & _guard3405;
wire _guard3407 = fsm_out == 1'd0;
wire _guard3408 = cond_wire12_out;
wire _guard3409 = _guard3407 & _guard3408;
wire _guard3410 = fsm_out == 1'd0;
wire _guard3411 = _guard3409 & _guard3410;
wire _guard3412 = _guard3406 | _guard3411;
wire _guard3413 = early_reset_static_par0_go_out;
wire _guard3414 = _guard3412 & _guard3413;
wire _guard3415 = fsm_out == 1'd0;
wire _guard3416 = cond_wire10_out;
wire _guard3417 = _guard3415 & _guard3416;
wire _guard3418 = fsm_out == 1'd0;
wire _guard3419 = _guard3417 & _guard3418;
wire _guard3420 = fsm_out == 1'd0;
wire _guard3421 = cond_wire12_out;
wire _guard3422 = _guard3420 & _guard3421;
wire _guard3423 = fsm_out == 1'd0;
wire _guard3424 = _guard3422 & _guard3423;
wire _guard3425 = _guard3419 | _guard3424;
wire _guard3426 = early_reset_static_par0_go_out;
wire _guard3427 = _guard3425 & _guard3426;
wire _guard3428 = cond_wire66_out;
wire _guard3429 = early_reset_static_par0_go_out;
wire _guard3430 = _guard3428 & _guard3429;
wire _guard3431 = cond_wire64_out;
wire _guard3432 = early_reset_static_par0_go_out;
wire _guard3433 = _guard3431 & _guard3432;
wire _guard3434 = fsm_out == 1'd0;
wire _guard3435 = cond_wire64_out;
wire _guard3436 = _guard3434 & _guard3435;
wire _guard3437 = fsm_out == 1'd0;
wire _guard3438 = _guard3436 & _guard3437;
wire _guard3439 = fsm_out == 1'd0;
wire _guard3440 = cond_wire66_out;
wire _guard3441 = _guard3439 & _guard3440;
wire _guard3442 = fsm_out == 1'd0;
wire _guard3443 = _guard3441 & _guard3442;
wire _guard3444 = _guard3438 | _guard3443;
wire _guard3445 = early_reset_static_par0_go_out;
wire _guard3446 = _guard3444 & _guard3445;
wire _guard3447 = fsm_out == 1'd0;
wire _guard3448 = cond_wire64_out;
wire _guard3449 = _guard3447 & _guard3448;
wire _guard3450 = fsm_out == 1'd0;
wire _guard3451 = _guard3449 & _guard3450;
wire _guard3452 = fsm_out == 1'd0;
wire _guard3453 = cond_wire66_out;
wire _guard3454 = _guard3452 & _guard3453;
wire _guard3455 = fsm_out == 1'd0;
wire _guard3456 = _guard3454 & _guard3455;
wire _guard3457 = _guard3451 | _guard3456;
wire _guard3458 = early_reset_static_par0_go_out;
wire _guard3459 = _guard3457 & _guard3458;
wire _guard3460 = fsm_out == 1'd0;
wire _guard3461 = cond_wire64_out;
wire _guard3462 = _guard3460 & _guard3461;
wire _guard3463 = fsm_out == 1'd0;
wire _guard3464 = _guard3462 & _guard3463;
wire _guard3465 = fsm_out == 1'd0;
wire _guard3466 = cond_wire66_out;
wire _guard3467 = _guard3465 & _guard3466;
wire _guard3468 = fsm_out == 1'd0;
wire _guard3469 = _guard3467 & _guard3468;
wire _guard3470 = _guard3464 | _guard3469;
wire _guard3471 = early_reset_static_par0_go_out;
wire _guard3472 = _guard3470 & _guard3471;
wire _guard3473 = cond_wire123_out;
wire _guard3474 = early_reset_static_par0_go_out;
wire _guard3475 = _guard3473 & _guard3474;
wire _guard3476 = cond_wire123_out;
wire _guard3477 = early_reset_static_par0_go_out;
wire _guard3478 = _guard3476 & _guard3477;
wire _guard3479 = cond_wire160_out;
wire _guard3480 = early_reset_static_par0_go_out;
wire _guard3481 = _guard3479 & _guard3480;
wire _guard3482 = cond_wire160_out;
wire _guard3483 = early_reset_static_par0_go_out;
wire _guard3484 = _guard3482 & _guard3483;
wire _guard3485 = cond_wire206_out;
wire _guard3486 = early_reset_static_par0_go_out;
wire _guard3487 = _guard3485 & _guard3486;
wire _guard3488 = cond_wire206_out;
wire _guard3489 = early_reset_static_par0_go_out;
wire _guard3490 = _guard3488 & _guard3489;
wire _guard3491 = cond_wire227_out;
wire _guard3492 = early_reset_static_par0_go_out;
wire _guard3493 = _guard3491 & _guard3492;
wire _guard3494 = cond_wire225_out;
wire _guard3495 = early_reset_static_par0_go_out;
wire _guard3496 = _guard3494 & _guard3495;
wire _guard3497 = fsm_out == 1'd0;
wire _guard3498 = cond_wire225_out;
wire _guard3499 = _guard3497 & _guard3498;
wire _guard3500 = fsm_out == 1'd0;
wire _guard3501 = _guard3499 & _guard3500;
wire _guard3502 = fsm_out == 1'd0;
wire _guard3503 = cond_wire227_out;
wire _guard3504 = _guard3502 & _guard3503;
wire _guard3505 = fsm_out == 1'd0;
wire _guard3506 = _guard3504 & _guard3505;
wire _guard3507 = _guard3501 | _guard3506;
wire _guard3508 = early_reset_static_par0_go_out;
wire _guard3509 = _guard3507 & _guard3508;
wire _guard3510 = fsm_out == 1'd0;
wire _guard3511 = cond_wire225_out;
wire _guard3512 = _guard3510 & _guard3511;
wire _guard3513 = fsm_out == 1'd0;
wire _guard3514 = _guard3512 & _guard3513;
wire _guard3515 = fsm_out == 1'd0;
wire _guard3516 = cond_wire227_out;
wire _guard3517 = _guard3515 & _guard3516;
wire _guard3518 = fsm_out == 1'd0;
wire _guard3519 = _guard3517 & _guard3518;
wire _guard3520 = _guard3514 | _guard3519;
wire _guard3521 = early_reset_static_par0_go_out;
wire _guard3522 = _guard3520 & _guard3521;
wire _guard3523 = fsm_out == 1'd0;
wire _guard3524 = cond_wire225_out;
wire _guard3525 = _guard3523 & _guard3524;
wire _guard3526 = fsm_out == 1'd0;
wire _guard3527 = _guard3525 & _guard3526;
wire _guard3528 = fsm_out == 1'd0;
wire _guard3529 = cond_wire227_out;
wire _guard3530 = _guard3528 & _guard3529;
wire _guard3531 = fsm_out == 1'd0;
wire _guard3532 = _guard3530 & _guard3531;
wire _guard3533 = _guard3527 | _guard3532;
wire _guard3534 = early_reset_static_par0_go_out;
wire _guard3535 = _guard3533 & _guard3534;
wire _guard3536 = cond_wire230_out;
wire _guard3537 = early_reset_static_par0_go_out;
wire _guard3538 = _guard3536 & _guard3537;
wire _guard3539 = cond_wire230_out;
wire _guard3540 = early_reset_static_par0_go_out;
wire _guard3541 = _guard3539 & _guard3540;
wire _guard3542 = cond_wire240_out;
wire _guard3543 = early_reset_static_par0_go_out;
wire _guard3544 = _guard3542 & _guard3543;
wire _guard3545 = cond_wire238_out;
wire _guard3546 = early_reset_static_par0_go_out;
wire _guard3547 = _guard3545 & _guard3546;
wire _guard3548 = fsm_out == 1'd0;
wire _guard3549 = cond_wire238_out;
wire _guard3550 = _guard3548 & _guard3549;
wire _guard3551 = fsm_out == 1'd0;
wire _guard3552 = _guard3550 & _guard3551;
wire _guard3553 = fsm_out == 1'd0;
wire _guard3554 = cond_wire240_out;
wire _guard3555 = _guard3553 & _guard3554;
wire _guard3556 = fsm_out == 1'd0;
wire _guard3557 = _guard3555 & _guard3556;
wire _guard3558 = _guard3552 | _guard3557;
wire _guard3559 = early_reset_static_par0_go_out;
wire _guard3560 = _guard3558 & _guard3559;
wire _guard3561 = fsm_out == 1'd0;
wire _guard3562 = cond_wire238_out;
wire _guard3563 = _guard3561 & _guard3562;
wire _guard3564 = fsm_out == 1'd0;
wire _guard3565 = _guard3563 & _guard3564;
wire _guard3566 = fsm_out == 1'd0;
wire _guard3567 = cond_wire240_out;
wire _guard3568 = _guard3566 & _guard3567;
wire _guard3569 = fsm_out == 1'd0;
wire _guard3570 = _guard3568 & _guard3569;
wire _guard3571 = _guard3565 | _guard3570;
wire _guard3572 = early_reset_static_par0_go_out;
wire _guard3573 = _guard3571 & _guard3572;
wire _guard3574 = fsm_out == 1'd0;
wire _guard3575 = cond_wire238_out;
wire _guard3576 = _guard3574 & _guard3575;
wire _guard3577 = fsm_out == 1'd0;
wire _guard3578 = _guard3576 & _guard3577;
wire _guard3579 = fsm_out == 1'd0;
wire _guard3580 = cond_wire240_out;
wire _guard3581 = _guard3579 & _guard3580;
wire _guard3582 = fsm_out == 1'd0;
wire _guard3583 = _guard3581 & _guard3582;
wire _guard3584 = _guard3578 | _guard3583;
wire _guard3585 = early_reset_static_par0_go_out;
wire _guard3586 = _guard3584 & _guard3585;
wire _guard3587 = cond_wire222_out;
wire _guard3588 = early_reset_static_par0_go_out;
wire _guard3589 = _guard3587 & _guard3588;
wire _guard3590 = cond_wire222_out;
wire _guard3591 = early_reset_static_par0_go_out;
wire _guard3592 = _guard3590 & _guard3591;
wire _guard3593 = fsm0_out == 5'd0;
wire _guard3594 = early_reset_static_seq_go_out;
wire _guard3595 = _guard3593 & _guard3594;
wire _guard3596 = cond_wire_out;
wire _guard3597 = early_reset_static_par0_go_out;
wire _guard3598 = _guard3596 & _guard3597;
wire _guard3599 = _guard3595 | _guard3598;
wire _guard3600 = fsm0_out == 5'd0;
wire _guard3601 = early_reset_static_seq_go_out;
wire _guard3602 = _guard3600 & _guard3601;
wire _guard3603 = cond_wire_out;
wire _guard3604 = early_reset_static_par0_go_out;
wire _guard3605 = _guard3603 & _guard3604;
wire _guard3606 = fsm0_out == 5'd0;
wire _guard3607 = early_reset_static_seq_go_out;
wire _guard3608 = _guard3606 & _guard3607;
wire _guard3609 = cond_wire19_out;
wire _guard3610 = early_reset_static_par0_go_out;
wire _guard3611 = _guard3609 & _guard3610;
wire _guard3612 = _guard3608 | _guard3611;
wire _guard3613 = fsm0_out == 5'd0;
wire _guard3614 = early_reset_static_seq_go_out;
wire _guard3615 = _guard3613 & _guard3614;
wire _guard3616 = cond_wire19_out;
wire _guard3617 = early_reset_static_par0_go_out;
wire _guard3618 = _guard3616 & _guard3617;
wire _guard3619 = fsm0_out == 5'd0;
wire _guard3620 = early_reset_static_seq_go_out;
wire _guard3621 = _guard3619 & _guard3620;
wire _guard3622 = cond_wire29_out;
wire _guard3623 = early_reset_static_par0_go_out;
wire _guard3624 = _guard3622 & _guard3623;
wire _guard3625 = _guard3621 | _guard3624;
wire _guard3626 = fsm0_out == 5'd0;
wire _guard3627 = early_reset_static_seq_go_out;
wire _guard3628 = _guard3626 & _guard3627;
wire _guard3629 = cond_wire29_out;
wire _guard3630 = early_reset_static_par0_go_out;
wire _guard3631 = _guard3629 & _guard3630;
wire _guard3632 = fsm0_out == 5'd0;
wire _guard3633 = early_reset_static_seq_go_out;
wire _guard3634 = _guard3632 & _guard3633;
wire _guard3635 = cond_wire39_out;
wire _guard3636 = early_reset_static_par0_go_out;
wire _guard3637 = _guard3635 & _guard3636;
wire _guard3638 = _guard3634 | _guard3637;
wire _guard3639 = cond_wire39_out;
wire _guard3640 = early_reset_static_par0_go_out;
wire _guard3641 = _guard3639 & _guard3640;
wire _guard3642 = fsm0_out == 5'd0;
wire _guard3643 = early_reset_static_seq_go_out;
wire _guard3644 = _guard3642 & _guard3643;
wire _guard3645 = cond_wire171_out;
wire _guard3646 = early_reset_static_par0_go_out;
wire _guard3647 = _guard3645 & _guard3646;
wire _guard3648 = cond_wire171_out;
wire _guard3649 = early_reset_static_par0_go_out;
wire _guard3650 = _guard3648 & _guard3649;
wire _guard3651 = early_reset_static_par0_go_out;
wire _guard3652 = early_reset_static_par0_go_out;
wire _guard3653 = early_reset_static_par0_go_out;
wire _guard3654 = early_reset_static_par0_go_out;
wire _guard3655 = early_reset_static_par0_go_out;
wire _guard3656 = early_reset_static_par0_go_out;
wire _guard3657 = fsm0_out == 5'd0;
wire _guard3658 = early_reset_static_seq_go_out;
wire _guard3659 = _guard3657 & _guard3658;
wire _guard3660 = early_reset_static_par0_go_out;
wire _guard3661 = _guard3659 | _guard3660;
wire _guard3662 = early_reset_static_par0_go_out;
wire _guard3663 = fsm0_out == 5'd0;
wire _guard3664 = early_reset_static_seq_go_out;
wire _guard3665 = _guard3663 & _guard3664;
wire _guard3666 = early_reset_static_par0_go_out;
wire _guard3667 = early_reset_static_par0_go_out;
wire _guard3668 = fsm0_out == 5'd0;
wire _guard3669 = early_reset_static_seq_go_out;
wire _guard3670 = _guard3668 & _guard3669;
wire _guard3671 = early_reset_static_par0_go_out;
wire _guard3672 = _guard3670 | _guard3671;
wire _guard3673 = fsm0_out == 5'd0;
wire _guard3674 = early_reset_static_seq_go_out;
wire _guard3675 = _guard3673 & _guard3674;
wire _guard3676 = early_reset_static_par0_go_out;
wire _guard3677 = early_reset_static_par0_go_out;
wire _guard3678 = early_reset_static_par0_go_out;
wire _guard3679 = early_reset_static_par0_go_out;
wire _guard3680 = early_reset_static_par0_go_out;
wire _guard3681 = early_reset_static_par0_go_out;
wire _guard3682 = early_reset_static_par0_go_out;
wire _guard3683 = early_reset_static_par0_go_out;
wire _guard3684 = early_reset_static_par0_go_out;
wire _guard3685 = early_reset_static_par0_go_out;
wire _guard3686 = early_reset_static_par0_go_out;
wire _guard3687 = early_reset_static_par0_go_out;
wire _guard3688 = early_reset_static_par0_go_out;
wire _guard3689 = early_reset_static_par0_go_out;
wire _guard3690 = early_reset_static_par0_go_out;
wire _guard3691 = early_reset_static_par0_go_out;
wire _guard3692 = early_reset_static_par0_go_out;
wire _guard3693 = early_reset_static_par0_go_out;
wire _guard3694 = early_reset_static_par0_go_out;
wire _guard3695 = early_reset_static_par0_go_out;
wire _guard3696 = early_reset_static_par0_go_out;
wire _guard3697 = early_reset_static_par0_go_out;
wire _guard3698 = early_reset_static_par0_go_out;
wire _guard3699 = early_reset_static_par0_go_out;
wire _guard3700 = early_reset_static_par0_go_out;
wire _guard3701 = early_reset_static_par0_go_out;
wire _guard3702 = early_reset_static_par0_go_out;
wire _guard3703 = early_reset_static_par0_go_out;
wire _guard3704 = ~_guard0;
wire _guard3705 = early_reset_static_par0_go_out;
wire _guard3706 = _guard3704 & _guard3705;
wire _guard3707 = early_reset_static_par0_go_out;
wire _guard3708 = early_reset_static_par0_go_out;
wire _guard3709 = early_reset_static_par0_go_out;
wire _guard3710 = early_reset_static_par0_go_out;
wire _guard3711 = early_reset_static_par0_go_out;
wire _guard3712 = early_reset_static_par0_go_out;
wire _guard3713 = ~_guard0;
wire _guard3714 = early_reset_static_par0_go_out;
wire _guard3715 = _guard3713 & _guard3714;
wire _guard3716 = early_reset_static_par0_go_out;
wire _guard3717 = early_reset_static_par0_go_out;
wire _guard3718 = early_reset_static_par0_go_out;
wire _guard3719 = early_reset_static_par0_go_out;
wire _guard3720 = early_reset_static_par0_go_out;
wire _guard3721 = early_reset_static_par0_go_out;
wire _guard3722 = early_reset_static_par0_go_out;
wire _guard3723 = early_reset_static_par0_go_out;
wire _guard3724 = early_reset_static_par0_go_out;
wire _guard3725 = early_reset_static_par0_go_out;
wire _guard3726 = ~_guard0;
wire _guard3727 = early_reset_static_par0_go_out;
wire _guard3728 = _guard3726 & _guard3727;
wire _guard3729 = early_reset_static_par0_go_out;
wire _guard3730 = ~_guard0;
wire _guard3731 = early_reset_static_par0_go_out;
wire _guard3732 = _guard3730 & _guard3731;
wire _guard3733 = ~_guard0;
wire _guard3734 = early_reset_static_par0_go_out;
wire _guard3735 = _guard3733 & _guard3734;
wire _guard3736 = early_reset_static_par0_go_out;
wire _guard3737 = ~_guard0;
wire _guard3738 = early_reset_static_par0_go_out;
wire _guard3739 = _guard3737 & _guard3738;
wire _guard3740 = early_reset_static_par0_go_out;
wire _guard3741 = early_reset_static_par0_go_out;
wire _guard3742 = ~_guard0;
wire _guard3743 = early_reset_static_par0_go_out;
wire _guard3744 = _guard3742 & _guard3743;
wire _guard3745 = early_reset_static_par0_go_out;
wire _guard3746 = ~_guard0;
wire _guard3747 = early_reset_static_par0_go_out;
wire _guard3748 = _guard3746 & _guard3747;
wire _guard3749 = early_reset_static_par0_go_out;
wire _guard3750 = ~_guard0;
wire _guard3751 = early_reset_static_par0_go_out;
wire _guard3752 = _guard3750 & _guard3751;
wire _guard3753 = early_reset_static_par0_go_out;
wire _guard3754 = early_reset_static_par0_go_out;
wire _guard3755 = ~_guard0;
wire _guard3756 = early_reset_static_par0_go_out;
wire _guard3757 = _guard3755 & _guard3756;
wire _guard3758 = early_reset_static_par0_go_out;
wire _guard3759 = early_reset_static_par0_go_out;
wire _guard3760 = early_reset_static_par0_go_out;
wire _guard3761 = early_reset_static_par0_go_out;
wire _guard3762 = early_reset_static_par0_go_out;
wire _guard3763 = early_reset_static_par0_go_out;
wire _guard3764 = early_reset_static_par0_go_out;
wire _guard3765 = early_reset_static_par0_go_out;
wire _guard3766 = early_reset_static_par0_go_out;
wire _guard3767 = early_reset_static_par0_go_out;
wire _guard3768 = early_reset_static_par0_go_out;
wire _guard3769 = early_reset_static_par0_go_out;
wire _guard3770 = early_reset_static_par0_go_out;
wire _guard3771 = early_reset_static_par0_go_out;
wire _guard3772 = early_reset_static_par0_go_out;
wire _guard3773 = early_reset_static_par0_go_out;
wire _guard3774 = ~_guard0;
wire _guard3775 = early_reset_static_par0_go_out;
wire _guard3776 = _guard3774 & _guard3775;
wire _guard3777 = early_reset_static_par0_go_out;
wire _guard3778 = ~_guard0;
wire _guard3779 = early_reset_static_par0_go_out;
wire _guard3780 = _guard3778 & _guard3779;
wire _guard3781 = ~_guard0;
wire _guard3782 = early_reset_static_par0_go_out;
wire _guard3783 = _guard3781 & _guard3782;
wire _guard3784 = early_reset_static_par0_go_out;
wire _guard3785 = early_reset_static_par0_go_out;
wire _guard3786 = early_reset_static_par0_go_out;
wire _guard3787 = early_reset_static_par0_go_out;
wire _guard3788 = ~_guard0;
wire _guard3789 = early_reset_static_par0_go_out;
wire _guard3790 = _guard3788 & _guard3789;
wire _guard3791 = cond_wire31_out;
wire _guard3792 = early_reset_static_par0_go_out;
wire _guard3793 = _guard3791 & _guard3792;
wire _guard3794 = cond_wire31_out;
wire _guard3795 = early_reset_static_par0_go_out;
wire _guard3796 = _guard3794 & _guard3795;
wire _guard3797 = cond_wire79_out;
wire _guard3798 = early_reset_static_par0_go_out;
wire _guard3799 = _guard3797 & _guard3798;
wire _guard3800 = cond_wire77_out;
wire _guard3801 = early_reset_static_par0_go_out;
wire _guard3802 = _guard3800 & _guard3801;
wire _guard3803 = fsm_out == 1'd0;
wire _guard3804 = cond_wire77_out;
wire _guard3805 = _guard3803 & _guard3804;
wire _guard3806 = fsm_out == 1'd0;
wire _guard3807 = _guard3805 & _guard3806;
wire _guard3808 = fsm_out == 1'd0;
wire _guard3809 = cond_wire79_out;
wire _guard3810 = _guard3808 & _guard3809;
wire _guard3811 = fsm_out == 1'd0;
wire _guard3812 = _guard3810 & _guard3811;
wire _guard3813 = _guard3807 | _guard3812;
wire _guard3814 = early_reset_static_par0_go_out;
wire _guard3815 = _guard3813 & _guard3814;
wire _guard3816 = fsm_out == 1'd0;
wire _guard3817 = cond_wire77_out;
wire _guard3818 = _guard3816 & _guard3817;
wire _guard3819 = fsm_out == 1'd0;
wire _guard3820 = _guard3818 & _guard3819;
wire _guard3821 = fsm_out == 1'd0;
wire _guard3822 = cond_wire79_out;
wire _guard3823 = _guard3821 & _guard3822;
wire _guard3824 = fsm_out == 1'd0;
wire _guard3825 = _guard3823 & _guard3824;
wire _guard3826 = _guard3820 | _guard3825;
wire _guard3827 = early_reset_static_par0_go_out;
wire _guard3828 = _guard3826 & _guard3827;
wire _guard3829 = fsm_out == 1'd0;
wire _guard3830 = cond_wire77_out;
wire _guard3831 = _guard3829 & _guard3830;
wire _guard3832 = fsm_out == 1'd0;
wire _guard3833 = _guard3831 & _guard3832;
wire _guard3834 = fsm_out == 1'd0;
wire _guard3835 = cond_wire79_out;
wire _guard3836 = _guard3834 & _guard3835;
wire _guard3837 = fsm_out == 1'd0;
wire _guard3838 = _guard3836 & _guard3837;
wire _guard3839 = _guard3833 | _guard3838;
wire _guard3840 = early_reset_static_par0_go_out;
wire _guard3841 = _guard3839 & _guard3840;
wire _guard3842 = cond_wire87_out;
wire _guard3843 = early_reset_static_par0_go_out;
wire _guard3844 = _guard3842 & _guard3843;
wire _guard3845 = cond_wire85_out;
wire _guard3846 = early_reset_static_par0_go_out;
wire _guard3847 = _guard3845 & _guard3846;
wire _guard3848 = fsm_out == 1'd0;
wire _guard3849 = cond_wire85_out;
wire _guard3850 = _guard3848 & _guard3849;
wire _guard3851 = fsm_out == 1'd0;
wire _guard3852 = _guard3850 & _guard3851;
wire _guard3853 = fsm_out == 1'd0;
wire _guard3854 = cond_wire87_out;
wire _guard3855 = _guard3853 & _guard3854;
wire _guard3856 = fsm_out == 1'd0;
wire _guard3857 = _guard3855 & _guard3856;
wire _guard3858 = _guard3852 | _guard3857;
wire _guard3859 = early_reset_static_par0_go_out;
wire _guard3860 = _guard3858 & _guard3859;
wire _guard3861 = fsm_out == 1'd0;
wire _guard3862 = cond_wire85_out;
wire _guard3863 = _guard3861 & _guard3862;
wire _guard3864 = fsm_out == 1'd0;
wire _guard3865 = _guard3863 & _guard3864;
wire _guard3866 = fsm_out == 1'd0;
wire _guard3867 = cond_wire87_out;
wire _guard3868 = _guard3866 & _guard3867;
wire _guard3869 = fsm_out == 1'd0;
wire _guard3870 = _guard3868 & _guard3869;
wire _guard3871 = _guard3865 | _guard3870;
wire _guard3872 = early_reset_static_par0_go_out;
wire _guard3873 = _guard3871 & _guard3872;
wire _guard3874 = fsm_out == 1'd0;
wire _guard3875 = cond_wire85_out;
wire _guard3876 = _guard3874 & _guard3875;
wire _guard3877 = fsm_out == 1'd0;
wire _guard3878 = _guard3876 & _guard3877;
wire _guard3879 = fsm_out == 1'd0;
wire _guard3880 = cond_wire87_out;
wire _guard3881 = _guard3879 & _guard3880;
wire _guard3882 = fsm_out == 1'd0;
wire _guard3883 = _guard3881 & _guard3882;
wire _guard3884 = _guard3878 | _guard3883;
wire _guard3885 = early_reset_static_par0_go_out;
wire _guard3886 = _guard3884 & _guard3885;
wire _guard3887 = cond_wire95_out;
wire _guard3888 = early_reset_static_par0_go_out;
wire _guard3889 = _guard3887 & _guard3888;
wire _guard3890 = cond_wire93_out;
wire _guard3891 = early_reset_static_par0_go_out;
wire _guard3892 = _guard3890 & _guard3891;
wire _guard3893 = fsm_out == 1'd0;
wire _guard3894 = cond_wire93_out;
wire _guard3895 = _guard3893 & _guard3894;
wire _guard3896 = fsm_out == 1'd0;
wire _guard3897 = _guard3895 & _guard3896;
wire _guard3898 = fsm_out == 1'd0;
wire _guard3899 = cond_wire95_out;
wire _guard3900 = _guard3898 & _guard3899;
wire _guard3901 = fsm_out == 1'd0;
wire _guard3902 = _guard3900 & _guard3901;
wire _guard3903 = _guard3897 | _guard3902;
wire _guard3904 = early_reset_static_par0_go_out;
wire _guard3905 = _guard3903 & _guard3904;
wire _guard3906 = fsm_out == 1'd0;
wire _guard3907 = cond_wire93_out;
wire _guard3908 = _guard3906 & _guard3907;
wire _guard3909 = fsm_out == 1'd0;
wire _guard3910 = _guard3908 & _guard3909;
wire _guard3911 = fsm_out == 1'd0;
wire _guard3912 = cond_wire95_out;
wire _guard3913 = _guard3911 & _guard3912;
wire _guard3914 = fsm_out == 1'd0;
wire _guard3915 = _guard3913 & _guard3914;
wire _guard3916 = _guard3910 | _guard3915;
wire _guard3917 = early_reset_static_par0_go_out;
wire _guard3918 = _guard3916 & _guard3917;
wire _guard3919 = fsm_out == 1'd0;
wire _guard3920 = cond_wire93_out;
wire _guard3921 = _guard3919 & _guard3920;
wire _guard3922 = fsm_out == 1'd0;
wire _guard3923 = _guard3921 & _guard3922;
wire _guard3924 = fsm_out == 1'd0;
wire _guard3925 = cond_wire95_out;
wire _guard3926 = _guard3924 & _guard3925;
wire _guard3927 = fsm_out == 1'd0;
wire _guard3928 = _guard3926 & _guard3927;
wire _guard3929 = _guard3923 | _guard3928;
wire _guard3930 = early_reset_static_par0_go_out;
wire _guard3931 = _guard3929 & _guard3930;
wire _guard3932 = cond_wire112_out;
wire _guard3933 = early_reset_static_par0_go_out;
wire _guard3934 = _guard3932 & _guard3933;
wire _guard3935 = cond_wire110_out;
wire _guard3936 = early_reset_static_par0_go_out;
wire _guard3937 = _guard3935 & _guard3936;
wire _guard3938 = fsm_out == 1'd0;
wire _guard3939 = cond_wire110_out;
wire _guard3940 = _guard3938 & _guard3939;
wire _guard3941 = fsm_out == 1'd0;
wire _guard3942 = _guard3940 & _guard3941;
wire _guard3943 = fsm_out == 1'd0;
wire _guard3944 = cond_wire112_out;
wire _guard3945 = _guard3943 & _guard3944;
wire _guard3946 = fsm_out == 1'd0;
wire _guard3947 = _guard3945 & _guard3946;
wire _guard3948 = _guard3942 | _guard3947;
wire _guard3949 = early_reset_static_par0_go_out;
wire _guard3950 = _guard3948 & _guard3949;
wire _guard3951 = fsm_out == 1'd0;
wire _guard3952 = cond_wire110_out;
wire _guard3953 = _guard3951 & _guard3952;
wire _guard3954 = fsm_out == 1'd0;
wire _guard3955 = _guard3953 & _guard3954;
wire _guard3956 = fsm_out == 1'd0;
wire _guard3957 = cond_wire112_out;
wire _guard3958 = _guard3956 & _guard3957;
wire _guard3959 = fsm_out == 1'd0;
wire _guard3960 = _guard3958 & _guard3959;
wire _guard3961 = _guard3955 | _guard3960;
wire _guard3962 = early_reset_static_par0_go_out;
wire _guard3963 = _guard3961 & _guard3962;
wire _guard3964 = fsm_out == 1'd0;
wire _guard3965 = cond_wire110_out;
wire _guard3966 = _guard3964 & _guard3965;
wire _guard3967 = fsm_out == 1'd0;
wire _guard3968 = _guard3966 & _guard3967;
wire _guard3969 = fsm_out == 1'd0;
wire _guard3970 = cond_wire112_out;
wire _guard3971 = _guard3969 & _guard3970;
wire _guard3972 = fsm_out == 1'd0;
wire _guard3973 = _guard3971 & _guard3972;
wire _guard3974 = _guard3968 | _guard3973;
wire _guard3975 = early_reset_static_par0_go_out;
wire _guard3976 = _guard3974 & _guard3975;
wire _guard3977 = cond_wire90_out;
wire _guard3978 = early_reset_static_par0_go_out;
wire _guard3979 = _guard3977 & _guard3978;
wire _guard3980 = cond_wire90_out;
wire _guard3981 = early_reset_static_par0_go_out;
wire _guard3982 = _guard3980 & _guard3981;
wire _guard3983 = cond_wire186_out;
wire _guard3984 = early_reset_static_par0_go_out;
wire _guard3985 = _guard3983 & _guard3984;
wire _guard3986 = cond_wire184_out;
wire _guard3987 = early_reset_static_par0_go_out;
wire _guard3988 = _guard3986 & _guard3987;
wire _guard3989 = fsm_out == 1'd0;
wire _guard3990 = cond_wire184_out;
wire _guard3991 = _guard3989 & _guard3990;
wire _guard3992 = fsm_out == 1'd0;
wire _guard3993 = _guard3991 & _guard3992;
wire _guard3994 = fsm_out == 1'd0;
wire _guard3995 = cond_wire186_out;
wire _guard3996 = _guard3994 & _guard3995;
wire _guard3997 = fsm_out == 1'd0;
wire _guard3998 = _guard3996 & _guard3997;
wire _guard3999 = _guard3993 | _guard3998;
wire _guard4000 = early_reset_static_par0_go_out;
wire _guard4001 = _guard3999 & _guard4000;
wire _guard4002 = fsm_out == 1'd0;
wire _guard4003 = cond_wire184_out;
wire _guard4004 = _guard4002 & _guard4003;
wire _guard4005 = fsm_out == 1'd0;
wire _guard4006 = _guard4004 & _guard4005;
wire _guard4007 = fsm_out == 1'd0;
wire _guard4008 = cond_wire186_out;
wire _guard4009 = _guard4007 & _guard4008;
wire _guard4010 = fsm_out == 1'd0;
wire _guard4011 = _guard4009 & _guard4010;
wire _guard4012 = _guard4006 | _guard4011;
wire _guard4013 = early_reset_static_par0_go_out;
wire _guard4014 = _guard4012 & _guard4013;
wire _guard4015 = fsm_out == 1'd0;
wire _guard4016 = cond_wire184_out;
wire _guard4017 = _guard4015 & _guard4016;
wire _guard4018 = fsm_out == 1'd0;
wire _guard4019 = _guard4017 & _guard4018;
wire _guard4020 = fsm_out == 1'd0;
wire _guard4021 = cond_wire186_out;
wire _guard4022 = _guard4020 & _guard4021;
wire _guard4023 = fsm_out == 1'd0;
wire _guard4024 = _guard4022 & _guard4023;
wire _guard4025 = _guard4019 | _guard4024;
wire _guard4026 = early_reset_static_par0_go_out;
wire _guard4027 = _guard4025 & _guard4026;
wire _guard4028 = cond_wire194_out;
wire _guard4029 = early_reset_static_par0_go_out;
wire _guard4030 = _guard4028 & _guard4029;
wire _guard4031 = cond_wire192_out;
wire _guard4032 = early_reset_static_par0_go_out;
wire _guard4033 = _guard4031 & _guard4032;
wire _guard4034 = fsm_out == 1'd0;
wire _guard4035 = cond_wire192_out;
wire _guard4036 = _guard4034 & _guard4035;
wire _guard4037 = fsm_out == 1'd0;
wire _guard4038 = _guard4036 & _guard4037;
wire _guard4039 = fsm_out == 1'd0;
wire _guard4040 = cond_wire194_out;
wire _guard4041 = _guard4039 & _guard4040;
wire _guard4042 = fsm_out == 1'd0;
wire _guard4043 = _guard4041 & _guard4042;
wire _guard4044 = _guard4038 | _guard4043;
wire _guard4045 = early_reset_static_par0_go_out;
wire _guard4046 = _guard4044 & _guard4045;
wire _guard4047 = fsm_out == 1'd0;
wire _guard4048 = cond_wire192_out;
wire _guard4049 = _guard4047 & _guard4048;
wire _guard4050 = fsm_out == 1'd0;
wire _guard4051 = _guard4049 & _guard4050;
wire _guard4052 = fsm_out == 1'd0;
wire _guard4053 = cond_wire194_out;
wire _guard4054 = _guard4052 & _guard4053;
wire _guard4055 = fsm_out == 1'd0;
wire _guard4056 = _guard4054 & _guard4055;
wire _guard4057 = _guard4051 | _guard4056;
wire _guard4058 = early_reset_static_par0_go_out;
wire _guard4059 = _guard4057 & _guard4058;
wire _guard4060 = fsm_out == 1'd0;
wire _guard4061 = cond_wire192_out;
wire _guard4062 = _guard4060 & _guard4061;
wire _guard4063 = fsm_out == 1'd0;
wire _guard4064 = _guard4062 & _guard4063;
wire _guard4065 = fsm_out == 1'd0;
wire _guard4066 = cond_wire194_out;
wire _guard4067 = _guard4065 & _guard4066;
wire _guard4068 = fsm_out == 1'd0;
wire _guard4069 = _guard4067 & _guard4068;
wire _guard4070 = _guard4064 | _guard4069;
wire _guard4071 = early_reset_static_par0_go_out;
wire _guard4072 = _guard4070 & _guard4071;
wire _guard4073 = cond_wire215_out;
wire _guard4074 = early_reset_static_par0_go_out;
wire _guard4075 = _guard4073 & _guard4074;
wire _guard4076 = cond_wire213_out;
wire _guard4077 = early_reset_static_par0_go_out;
wire _guard4078 = _guard4076 & _guard4077;
wire _guard4079 = fsm_out == 1'd0;
wire _guard4080 = cond_wire213_out;
wire _guard4081 = _guard4079 & _guard4080;
wire _guard4082 = fsm_out == 1'd0;
wire _guard4083 = _guard4081 & _guard4082;
wire _guard4084 = fsm_out == 1'd0;
wire _guard4085 = cond_wire215_out;
wire _guard4086 = _guard4084 & _guard4085;
wire _guard4087 = fsm_out == 1'd0;
wire _guard4088 = _guard4086 & _guard4087;
wire _guard4089 = _guard4083 | _guard4088;
wire _guard4090 = early_reset_static_par0_go_out;
wire _guard4091 = _guard4089 & _guard4090;
wire _guard4092 = fsm_out == 1'd0;
wire _guard4093 = cond_wire213_out;
wire _guard4094 = _guard4092 & _guard4093;
wire _guard4095 = fsm_out == 1'd0;
wire _guard4096 = _guard4094 & _guard4095;
wire _guard4097 = fsm_out == 1'd0;
wire _guard4098 = cond_wire215_out;
wire _guard4099 = _guard4097 & _guard4098;
wire _guard4100 = fsm_out == 1'd0;
wire _guard4101 = _guard4099 & _guard4100;
wire _guard4102 = _guard4096 | _guard4101;
wire _guard4103 = early_reset_static_par0_go_out;
wire _guard4104 = _guard4102 & _guard4103;
wire _guard4105 = fsm_out == 1'd0;
wire _guard4106 = cond_wire213_out;
wire _guard4107 = _guard4105 & _guard4106;
wire _guard4108 = fsm_out == 1'd0;
wire _guard4109 = _guard4107 & _guard4108;
wire _guard4110 = fsm_out == 1'd0;
wire _guard4111 = cond_wire215_out;
wire _guard4112 = _guard4110 & _guard4111;
wire _guard4113 = fsm_out == 1'd0;
wire _guard4114 = _guard4112 & _guard4113;
wire _guard4115 = _guard4109 | _guard4114;
wire _guard4116 = early_reset_static_par0_go_out;
wire _guard4117 = _guard4115 & _guard4116;
wire _guard4118 = cond_wire219_out;
wire _guard4119 = early_reset_static_par0_go_out;
wire _guard4120 = _guard4118 & _guard4119;
wire _guard4121 = cond_wire217_out;
wire _guard4122 = early_reset_static_par0_go_out;
wire _guard4123 = _guard4121 & _guard4122;
wire _guard4124 = fsm_out == 1'd0;
wire _guard4125 = cond_wire217_out;
wire _guard4126 = _guard4124 & _guard4125;
wire _guard4127 = fsm_out == 1'd0;
wire _guard4128 = _guard4126 & _guard4127;
wire _guard4129 = fsm_out == 1'd0;
wire _guard4130 = cond_wire219_out;
wire _guard4131 = _guard4129 & _guard4130;
wire _guard4132 = fsm_out == 1'd0;
wire _guard4133 = _guard4131 & _guard4132;
wire _guard4134 = _guard4128 | _guard4133;
wire _guard4135 = early_reset_static_par0_go_out;
wire _guard4136 = _guard4134 & _guard4135;
wire _guard4137 = fsm_out == 1'd0;
wire _guard4138 = cond_wire217_out;
wire _guard4139 = _guard4137 & _guard4138;
wire _guard4140 = fsm_out == 1'd0;
wire _guard4141 = _guard4139 & _guard4140;
wire _guard4142 = fsm_out == 1'd0;
wire _guard4143 = cond_wire219_out;
wire _guard4144 = _guard4142 & _guard4143;
wire _guard4145 = fsm_out == 1'd0;
wire _guard4146 = _guard4144 & _guard4145;
wire _guard4147 = _guard4141 | _guard4146;
wire _guard4148 = early_reset_static_par0_go_out;
wire _guard4149 = _guard4147 & _guard4148;
wire _guard4150 = fsm_out == 1'd0;
wire _guard4151 = cond_wire217_out;
wire _guard4152 = _guard4150 & _guard4151;
wire _guard4153 = fsm_out == 1'd0;
wire _guard4154 = _guard4152 & _guard4153;
wire _guard4155 = fsm_out == 1'd0;
wire _guard4156 = cond_wire219_out;
wire _guard4157 = _guard4155 & _guard4156;
wire _guard4158 = fsm_out == 1'd0;
wire _guard4159 = _guard4157 & _guard4158;
wire _guard4160 = _guard4154 | _guard4159;
wire _guard4161 = early_reset_static_par0_go_out;
wire _guard4162 = _guard4160 & _guard4161;
wire _guard4163 = cond_wire239_out;
wire _guard4164 = early_reset_static_par0_go_out;
wire _guard4165 = _guard4163 & _guard4164;
wire _guard4166 = cond_wire239_out;
wire _guard4167 = early_reset_static_par0_go_out;
wire _guard4168 = _guard4166 & _guard4167;
wire _guard4169 = cond_wire247_out;
wire _guard4170 = early_reset_static_par0_go_out;
wire _guard4171 = _guard4169 & _guard4170;
wire _guard4172 = cond_wire247_out;
wire _guard4173 = early_reset_static_par0_go_out;
wire _guard4174 = _guard4172 & _guard4173;
wire _guard4175 = cond_wire226_out;
wire _guard4176 = early_reset_static_par0_go_out;
wire _guard4177 = _guard4175 & _guard4176;
wire _guard4178 = cond_wire226_out;
wire _guard4179 = early_reset_static_par0_go_out;
wire _guard4180 = _guard4178 & _guard4179;
wire _guard4181 = cond_wire19_out;
wire _guard4182 = early_reset_static_par0_go_out;
wire _guard4183 = _guard4181 & _guard4182;
wire _guard4184 = cond_wire19_out;
wire _guard4185 = early_reset_static_par0_go_out;
wire _guard4186 = _guard4184 & _guard4185;
wire _guard4187 = fsm0_out == 5'd0;
wire _guard4188 = early_reset_static_seq_go_out;
wire _guard4189 = _guard4187 & _guard4188;
wire _guard4190 = cond_wire24_out;
wire _guard4191 = early_reset_static_par0_go_out;
wire _guard4192 = _guard4190 & _guard4191;
wire _guard4193 = _guard4189 | _guard4192;
wire _guard4194 = fsm0_out == 5'd0;
wire _guard4195 = early_reset_static_seq_go_out;
wire _guard4196 = _guard4194 & _guard4195;
wire _guard4197 = cond_wire24_out;
wire _guard4198 = early_reset_static_par0_go_out;
wire _guard4199 = _guard4197 & _guard4198;
wire _guard4200 = cond_wire29_out;
wire _guard4201 = early_reset_static_par0_go_out;
wire _guard4202 = _guard4200 & _guard4201;
wire _guard4203 = cond_wire29_out;
wire _guard4204 = early_reset_static_par0_go_out;
wire _guard4205 = _guard4203 & _guard4204;
wire _guard4206 = early_reset_static_par0_go_out;
wire _guard4207 = early_reset_static_par0_go_out;
wire _guard4208 = early_reset_static_par0_go_out;
wire _guard4209 = early_reset_static_par0_go_out;
wire _guard4210 = fsm0_out == 5'd0;
wire _guard4211 = early_reset_static_seq_go_out;
wire _guard4212 = _guard4210 & _guard4211;
wire _guard4213 = early_reset_static_par0_go_out;
wire _guard4214 = _guard4212 | _guard4213;
wire _guard4215 = fsm0_out == 5'd0;
wire _guard4216 = early_reset_static_seq_go_out;
wire _guard4217 = _guard4215 & _guard4216;
wire _guard4218 = early_reset_static_par0_go_out;
wire _guard4219 = early_reset_static_par0_go_out;
wire _guard4220 = early_reset_static_par0_go_out;
wire _guard4221 = fsm0_out == 5'd0;
wire _guard4222 = early_reset_static_seq_go_out;
wire _guard4223 = _guard4221 & _guard4222;
wire _guard4224 = early_reset_static_par0_go_out;
wire _guard4225 = _guard4223 | _guard4224;
wire _guard4226 = early_reset_static_par0_go_out;
wire _guard4227 = fsm0_out == 5'd0;
wire _guard4228 = early_reset_static_seq_go_out;
wire _guard4229 = _guard4227 & _guard4228;
wire _guard4230 = early_reset_static_par0_go_out;
wire _guard4231 = early_reset_static_par0_go_out;
wire _guard4232 = fsm0_out == 5'd0;
wire _guard4233 = early_reset_static_seq_go_out;
wire _guard4234 = _guard4232 & _guard4233;
wire _guard4235 = early_reset_static_par0_go_out;
wire _guard4236 = _guard4234 | _guard4235;
wire _guard4237 = fsm0_out == 5'd0;
wire _guard4238 = early_reset_static_seq_go_out;
wire _guard4239 = _guard4237 & _guard4238;
wire _guard4240 = early_reset_static_par0_go_out;
wire _guard4241 = early_reset_static_par0_go_out;
wire _guard4242 = early_reset_static_par0_go_out;
wire _guard4243 = ~_guard0;
wire _guard4244 = early_reset_static_par0_go_out;
wire _guard4245 = _guard4243 & _guard4244;
wire _guard4246 = early_reset_static_par0_go_out;
wire _guard4247 = early_reset_static_par0_go_out;
wire _guard4248 = early_reset_static_par0_go_out;
wire _guard4249 = early_reset_static_par0_go_out;
wire _guard4250 = early_reset_static_par0_go_out;
wire _guard4251 = early_reset_static_par0_go_out;
wire _guard4252 = ~_guard0;
wire _guard4253 = early_reset_static_par0_go_out;
wire _guard4254 = _guard4252 & _guard4253;
wire _guard4255 = early_reset_static_par0_go_out;
wire _guard4256 = early_reset_static_par0_go_out;
wire _guard4257 = early_reset_static_par0_go_out;
wire _guard4258 = early_reset_static_par0_go_out;
wire _guard4259 = early_reset_static_par0_go_out;
wire _guard4260 = early_reset_static_par0_go_out;
wire _guard4261 = early_reset_static_par0_go_out;
wire _guard4262 = early_reset_static_par0_go_out;
wire _guard4263 = early_reset_static_par0_go_out;
wire _guard4264 = early_reset_static_par0_go_out;
wire _guard4265 = early_reset_static_par0_go_out;
wire _guard4266 = early_reset_static_par0_go_out;
wire _guard4267 = ~_guard0;
wire _guard4268 = early_reset_static_par0_go_out;
wire _guard4269 = _guard4267 & _guard4268;
wire _guard4270 = early_reset_static_par0_go_out;
wire _guard4271 = early_reset_static_par0_go_out;
wire _guard4272 = ~_guard0;
wire _guard4273 = early_reset_static_par0_go_out;
wire _guard4274 = _guard4272 & _guard4273;
wire _guard4275 = early_reset_static_par0_go_out;
wire _guard4276 = ~_guard0;
wire _guard4277 = early_reset_static_par0_go_out;
wire _guard4278 = _guard4276 & _guard4277;
wire _guard4279 = early_reset_static_par0_go_out;
wire _guard4280 = early_reset_static_par0_go_out;
wire _guard4281 = early_reset_static_par0_go_out;
wire _guard4282 = early_reset_static_par0_go_out;
wire _guard4283 = early_reset_static_par0_go_out;
wire _guard4284 = early_reset_static_par0_go_out;
wire _guard4285 = early_reset_static_par0_go_out;
wire _guard4286 = ~_guard0;
wire _guard4287 = early_reset_static_par0_go_out;
wire _guard4288 = _guard4286 & _guard4287;
wire _guard4289 = early_reset_static_par0_go_out;
wire _guard4290 = early_reset_static_par0_go_out;
wire _guard4291 = early_reset_static_par0_go_out;
wire _guard4292 = early_reset_static_par0_go_out;
wire _guard4293 = early_reset_static_par0_go_out;
wire _guard4294 = ~_guard0;
wire _guard4295 = early_reset_static_par0_go_out;
wire _guard4296 = _guard4294 & _guard4295;
wire _guard4297 = early_reset_static_par0_go_out;
wire _guard4298 = early_reset_static_par0_go_out;
wire _guard4299 = ~_guard0;
wire _guard4300 = early_reset_static_par0_go_out;
wire _guard4301 = _guard4299 & _guard4300;
wire _guard4302 = early_reset_static_par0_go_out;
wire _guard4303 = early_reset_static_par0_go_out;
wire _guard4304 = early_reset_static_par0_go_out;
wire _guard4305 = early_reset_static_par0_go_out;
wire _guard4306 = early_reset_static_par0_go_out;
wire _guard4307 = early_reset_static_par0_go_out;
wire _guard4308 = ~_guard0;
wire _guard4309 = early_reset_static_par0_go_out;
wire _guard4310 = _guard4308 & _guard4309;
wire _guard4311 = early_reset_static_par0_go_out;
wire _guard4312 = early_reset_static_par0_go_out;
wire _guard4313 = early_reset_static_par0_go_out;
wire _guard4314 = early_reset_static_par0_go_out;
wire _guard4315 = early_reset_static_seq_go_out;
wire _guard4316 = fsm0_out != 5'd28;
wire _guard4317 = early_reset_static_seq_go_out;
wire _guard4318 = _guard4316 & _guard4317;
wire _guard4319 = fsm0_out == 5'd28;
wire _guard4320 = early_reset_static_seq_go_out;
wire _guard4321 = _guard4319 & _guard4320;
wire _guard4322 = cond_wire62_out;
wire _guard4323 = early_reset_static_par0_go_out;
wire _guard4324 = _guard4322 & _guard4323;
wire _guard4325 = cond_wire60_out;
wire _guard4326 = early_reset_static_par0_go_out;
wire _guard4327 = _guard4325 & _guard4326;
wire _guard4328 = fsm_out == 1'd0;
wire _guard4329 = cond_wire60_out;
wire _guard4330 = _guard4328 & _guard4329;
wire _guard4331 = fsm_out == 1'd0;
wire _guard4332 = _guard4330 & _guard4331;
wire _guard4333 = fsm_out == 1'd0;
wire _guard4334 = cond_wire62_out;
wire _guard4335 = _guard4333 & _guard4334;
wire _guard4336 = fsm_out == 1'd0;
wire _guard4337 = _guard4335 & _guard4336;
wire _guard4338 = _guard4332 | _guard4337;
wire _guard4339 = early_reset_static_par0_go_out;
wire _guard4340 = _guard4338 & _guard4339;
wire _guard4341 = fsm_out == 1'd0;
wire _guard4342 = cond_wire60_out;
wire _guard4343 = _guard4341 & _guard4342;
wire _guard4344 = fsm_out == 1'd0;
wire _guard4345 = _guard4343 & _guard4344;
wire _guard4346 = fsm_out == 1'd0;
wire _guard4347 = cond_wire62_out;
wire _guard4348 = _guard4346 & _guard4347;
wire _guard4349 = fsm_out == 1'd0;
wire _guard4350 = _guard4348 & _guard4349;
wire _guard4351 = _guard4345 | _guard4350;
wire _guard4352 = early_reset_static_par0_go_out;
wire _guard4353 = _guard4351 & _guard4352;
wire _guard4354 = fsm_out == 1'd0;
wire _guard4355 = cond_wire60_out;
wire _guard4356 = _guard4354 & _guard4355;
wire _guard4357 = fsm_out == 1'd0;
wire _guard4358 = _guard4356 & _guard4357;
wire _guard4359 = fsm_out == 1'd0;
wire _guard4360 = cond_wire62_out;
wire _guard4361 = _guard4359 & _guard4360;
wire _guard4362 = fsm_out == 1'd0;
wire _guard4363 = _guard4361 & _guard4362;
wire _guard4364 = _guard4358 | _guard4363;
wire _guard4365 = early_reset_static_par0_go_out;
wire _guard4366 = _guard4364 & _guard4365;
wire _guard4367 = cond_wire31_out;
wire _guard4368 = early_reset_static_par0_go_out;
wire _guard4369 = _guard4367 & _guard4368;
wire _guard4370 = cond_wire31_out;
wire _guard4371 = early_reset_static_par0_go_out;
wire _guard4372 = _guard4370 & _guard4371;
wire _guard4373 = cond_wire41_out;
wire _guard4374 = early_reset_static_par0_go_out;
wire _guard4375 = _guard4373 & _guard4374;
wire _guard4376 = cond_wire41_out;
wire _guard4377 = early_reset_static_par0_go_out;
wire _guard4378 = _guard4376 & _guard4377;
wire _guard4379 = cond_wire74_out;
wire _guard4380 = early_reset_static_par0_go_out;
wire _guard4381 = _guard4379 & _guard4380;
wire _guard4382 = cond_wire74_out;
wire _guard4383 = early_reset_static_par0_go_out;
wire _guard4384 = _guard4382 & _guard4383;
wire _guard4385 = cond_wire78_out;
wire _guard4386 = early_reset_static_par0_go_out;
wire _guard4387 = _guard4385 & _guard4386;
wire _guard4388 = cond_wire78_out;
wire _guard4389 = early_reset_static_par0_go_out;
wire _guard4390 = _guard4388 & _guard4389;
wire _guard4391 = cond_wire165_out;
wire _guard4392 = early_reset_static_par0_go_out;
wire _guard4393 = _guard4391 & _guard4392;
wire _guard4394 = cond_wire163_out;
wire _guard4395 = early_reset_static_par0_go_out;
wire _guard4396 = _guard4394 & _guard4395;
wire _guard4397 = fsm_out == 1'd0;
wire _guard4398 = cond_wire163_out;
wire _guard4399 = _guard4397 & _guard4398;
wire _guard4400 = fsm_out == 1'd0;
wire _guard4401 = _guard4399 & _guard4400;
wire _guard4402 = fsm_out == 1'd0;
wire _guard4403 = cond_wire165_out;
wire _guard4404 = _guard4402 & _guard4403;
wire _guard4405 = fsm_out == 1'd0;
wire _guard4406 = _guard4404 & _guard4405;
wire _guard4407 = _guard4401 | _guard4406;
wire _guard4408 = early_reset_static_par0_go_out;
wire _guard4409 = _guard4407 & _guard4408;
wire _guard4410 = fsm_out == 1'd0;
wire _guard4411 = cond_wire163_out;
wire _guard4412 = _guard4410 & _guard4411;
wire _guard4413 = fsm_out == 1'd0;
wire _guard4414 = _guard4412 & _guard4413;
wire _guard4415 = fsm_out == 1'd0;
wire _guard4416 = cond_wire165_out;
wire _guard4417 = _guard4415 & _guard4416;
wire _guard4418 = fsm_out == 1'd0;
wire _guard4419 = _guard4417 & _guard4418;
wire _guard4420 = _guard4414 | _guard4419;
wire _guard4421 = early_reset_static_par0_go_out;
wire _guard4422 = _guard4420 & _guard4421;
wire _guard4423 = fsm_out == 1'd0;
wire _guard4424 = cond_wire163_out;
wire _guard4425 = _guard4423 & _guard4424;
wire _guard4426 = fsm_out == 1'd0;
wire _guard4427 = _guard4425 & _guard4426;
wire _guard4428 = fsm_out == 1'd0;
wire _guard4429 = cond_wire165_out;
wire _guard4430 = _guard4428 & _guard4429;
wire _guard4431 = fsm_out == 1'd0;
wire _guard4432 = _guard4430 & _guard4431;
wire _guard4433 = _guard4427 | _guard4432;
wire _guard4434 = early_reset_static_par0_go_out;
wire _guard4435 = _guard4433 & _guard4434;
wire _guard4436 = cond_wire148_out;
wire _guard4437 = early_reset_static_par0_go_out;
wire _guard4438 = _guard4436 & _guard4437;
wire _guard4439 = cond_wire148_out;
wire _guard4440 = early_reset_static_par0_go_out;
wire _guard4441 = _guard4439 & _guard4440;
wire _guard4442 = cond_wire156_out;
wire _guard4443 = early_reset_static_par0_go_out;
wire _guard4444 = _guard4442 & _guard4443;
wire _guard4445 = cond_wire156_out;
wire _guard4446 = early_reset_static_par0_go_out;
wire _guard4447 = _guard4445 & _guard4446;
wire _guard4448 = cond_wire263_out;
wire _guard4449 = early_reset_static_par0_go_out;
wire _guard4450 = _guard4448 & _guard4449;
wire _guard4451 = cond_wire263_out;
wire _guard4452 = early_reset_static_par0_go_out;
wire _guard4453 = _guard4451 & _guard4452;
wire _guard4454 = cond_wire34_out;
wire _guard4455 = early_reset_static_par0_go_out;
wire _guard4456 = _guard4454 & _guard4455;
wire _guard4457 = cond_wire34_out;
wire _guard4458 = early_reset_static_par0_go_out;
wire _guard4459 = _guard4457 & _guard4458;
wire _guard4460 = fsm0_out == 5'd0;
wire _guard4461 = early_reset_static_seq_go_out;
wire _guard4462 = _guard4460 & _guard4461;
wire _guard4463 = cond_wire138_out;
wire _guard4464 = early_reset_static_par0_go_out;
wire _guard4465 = _guard4463 & _guard4464;
wire _guard4466 = _guard4462 | _guard4465;
wire _guard4467 = fsm0_out == 5'd0;
wire _guard4468 = early_reset_static_seq_go_out;
wire _guard4469 = _guard4467 & _guard4468;
wire _guard4470 = cond_wire138_out;
wire _guard4471 = early_reset_static_par0_go_out;
wire _guard4472 = _guard4470 & _guard4471;
wire _guard4473 = fsm0_out == 5'd0;
wire _guard4474 = early_reset_static_seq_go_out;
wire _guard4475 = _guard4473 & _guard4474;
wire _guard4476 = early_reset_static_par0_go_out;
wire _guard4477 = _guard4475 | _guard4476;
wire _guard4478 = fsm0_out == 5'd0;
wire _guard4479 = early_reset_static_seq_go_out;
wire _guard4480 = _guard4478 & _guard4479;
wire _guard4481 = early_reset_static_par0_go_out;
wire _guard4482 = early_reset_static_par0_go_out;
wire _guard4483 = early_reset_static_par0_go_out;
wire _guard4484 = early_reset_static_par0_go_out;
wire _guard4485 = early_reset_static_par0_go_out;
wire _guard4486 = fsm0_out == 5'd0;
wire _guard4487 = early_reset_static_seq_go_out;
wire _guard4488 = _guard4486 & _guard4487;
wire _guard4489 = early_reset_static_par0_go_out;
wire _guard4490 = _guard4488 | _guard4489;
wire _guard4491 = fsm0_out == 5'd0;
wire _guard4492 = early_reset_static_seq_go_out;
wire _guard4493 = _guard4491 & _guard4492;
wire _guard4494 = early_reset_static_par0_go_out;
wire _guard4495 = fsm0_out == 5'd0;
wire _guard4496 = early_reset_static_seq_go_out;
wire _guard4497 = _guard4495 & _guard4496;
wire _guard4498 = early_reset_static_par0_go_out;
wire _guard4499 = _guard4497 | _guard4498;
wire _guard4500 = early_reset_static_par0_go_out;
wire _guard4501 = fsm0_out == 5'd0;
wire _guard4502 = early_reset_static_seq_go_out;
wire _guard4503 = _guard4501 & _guard4502;
wire _guard4504 = early_reset_static_par0_go_out;
wire _guard4505 = early_reset_static_par0_go_out;
wire _guard4506 = early_reset_static_par0_go_out;
wire _guard4507 = early_reset_static_par0_go_out;
wire _guard4508 = early_reset_static_par0_go_out;
wire _guard4509 = ~_guard0;
wire _guard4510 = early_reset_static_par0_go_out;
wire _guard4511 = _guard4509 & _guard4510;
wire _guard4512 = early_reset_static_par0_go_out;
wire _guard4513 = early_reset_static_par0_go_out;
wire _guard4514 = early_reset_static_par0_go_out;
wire _guard4515 = early_reset_static_par0_go_out;
wire _guard4516 = early_reset_static_par0_go_out;
wire _guard4517 = ~_guard0;
wire _guard4518 = early_reset_static_par0_go_out;
wire _guard4519 = _guard4517 & _guard4518;
wire _guard4520 = early_reset_static_par0_go_out;
wire _guard4521 = early_reset_static_par0_go_out;
wire _guard4522 = early_reset_static_par0_go_out;
wire _guard4523 = early_reset_static_par0_go_out;
wire _guard4524 = ~_guard0;
wire _guard4525 = early_reset_static_par0_go_out;
wire _guard4526 = _guard4524 & _guard4525;
wire _guard4527 = early_reset_static_par0_go_out;
wire _guard4528 = early_reset_static_par0_go_out;
wire _guard4529 = early_reset_static_par0_go_out;
wire _guard4530 = early_reset_static_par0_go_out;
wire _guard4531 = ~_guard0;
wire _guard4532 = early_reset_static_par0_go_out;
wire _guard4533 = _guard4531 & _guard4532;
wire _guard4534 = early_reset_static_par0_go_out;
wire _guard4535 = ~_guard0;
wire _guard4536 = early_reset_static_par0_go_out;
wire _guard4537 = _guard4535 & _guard4536;
wire _guard4538 = ~_guard0;
wire _guard4539 = early_reset_static_par0_go_out;
wire _guard4540 = _guard4538 & _guard4539;
wire _guard4541 = early_reset_static_par0_go_out;
wire _guard4542 = early_reset_static_par0_go_out;
wire _guard4543 = ~_guard0;
wire _guard4544 = early_reset_static_par0_go_out;
wire _guard4545 = _guard4543 & _guard4544;
wire _guard4546 = early_reset_static_par0_go_out;
wire _guard4547 = early_reset_static_par0_go_out;
wire _guard4548 = early_reset_static_par0_go_out;
wire _guard4549 = ~_guard0;
wire _guard4550 = early_reset_static_par0_go_out;
wire _guard4551 = _guard4549 & _guard4550;
wire _guard4552 = early_reset_static_par0_go_out;
wire _guard4553 = ~_guard0;
wire _guard4554 = early_reset_static_par0_go_out;
wire _guard4555 = _guard4553 & _guard4554;
wire _guard4556 = early_reset_static_par0_go_out;
wire _guard4557 = early_reset_static_par0_go_out;
wire _guard4558 = ~_guard0;
wire _guard4559 = early_reset_static_par0_go_out;
wire _guard4560 = _guard4558 & _guard4559;
wire _guard4561 = early_reset_static_par0_go_out;
wire _guard4562 = early_reset_static_par0_go_out;
wire _guard4563 = early_reset_static_par0_go_out;
wire _guard4564 = early_reset_static_par0_go_out;
wire _guard4565 = ~_guard0;
wire _guard4566 = early_reset_static_par0_go_out;
wire _guard4567 = _guard4565 & _guard4566;
wire _guard4568 = early_reset_static_par0_go_out;
wire _guard4569 = ~_guard0;
wire _guard4570 = early_reset_static_par0_go_out;
wire _guard4571 = _guard4569 & _guard4570;
wire _guard4572 = early_reset_static_par0_go_out;
wire _guard4573 = ~_guard0;
wire _guard4574 = early_reset_static_par0_go_out;
wire _guard4575 = _guard4573 & _guard4574;
wire _guard4576 = ~_guard0;
wire _guard4577 = early_reset_static_par0_go_out;
wire _guard4578 = _guard4576 & _guard4577;
wire _guard4579 = early_reset_static_par0_go_out;
wire _guard4580 = early_reset_static_par0_go_out;
wire _guard4581 = early_reset_static_par0_go_out;
wire _guard4582 = early_reset_static_par0_go_out;
wire _guard4583 = early_reset_static_par0_go_out;
wire _guard4584 = early_reset_static_par0_go_out;
wire _guard4585 = early_reset_static_par0_go_out;
wire _guard4586 = early_reset_static_par0_go_out;
wire _guard4587 = ~_guard0;
wire _guard4588 = early_reset_static_par0_go_out;
wire _guard4589 = _guard4587 & _guard4588;
wire _guard4590 = ~_guard0;
wire _guard4591 = early_reset_static_par0_go_out;
wire _guard4592 = _guard4590 & _guard4591;
wire _guard4593 = early_reset_static_par0_go_out;
wire _guard4594 = early_reset_static_par0_go_out;
wire _guard4595 = early_reset_static_par0_go_out;
wire _guard4596 = early_reset_static_par0_go_out;
wire _guard4597 = early_reset_static_par0_go_out;
wire _guard4598 = early_reset_static_par0_go_out;
wire _guard4599 = early_reset_static_par0_go_out;
wire _guard4600 = early_reset_static_par0_go_out;
wire _guard4601 = ~_guard0;
wire _guard4602 = early_reset_static_par0_go_out;
wire _guard4603 = _guard4601 & _guard4602;
wire _guard4604 = early_reset_static_par0_go_out;
wire _guard4605 = ~_guard0;
wire _guard4606 = early_reset_static_par0_go_out;
wire _guard4607 = _guard4605 & _guard4606;
wire _guard4608 = early_reset_static_par0_go_out;
wire _guard4609 = early_reset_static_par0_go_out;
wire _guard4610 = early_reset_static_par0_go_out;
wire _guard4611 = early_reset_static_par0_go_out;
wire _guard4612 = early_reset_static_par0_go_out;
wire _guard4613 = early_reset_static_par0_go_out;
wire _guard4614 = early_reset_static_par0_go_out;
wire _guard4615 = early_reset_static_par0_go_out;
wire _guard4616 = fsm0_out == 5'd0;
wire _guard4617 = signal_reg_out;
wire _guard4618 = _guard4616 & _guard4617;
wire _guard4619 = cond_wire4_out;
wire _guard4620 = early_reset_static_par0_go_out;
wire _guard4621 = _guard4619 & _guard4620;
wire _guard4622 = cond_wire4_out;
wire _guard4623 = early_reset_static_par0_go_out;
wire _guard4624 = _guard4622 & _guard4623;
wire _guard4625 = cond_wire6_out;
wire _guard4626 = early_reset_static_par0_go_out;
wire _guard4627 = _guard4625 & _guard4626;
wire _guard4628 = cond_wire6_out;
wire _guard4629 = early_reset_static_par0_go_out;
wire _guard4630 = _guard4628 & _guard4629;
wire _guard4631 = cond_wire22_out;
wire _guard4632 = early_reset_static_par0_go_out;
wire _guard4633 = _guard4631 & _guard4632;
wire _guard4634 = cond_wire20_out;
wire _guard4635 = early_reset_static_par0_go_out;
wire _guard4636 = _guard4634 & _guard4635;
wire _guard4637 = fsm_out == 1'd0;
wire _guard4638 = cond_wire20_out;
wire _guard4639 = _guard4637 & _guard4638;
wire _guard4640 = fsm_out == 1'd0;
wire _guard4641 = _guard4639 & _guard4640;
wire _guard4642 = fsm_out == 1'd0;
wire _guard4643 = cond_wire22_out;
wire _guard4644 = _guard4642 & _guard4643;
wire _guard4645 = fsm_out == 1'd0;
wire _guard4646 = _guard4644 & _guard4645;
wire _guard4647 = _guard4641 | _guard4646;
wire _guard4648 = early_reset_static_par0_go_out;
wire _guard4649 = _guard4647 & _guard4648;
wire _guard4650 = fsm_out == 1'd0;
wire _guard4651 = cond_wire20_out;
wire _guard4652 = _guard4650 & _guard4651;
wire _guard4653 = fsm_out == 1'd0;
wire _guard4654 = _guard4652 & _guard4653;
wire _guard4655 = fsm_out == 1'd0;
wire _guard4656 = cond_wire22_out;
wire _guard4657 = _guard4655 & _guard4656;
wire _guard4658 = fsm_out == 1'd0;
wire _guard4659 = _guard4657 & _guard4658;
wire _guard4660 = _guard4654 | _guard4659;
wire _guard4661 = early_reset_static_par0_go_out;
wire _guard4662 = _guard4660 & _guard4661;
wire _guard4663 = fsm_out == 1'd0;
wire _guard4664 = cond_wire20_out;
wire _guard4665 = _guard4663 & _guard4664;
wire _guard4666 = fsm_out == 1'd0;
wire _guard4667 = _guard4665 & _guard4666;
wire _guard4668 = fsm_out == 1'd0;
wire _guard4669 = cond_wire22_out;
wire _guard4670 = _guard4668 & _guard4669;
wire _guard4671 = fsm_out == 1'd0;
wire _guard4672 = _guard4670 & _guard4671;
wire _guard4673 = _guard4667 | _guard4672;
wire _guard4674 = early_reset_static_par0_go_out;
wire _guard4675 = _guard4673 & _guard4674;
wire _guard4676 = cond_wire53_out;
wire _guard4677 = early_reset_static_par0_go_out;
wire _guard4678 = _guard4676 & _guard4677;
wire _guard4679 = cond_wire53_out;
wire _guard4680 = early_reset_static_par0_go_out;
wire _guard4681 = _guard4679 & _guard4680;
wire _guard4682 = cond_wire99_out;
wire _guard4683 = early_reset_static_par0_go_out;
wire _guard4684 = _guard4682 & _guard4683;
wire _guard4685 = cond_wire97_out;
wire _guard4686 = early_reset_static_par0_go_out;
wire _guard4687 = _guard4685 & _guard4686;
wire _guard4688 = fsm_out == 1'd0;
wire _guard4689 = cond_wire97_out;
wire _guard4690 = _guard4688 & _guard4689;
wire _guard4691 = fsm_out == 1'd0;
wire _guard4692 = _guard4690 & _guard4691;
wire _guard4693 = fsm_out == 1'd0;
wire _guard4694 = cond_wire99_out;
wire _guard4695 = _guard4693 & _guard4694;
wire _guard4696 = fsm_out == 1'd0;
wire _guard4697 = _guard4695 & _guard4696;
wire _guard4698 = _guard4692 | _guard4697;
wire _guard4699 = early_reset_static_par0_go_out;
wire _guard4700 = _guard4698 & _guard4699;
wire _guard4701 = fsm_out == 1'd0;
wire _guard4702 = cond_wire97_out;
wire _guard4703 = _guard4701 & _guard4702;
wire _guard4704 = fsm_out == 1'd0;
wire _guard4705 = _guard4703 & _guard4704;
wire _guard4706 = fsm_out == 1'd0;
wire _guard4707 = cond_wire99_out;
wire _guard4708 = _guard4706 & _guard4707;
wire _guard4709 = fsm_out == 1'd0;
wire _guard4710 = _guard4708 & _guard4709;
wire _guard4711 = _guard4705 | _guard4710;
wire _guard4712 = early_reset_static_par0_go_out;
wire _guard4713 = _guard4711 & _guard4712;
wire _guard4714 = fsm_out == 1'd0;
wire _guard4715 = cond_wire97_out;
wire _guard4716 = _guard4714 & _guard4715;
wire _guard4717 = fsm_out == 1'd0;
wire _guard4718 = _guard4716 & _guard4717;
wire _guard4719 = fsm_out == 1'd0;
wire _guard4720 = cond_wire99_out;
wire _guard4721 = _guard4719 & _guard4720;
wire _guard4722 = fsm_out == 1'd0;
wire _guard4723 = _guard4721 & _guard4722;
wire _guard4724 = _guard4718 | _guard4723;
wire _guard4725 = early_reset_static_par0_go_out;
wire _guard4726 = _guard4724 & _guard4725;
wire _guard4727 = cond_wire105_out;
wire _guard4728 = early_reset_static_par0_go_out;
wire _guard4729 = _guard4727 & _guard4728;
wire _guard4730 = cond_wire105_out;
wire _guard4731 = early_reset_static_par0_go_out;
wire _guard4732 = _guard4730 & _guard4731;
wire _guard4733 = cond_wire149_out;
wire _guard4734 = early_reset_static_par0_go_out;
wire _guard4735 = _guard4733 & _guard4734;
wire _guard4736 = cond_wire147_out;
wire _guard4737 = early_reset_static_par0_go_out;
wire _guard4738 = _guard4736 & _guard4737;
wire _guard4739 = fsm_out == 1'd0;
wire _guard4740 = cond_wire147_out;
wire _guard4741 = _guard4739 & _guard4740;
wire _guard4742 = fsm_out == 1'd0;
wire _guard4743 = _guard4741 & _guard4742;
wire _guard4744 = fsm_out == 1'd0;
wire _guard4745 = cond_wire149_out;
wire _guard4746 = _guard4744 & _guard4745;
wire _guard4747 = fsm_out == 1'd0;
wire _guard4748 = _guard4746 & _guard4747;
wire _guard4749 = _guard4743 | _guard4748;
wire _guard4750 = early_reset_static_par0_go_out;
wire _guard4751 = _guard4749 & _guard4750;
wire _guard4752 = fsm_out == 1'd0;
wire _guard4753 = cond_wire147_out;
wire _guard4754 = _guard4752 & _guard4753;
wire _guard4755 = fsm_out == 1'd0;
wire _guard4756 = _guard4754 & _guard4755;
wire _guard4757 = fsm_out == 1'd0;
wire _guard4758 = cond_wire149_out;
wire _guard4759 = _guard4757 & _guard4758;
wire _guard4760 = fsm_out == 1'd0;
wire _guard4761 = _guard4759 & _guard4760;
wire _guard4762 = _guard4756 | _guard4761;
wire _guard4763 = early_reset_static_par0_go_out;
wire _guard4764 = _guard4762 & _guard4763;
wire _guard4765 = fsm_out == 1'd0;
wire _guard4766 = cond_wire147_out;
wire _guard4767 = _guard4765 & _guard4766;
wire _guard4768 = fsm_out == 1'd0;
wire _guard4769 = _guard4767 & _guard4768;
wire _guard4770 = fsm_out == 1'd0;
wire _guard4771 = cond_wire149_out;
wire _guard4772 = _guard4770 & _guard4771;
wire _guard4773 = fsm_out == 1'd0;
wire _guard4774 = _guard4772 & _guard4773;
wire _guard4775 = _guard4769 | _guard4774;
wire _guard4776 = early_reset_static_par0_go_out;
wire _guard4777 = _guard4775 & _guard4776;
wire _guard4778 = cond_wire144_out;
wire _guard4779 = early_reset_static_par0_go_out;
wire _guard4780 = _guard4778 & _guard4779;
wire _guard4781 = cond_wire144_out;
wire _guard4782 = early_reset_static_par0_go_out;
wire _guard4783 = _guard4781 & _guard4782;
wire _guard4784 = cond_wire185_out;
wire _guard4785 = early_reset_static_par0_go_out;
wire _guard4786 = _guard4784 & _guard4785;
wire _guard4787 = cond_wire185_out;
wire _guard4788 = early_reset_static_par0_go_out;
wire _guard4789 = _guard4787 & _guard4788;
wire _guard4790 = cond_wire235_out;
wire _guard4791 = early_reset_static_par0_go_out;
wire _guard4792 = _guard4790 & _guard4791;
wire _guard4793 = cond_wire233_out;
wire _guard4794 = early_reset_static_par0_go_out;
wire _guard4795 = _guard4793 & _guard4794;
wire _guard4796 = fsm_out == 1'd0;
wire _guard4797 = cond_wire233_out;
wire _guard4798 = _guard4796 & _guard4797;
wire _guard4799 = fsm_out == 1'd0;
wire _guard4800 = _guard4798 & _guard4799;
wire _guard4801 = fsm_out == 1'd0;
wire _guard4802 = cond_wire235_out;
wire _guard4803 = _guard4801 & _guard4802;
wire _guard4804 = fsm_out == 1'd0;
wire _guard4805 = _guard4803 & _guard4804;
wire _guard4806 = _guard4800 | _guard4805;
wire _guard4807 = early_reset_static_par0_go_out;
wire _guard4808 = _guard4806 & _guard4807;
wire _guard4809 = fsm_out == 1'd0;
wire _guard4810 = cond_wire233_out;
wire _guard4811 = _guard4809 & _guard4810;
wire _guard4812 = fsm_out == 1'd0;
wire _guard4813 = _guard4811 & _guard4812;
wire _guard4814 = fsm_out == 1'd0;
wire _guard4815 = cond_wire235_out;
wire _guard4816 = _guard4814 & _guard4815;
wire _guard4817 = fsm_out == 1'd0;
wire _guard4818 = _guard4816 & _guard4817;
wire _guard4819 = _guard4813 | _guard4818;
wire _guard4820 = early_reset_static_par0_go_out;
wire _guard4821 = _guard4819 & _guard4820;
wire _guard4822 = fsm_out == 1'd0;
wire _guard4823 = cond_wire233_out;
wire _guard4824 = _guard4822 & _guard4823;
wire _guard4825 = fsm_out == 1'd0;
wire _guard4826 = _guard4824 & _guard4825;
wire _guard4827 = fsm_out == 1'd0;
wire _guard4828 = cond_wire235_out;
wire _guard4829 = _guard4827 & _guard4828;
wire _guard4830 = fsm_out == 1'd0;
wire _guard4831 = _guard4829 & _guard4830;
wire _guard4832 = _guard4826 | _guard4831;
wire _guard4833 = early_reset_static_par0_go_out;
wire _guard4834 = _guard4832 & _guard4833;
wire _guard4835 = cond_wire237_out;
wire _guard4836 = early_reset_static_par0_go_out;
wire _guard4837 = _guard4835 & _guard4836;
wire _guard4838 = cond_wire237_out;
wire _guard4839 = early_reset_static_par0_go_out;
wire _guard4840 = _guard4838 & _guard4839;
wire _guard4841 = fsm0_out == 5'd0;
wire _guard4842 = early_reset_static_seq_go_out;
wire _guard4843 = _guard4841 & _guard4842;
wire _guard4844 = early_reset_static_par0_go_out;
wire _guard4845 = _guard4843 | _guard4844;
wire _guard4846 = early_reset_static_par0_go_out;
wire _guard4847 = fsm0_out == 5'd0;
wire _guard4848 = early_reset_static_seq_go_out;
wire _guard4849 = _guard4847 & _guard4848;
wire _guard4850 = early_reset_static_par0_go_out;
wire _guard4851 = early_reset_static_par0_go_out;
wire _guard4852 = early_reset_static_par0_go_out;
wire _guard4853 = early_reset_static_par0_go_out;
wire _guard4854 = fsm0_out == 5'd0;
wire _guard4855 = early_reset_static_seq_go_out;
wire _guard4856 = _guard4854 & _guard4855;
wire _guard4857 = early_reset_static_par0_go_out;
wire _guard4858 = _guard4856 | _guard4857;
wire _guard4859 = fsm0_out == 5'd0;
wire _guard4860 = early_reset_static_seq_go_out;
wire _guard4861 = _guard4859 & _guard4860;
wire _guard4862 = early_reset_static_par0_go_out;
wire _guard4863 = early_reset_static_par0_go_out;
wire _guard4864 = early_reset_static_par0_go_out;
wire _guard4865 = early_reset_static_par0_go_out;
wire _guard4866 = early_reset_static_par0_go_out;
wire _guard4867 = early_reset_static_par0_go_out;
wire _guard4868 = early_reset_static_par0_go_out;
wire _guard4869 = early_reset_static_par0_go_out;
wire _guard4870 = early_reset_static_par0_go_out;
wire _guard4871 = fsm0_out == 5'd0;
wire _guard4872 = early_reset_static_seq_go_out;
wire _guard4873 = _guard4871 & _guard4872;
wire _guard4874 = early_reset_static_par0_go_out;
wire _guard4875 = _guard4873 | _guard4874;
wire _guard4876 = early_reset_static_par0_go_out;
wire _guard4877 = fsm0_out == 5'd0;
wire _guard4878 = early_reset_static_seq_go_out;
wire _guard4879 = _guard4877 & _guard4878;
wire _guard4880 = fsm0_out == 5'd0;
wire _guard4881 = early_reset_static_seq_go_out;
wire _guard4882 = _guard4880 & _guard4881;
wire _guard4883 = early_reset_static_par0_go_out;
wire _guard4884 = _guard4882 | _guard4883;
wire _guard4885 = fsm0_out == 5'd0;
wire _guard4886 = early_reset_static_seq_go_out;
wire _guard4887 = _guard4885 & _guard4886;
wire _guard4888 = early_reset_static_par0_go_out;
wire _guard4889 = fsm0_out == 5'd0;
wire _guard4890 = early_reset_static_seq_go_out;
wire _guard4891 = _guard4889 & _guard4890;
wire _guard4892 = early_reset_static_par0_go_out;
wire _guard4893 = _guard4891 | _guard4892;
wire _guard4894 = early_reset_static_par0_go_out;
wire _guard4895 = fsm0_out == 5'd0;
wire _guard4896 = early_reset_static_seq_go_out;
wire _guard4897 = _guard4895 & _guard4896;
wire _guard4898 = early_reset_static_par0_go_out;
wire _guard4899 = early_reset_static_par0_go_out;
wire _guard4900 = fsm0_out == 5'd0;
wire _guard4901 = early_reset_static_seq_go_out;
wire _guard4902 = _guard4900 & _guard4901;
wire _guard4903 = early_reset_static_par0_go_out;
wire _guard4904 = _guard4902 | _guard4903;
wire _guard4905 = early_reset_static_par0_go_out;
wire _guard4906 = fsm0_out == 5'd0;
wire _guard4907 = early_reset_static_seq_go_out;
wire _guard4908 = _guard4906 & _guard4907;
wire _guard4909 = early_reset_static_par0_go_out;
wire _guard4910 = early_reset_static_par0_go_out;
wire _guard4911 = early_reset_static_par0_go_out;
wire _guard4912 = early_reset_static_par0_go_out;
wire _guard4913 = early_reset_static_par0_go_out;
wire _guard4914 = early_reset_static_par0_go_out;
wire _guard4915 = ~_guard0;
wire _guard4916 = early_reset_static_par0_go_out;
wire _guard4917 = _guard4915 & _guard4916;
wire _guard4918 = early_reset_static_par0_go_out;
wire _guard4919 = early_reset_static_par0_go_out;
wire _guard4920 = early_reset_static_par0_go_out;
wire _guard4921 = early_reset_static_par0_go_out;
wire _guard4922 = ~_guard0;
wire _guard4923 = early_reset_static_par0_go_out;
wire _guard4924 = _guard4922 & _guard4923;
wire _guard4925 = early_reset_static_par0_go_out;
wire _guard4926 = early_reset_static_par0_go_out;
wire _guard4927 = early_reset_static_par0_go_out;
wire _guard4928 = ~_guard0;
wire _guard4929 = early_reset_static_par0_go_out;
wire _guard4930 = _guard4928 & _guard4929;
wire _guard4931 = early_reset_static_par0_go_out;
wire _guard4932 = early_reset_static_par0_go_out;
wire _guard4933 = ~_guard0;
wire _guard4934 = early_reset_static_par0_go_out;
wire _guard4935 = _guard4933 & _guard4934;
wire _guard4936 = early_reset_static_par0_go_out;
wire _guard4937 = ~_guard0;
wire _guard4938 = early_reset_static_par0_go_out;
wire _guard4939 = _guard4937 & _guard4938;
wire _guard4940 = early_reset_static_par0_go_out;
wire _guard4941 = early_reset_static_par0_go_out;
wire _guard4942 = ~_guard0;
wire _guard4943 = early_reset_static_par0_go_out;
wire _guard4944 = _guard4942 & _guard4943;
wire _guard4945 = early_reset_static_par0_go_out;
wire _guard4946 = early_reset_static_par0_go_out;
wire _guard4947 = early_reset_static_par0_go_out;
wire _guard4948 = early_reset_static_par0_go_out;
wire _guard4949 = ~_guard0;
wire _guard4950 = early_reset_static_par0_go_out;
wire _guard4951 = _guard4949 & _guard4950;
wire _guard4952 = early_reset_static_par0_go_out;
wire _guard4953 = early_reset_static_par0_go_out;
wire _guard4954 = early_reset_static_par0_go_out;
wire _guard4955 = early_reset_static_par0_go_out;
wire _guard4956 = early_reset_static_par0_go_out;
wire _guard4957 = early_reset_static_par0_go_out;
wire _guard4958 = ~_guard0;
wire _guard4959 = early_reset_static_par0_go_out;
wire _guard4960 = _guard4958 & _guard4959;
wire _guard4961 = early_reset_static_par0_go_out;
wire _guard4962 = early_reset_static_par0_go_out;
wire _guard4963 = early_reset_static_par0_go_out;
wire _guard4964 = early_reset_static_par0_go_out;
wire _guard4965 = early_reset_static_par0_go_out;
wire _guard4966 = ~_guard0;
wire _guard4967 = early_reset_static_par0_go_out;
wire _guard4968 = _guard4966 & _guard4967;
wire _guard4969 = ~_guard0;
wire _guard4970 = early_reset_static_par0_go_out;
wire _guard4971 = _guard4969 & _guard4970;
wire _guard4972 = early_reset_static_par0_go_out;
wire _guard4973 = ~_guard0;
wire _guard4974 = early_reset_static_par0_go_out;
wire _guard4975 = _guard4973 & _guard4974;
wire _guard4976 = early_reset_static_par0_go_out;
wire _guard4977 = early_reset_static_par0_go_out;
wire _guard4978 = early_reset_static_par0_go_out;
wire _guard4979 = early_reset_static_par0_go_out;
wire _guard4980 = ~_guard0;
wire _guard4981 = early_reset_static_par0_go_out;
wire _guard4982 = _guard4980 & _guard4981;
wire _guard4983 = early_reset_static_par0_go_out;
wire _guard4984 = early_reset_static_par0_go_out;
wire _guard4985 = early_reset_static_par0_go_out;
wire _guard4986 = early_reset_static_par0_go_out;
wire _guard4987 = early_reset_static_par0_go_out;
wire _guard4988 = ~_guard0;
wire _guard4989 = early_reset_static_par0_go_out;
wire _guard4990 = _guard4988 & _guard4989;
wire _guard4991 = early_reset_static_par0_go_out;
wire _guard4992 = ~_guard0;
wire _guard4993 = early_reset_static_par0_go_out;
wire _guard4994 = _guard4992 & _guard4993;
wire _guard4995 = ~_guard0;
wire _guard4996 = early_reset_static_par0_go_out;
wire _guard4997 = _guard4995 & _guard4996;
wire _guard4998 = early_reset_static_par0_go_out;
wire _guard4999 = ~_guard0;
wire _guard5000 = early_reset_static_par0_go_out;
wire _guard5001 = _guard4999 & _guard5000;
wire _guard5002 = early_reset_static_par0_go_out;
wire _guard5003 = early_reset_static_par0_go_out;
wire _guard5004 = early_reset_static_par0_go_out;
wire _guard5005 = early_reset_static_par0_go_out;
wire _guard5006 = early_reset_static_par0_go_out;
wire _guard5007 = early_reset_static_par0_go_out;
wire _guard5008 = early_reset_static_par0_go_out;
wire _guard5009 = early_reset_static_par0_go_out;
wire _guard5010 = ~_guard0;
wire _guard5011 = early_reset_static_par0_go_out;
wire _guard5012 = _guard5010 & _guard5011;
wire _guard5013 = early_reset_static_par0_go_out;
wire _guard5014 = early_reset_static_par0_go_out;
wire _guard5015 = early_reset_static_par0_go_out;
wire _guard5016 = ~_guard0;
wire _guard5017 = early_reset_static_par0_go_out;
wire _guard5018 = _guard5016 & _guard5017;
wire _guard5019 = ~_guard0;
wire _guard5020 = early_reset_static_par0_go_out;
wire _guard5021 = _guard5019 & _guard5020;
wire _guard5022 = early_reset_static_par0_go_out;
wire _guard5023 = ~_guard0;
wire _guard5024 = early_reset_static_par0_go_out;
wire _guard5025 = _guard5023 & _guard5024;
wire _guard5026 = early_reset_static_par0_go_out;
wire _guard5027 = early_reset_static_par0_go_out;
wire _guard5028 = early_reset_static_par0_go_out;
wire _guard5029 = ~_guard0;
wire _guard5030 = early_reset_static_par0_go_out;
wire _guard5031 = _guard5029 & _guard5030;
wire _guard5032 = early_reset_static_par0_go_out;
wire _guard5033 = early_reset_static_par0_go_out;
wire _guard5034 = early_reset_static_par0_go_out;
wire _guard5035 = early_reset_static_par0_go_out;
wire _guard5036 = early_reset_static_par0_go_out;
wire _guard5037 = early_reset_static_par0_go_out;
wire _guard5038 = ~_guard0;
wire _guard5039 = early_reset_static_par0_go_out;
wire _guard5040 = _guard5038 & _guard5039;
wire _guard5041 = ~_guard0;
wire _guard5042 = early_reset_static_par0_go_out;
wire _guard5043 = _guard5041 & _guard5042;
wire _guard5044 = early_reset_static_par0_go_out;
wire _guard5045 = ~_guard0;
wire _guard5046 = early_reset_static_par0_go_out;
wire _guard5047 = _guard5045 & _guard5046;
wire _guard5048 = early_reset_static_par0_go_out;
wire _guard5049 = early_reset_static_par0_go_out;
wire _guard5050 = ~_guard0;
wire _guard5051 = early_reset_static_par0_go_out;
wire _guard5052 = _guard5050 & _guard5051;
wire _guard5053 = early_reset_static_par0_go_out;
wire _guard5054 = early_reset_static_par0_go_out;
wire _guard5055 = wrapper_early_reset_static_seq_go_out;
wire _guard5056 = cond_wire9_out;
wire _guard5057 = early_reset_static_par0_go_out;
wire _guard5058 = _guard5056 & _guard5057;
wire _guard5059 = cond_wire9_out;
wire _guard5060 = early_reset_static_par0_go_out;
wire _guard5061 = _guard5059 & _guard5060;
wire _guard5062 = cond_wire6_out;
wire _guard5063 = early_reset_static_par0_go_out;
wire _guard5064 = _guard5062 & _guard5063;
wire _guard5065 = cond_wire6_out;
wire _guard5066 = early_reset_static_par0_go_out;
wire _guard5067 = _guard5065 & _guard5066;
wire _guard5068 = cond_wire111_out;
wire _guard5069 = early_reset_static_par0_go_out;
wire _guard5070 = _guard5068 & _guard5069;
wire _guard5071 = cond_wire111_out;
wire _guard5072 = early_reset_static_par0_go_out;
wire _guard5073 = _guard5071 & _guard5072;
wire _guard5074 = cond_wire119_out;
wire _guard5075 = early_reset_static_par0_go_out;
wire _guard5076 = _guard5074 & _guard5075;
wire _guard5077 = cond_wire119_out;
wire _guard5078 = early_reset_static_par0_go_out;
wire _guard5079 = _guard5077 & _guard5078;
wire _guard5080 = cond_wire111_out;
wire _guard5081 = early_reset_static_par0_go_out;
wire _guard5082 = _guard5080 & _guard5081;
wire _guard5083 = cond_wire111_out;
wire _guard5084 = early_reset_static_par0_go_out;
wire _guard5085 = _guard5083 & _guard5084;
wire _guard5086 = cond_wire115_out;
wire _guard5087 = early_reset_static_par0_go_out;
wire _guard5088 = _guard5086 & _guard5087;
wire _guard5089 = cond_wire115_out;
wire _guard5090 = early_reset_static_par0_go_out;
wire _guard5091 = _guard5089 & _guard5090;
wire _guard5092 = cond_wire189_out;
wire _guard5093 = early_reset_static_par0_go_out;
wire _guard5094 = _guard5092 & _guard5093;
wire _guard5095 = cond_wire189_out;
wire _guard5096 = early_reset_static_par0_go_out;
wire _guard5097 = _guard5095 & _guard5096;
wire _guard5098 = cond_wire193_out;
wire _guard5099 = early_reset_static_par0_go_out;
wire _guard5100 = _guard5098 & _guard5099;
wire _guard5101 = cond_wire193_out;
wire _guard5102 = early_reset_static_par0_go_out;
wire _guard5103 = _guard5101 & _guard5102;
wire _guard5104 = cond_wire226_out;
wire _guard5105 = early_reset_static_par0_go_out;
wire _guard5106 = _guard5104 & _guard5105;
wire _guard5107 = cond_wire226_out;
wire _guard5108 = early_reset_static_par0_go_out;
wire _guard5109 = _guard5107 & _guard5108;
wire _guard5110 = cond_wire243_out;
wire _guard5111 = early_reset_static_par0_go_out;
wire _guard5112 = _guard5110 & _guard5111;
wire _guard5113 = cond_wire243_out;
wire _guard5114 = early_reset_static_par0_go_out;
wire _guard5115 = _guard5113 & _guard5114;
wire _guard5116 = cond_wire260_out;
wire _guard5117 = early_reset_static_par0_go_out;
wire _guard5118 = _guard5116 & _guard5117;
wire _guard5119 = cond_wire258_out;
wire _guard5120 = early_reset_static_par0_go_out;
wire _guard5121 = _guard5119 & _guard5120;
wire _guard5122 = fsm_out == 1'd0;
wire _guard5123 = cond_wire258_out;
wire _guard5124 = _guard5122 & _guard5123;
wire _guard5125 = fsm_out == 1'd0;
wire _guard5126 = _guard5124 & _guard5125;
wire _guard5127 = fsm_out == 1'd0;
wire _guard5128 = cond_wire260_out;
wire _guard5129 = _guard5127 & _guard5128;
wire _guard5130 = fsm_out == 1'd0;
wire _guard5131 = _guard5129 & _guard5130;
wire _guard5132 = _guard5126 | _guard5131;
wire _guard5133 = early_reset_static_par0_go_out;
wire _guard5134 = _guard5132 & _guard5133;
wire _guard5135 = fsm_out == 1'd0;
wire _guard5136 = cond_wire258_out;
wire _guard5137 = _guard5135 & _guard5136;
wire _guard5138 = fsm_out == 1'd0;
wire _guard5139 = _guard5137 & _guard5138;
wire _guard5140 = fsm_out == 1'd0;
wire _guard5141 = cond_wire260_out;
wire _guard5142 = _guard5140 & _guard5141;
wire _guard5143 = fsm_out == 1'd0;
wire _guard5144 = _guard5142 & _guard5143;
wire _guard5145 = _guard5139 | _guard5144;
wire _guard5146 = early_reset_static_par0_go_out;
wire _guard5147 = _guard5145 & _guard5146;
wire _guard5148 = fsm_out == 1'd0;
wire _guard5149 = cond_wire258_out;
wire _guard5150 = _guard5148 & _guard5149;
wire _guard5151 = fsm_out == 1'd0;
wire _guard5152 = _guard5150 & _guard5151;
wire _guard5153 = fsm_out == 1'd0;
wire _guard5154 = cond_wire260_out;
wire _guard5155 = _guard5153 & _guard5154;
wire _guard5156 = fsm_out == 1'd0;
wire _guard5157 = _guard5155 & _guard5156;
wire _guard5158 = _guard5152 | _guard5157;
wire _guard5159 = early_reset_static_par0_go_out;
wire _guard5160 = _guard5158 & _guard5159;
wire _guard5161 = cond_wire264_out;
wire _guard5162 = early_reset_static_par0_go_out;
wire _guard5163 = _guard5161 & _guard5162;
wire _guard5164 = cond_wire262_out;
wire _guard5165 = early_reset_static_par0_go_out;
wire _guard5166 = _guard5164 & _guard5165;
wire _guard5167 = fsm_out == 1'd0;
wire _guard5168 = cond_wire262_out;
wire _guard5169 = _guard5167 & _guard5168;
wire _guard5170 = fsm_out == 1'd0;
wire _guard5171 = _guard5169 & _guard5170;
wire _guard5172 = fsm_out == 1'd0;
wire _guard5173 = cond_wire264_out;
wire _guard5174 = _guard5172 & _guard5173;
wire _guard5175 = fsm_out == 1'd0;
wire _guard5176 = _guard5174 & _guard5175;
wire _guard5177 = _guard5171 | _guard5176;
wire _guard5178 = early_reset_static_par0_go_out;
wire _guard5179 = _guard5177 & _guard5178;
wire _guard5180 = fsm_out == 1'd0;
wire _guard5181 = cond_wire262_out;
wire _guard5182 = _guard5180 & _guard5181;
wire _guard5183 = fsm_out == 1'd0;
wire _guard5184 = _guard5182 & _guard5183;
wire _guard5185 = fsm_out == 1'd0;
wire _guard5186 = cond_wire264_out;
wire _guard5187 = _guard5185 & _guard5186;
wire _guard5188 = fsm_out == 1'd0;
wire _guard5189 = _guard5187 & _guard5188;
wire _guard5190 = _guard5184 | _guard5189;
wire _guard5191 = early_reset_static_par0_go_out;
wire _guard5192 = _guard5190 & _guard5191;
wire _guard5193 = fsm_out == 1'd0;
wire _guard5194 = cond_wire262_out;
wire _guard5195 = _guard5193 & _guard5194;
wire _guard5196 = fsm_out == 1'd0;
wire _guard5197 = _guard5195 & _guard5196;
wire _guard5198 = fsm_out == 1'd0;
wire _guard5199 = cond_wire264_out;
wire _guard5200 = _guard5198 & _guard5199;
wire _guard5201 = fsm_out == 1'd0;
wire _guard5202 = _guard5200 & _guard5201;
wire _guard5203 = _guard5197 | _guard5202;
wire _guard5204 = early_reset_static_par0_go_out;
wire _guard5205 = _guard5203 & _guard5204;
wire _guard5206 = cond_wire_out;
wire _guard5207 = early_reset_static_par0_go_out;
wire _guard5208 = _guard5206 & _guard5207;
wire _guard5209 = cond_wire_out;
wire _guard5210 = early_reset_static_par0_go_out;
wire _guard5211 = _guard5209 & _guard5210;
wire _guard5212 = cond_wire_out;
wire _guard5213 = early_reset_static_par0_go_out;
wire _guard5214 = _guard5212 & _guard5213;
wire _guard5215 = cond_wire_out;
wire _guard5216 = early_reset_static_par0_go_out;
wire _guard5217 = _guard5215 & _guard5216;
wire _guard5218 = early_reset_static_par0_go_out;
wire _guard5219 = early_reset_static_par0_go_out;
wire _guard5220 = early_reset_static_par0_go_out;
wire _guard5221 = early_reset_static_par0_go_out;
wire _guard5222 = early_reset_static_par0_go_out;
wire _guard5223 = early_reset_static_par0_go_out;
wire _guard5224 = early_reset_static_par0_go_out;
wire _guard5225 = early_reset_static_par0_go_out;
wire _guard5226 = early_reset_static_par0_go_out;
wire _guard5227 = early_reset_static_par0_go_out;
wire _guard5228 = early_reset_static_par0_go_out;
wire _guard5229 = early_reset_static_par0_go_out;
wire _guard5230 = early_reset_static_par0_go_out;
wire _guard5231 = early_reset_static_par0_go_out;
wire _guard5232 = early_reset_static_par0_go_out;
wire _guard5233 = early_reset_static_par0_go_out;
wire _guard5234 = early_reset_static_par0_go_out;
wire _guard5235 = early_reset_static_par0_go_out;
wire _guard5236 = early_reset_static_par0_go_out;
wire _guard5237 = early_reset_static_par0_go_out;
wire _guard5238 = early_reset_static_par0_go_out;
wire _guard5239 = early_reset_static_par0_go_out;
wire _guard5240 = early_reset_static_par0_go_out;
wire _guard5241 = early_reset_static_par0_go_out;
wire _guard5242 = early_reset_static_par0_go_out;
wire _guard5243 = ~_guard0;
wire _guard5244 = early_reset_static_par0_go_out;
wire _guard5245 = _guard5243 & _guard5244;
wire _guard5246 = ~_guard0;
wire _guard5247 = early_reset_static_par0_go_out;
wire _guard5248 = _guard5246 & _guard5247;
wire _guard5249 = early_reset_static_par0_go_out;
wire _guard5250 = early_reset_static_par0_go_out;
wire _guard5251 = early_reset_static_par0_go_out;
wire _guard5252 = ~_guard0;
wire _guard5253 = early_reset_static_par0_go_out;
wire _guard5254 = _guard5252 & _guard5253;
wire _guard5255 = early_reset_static_par0_go_out;
wire _guard5256 = early_reset_static_par0_go_out;
wire _guard5257 = early_reset_static_par0_go_out;
wire _guard5258 = early_reset_static_par0_go_out;
wire _guard5259 = early_reset_static_par0_go_out;
wire _guard5260 = early_reset_static_par0_go_out;
wire _guard5261 = early_reset_static_par0_go_out;
wire _guard5262 = early_reset_static_par0_go_out;
wire _guard5263 = early_reset_static_par0_go_out;
wire _guard5264 = ~_guard0;
wire _guard5265 = early_reset_static_par0_go_out;
wire _guard5266 = _guard5264 & _guard5265;
wire _guard5267 = early_reset_static_par0_go_out;
wire _guard5268 = ~_guard0;
wire _guard5269 = early_reset_static_par0_go_out;
wire _guard5270 = _guard5268 & _guard5269;
wire _guard5271 = early_reset_static_par0_go_out;
wire _guard5272 = early_reset_static_par0_go_out;
wire _guard5273 = early_reset_static_par0_go_out;
wire _guard5274 = early_reset_static_par0_go_out;
wire _guard5275 = ~_guard0;
wire _guard5276 = early_reset_static_par0_go_out;
wire _guard5277 = _guard5275 & _guard5276;
wire _guard5278 = ~_guard0;
wire _guard5279 = early_reset_static_par0_go_out;
wire _guard5280 = _guard5278 & _guard5279;
wire _guard5281 = early_reset_static_par0_go_out;
wire _guard5282 = early_reset_static_par0_go_out;
wire _guard5283 = early_reset_static_par0_go_out;
wire _guard5284 = early_reset_static_par0_go_out;
wire _guard5285 = early_reset_static_par0_go_out;
wire _guard5286 = early_reset_static_par0_go_out;
wire _guard5287 = ~_guard0;
wire _guard5288 = early_reset_static_par0_go_out;
wire _guard5289 = _guard5287 & _guard5288;
wire _guard5290 = early_reset_static_par0_go_out;
wire _guard5291 = early_reset_static_par0_go_out;
wire _guard5292 = early_reset_static_par0_go_out;
wire _guard5293 = early_reset_static_par0_go_out;
wire _guard5294 = ~_guard0;
wire _guard5295 = early_reset_static_par0_go_out;
wire _guard5296 = _guard5294 & _guard5295;
wire _guard5297 = early_reset_static_par0_go_out;
wire _guard5298 = early_reset_static_par0_go_out;
wire _guard5299 = early_reset_static_par0_go_out;
wire _guard5300 = early_reset_static_par0_go_out;
wire _guard5301 = early_reset_static_par0_go_out;
wire _guard5302 = early_reset_static_par0_go_out;
wire _guard5303 = ~_guard0;
wire _guard5304 = early_reset_static_par0_go_out;
wire _guard5305 = _guard5303 & _guard5304;
wire _guard5306 = early_reset_static_par0_go_out;
wire _guard5307 = ~_guard0;
wire _guard5308 = early_reset_static_par0_go_out;
wire _guard5309 = _guard5307 & _guard5308;
wire _guard5310 = early_reset_static_par0_go_out;
wire _guard5311 = ~_guard0;
wire _guard5312 = early_reset_static_par0_go_out;
wire _guard5313 = _guard5311 & _guard5312;
wire _guard5314 = early_reset_static_par0_go_out;
wire _guard5315 = early_reset_static_par0_go_out;
wire _guard5316 = ~_guard0;
wire _guard5317 = early_reset_static_par0_go_out;
wire _guard5318 = _guard5316 & _guard5317;
wire _guard5319 = early_reset_static_par0_go_out;
wire _guard5320 = early_reset_static_par0_go_out;
wire _guard5321 = ~_guard0;
wire _guard5322 = early_reset_static_par0_go_out;
wire _guard5323 = _guard5321 & _guard5322;
wire _guard5324 = early_reset_static_par0_go_out;
wire _guard5325 = early_reset_static_par0_go_out;
wire _guard5326 = ~_guard0;
wire _guard5327 = early_reset_static_par0_go_out;
wire _guard5328 = _guard5326 & _guard5327;
wire _guard5329 = early_reset_static_par0_go_out;
wire _guard5330 = early_reset_static_par0_go_out;
wire _guard5331 = early_reset_static_par0_go_out;
wire _guard5332 = early_reset_static_par0_go_out;
wire _guard5333 = ~_guard0;
wire _guard5334 = early_reset_static_par0_go_out;
wire _guard5335 = _guard5333 & _guard5334;
wire _guard5336 = early_reset_static_par0_go_out;
wire _guard5337 = early_reset_static_par0_go_out;
wire _guard5338 = ~_guard0;
wire _guard5339 = early_reset_static_par0_go_out;
wire _guard5340 = _guard5338 & _guard5339;
wire _guard5341 = early_reset_static_par0_go_out;
wire _guard5342 = early_reset_static_par0_go_out;
wire _guard5343 = ~_guard0;
wire _guard5344 = early_reset_static_par0_go_out;
wire _guard5345 = _guard5343 & _guard5344;
wire _guard5346 = early_reset_static_par0_go_out;
wire _guard5347 = early_reset_static_par0_go_out;
wire _guard5348 = early_reset_static_par0_go_out;
wire _guard5349 = ~_guard0;
wire _guard5350 = early_reset_static_par0_go_out;
wire _guard5351 = _guard5349 & _guard5350;
wire _guard5352 = ~_guard0;
wire _guard5353 = early_reset_static_par0_go_out;
wire _guard5354 = _guard5352 & _guard5353;
wire _guard5355 = early_reset_static_par0_go_out;
wire _guard5356 = early_reset_static_par0_go_out;
wire _guard5357 = ~_guard0;
wire _guard5358 = early_reset_static_par0_go_out;
wire _guard5359 = _guard5357 & _guard5358;
wire _guard5360 = early_reset_static_par0_go_out;
wire _guard5361 = early_reset_static_par0_go_out;
wire _guard5362 = fsm0_out == 5'd0;
wire _guard5363 = signal_reg_out;
wire _guard5364 = _guard5362 & _guard5363;
wire _guard5365 = fsm0_out == 5'd0;
wire _guard5366 = signal_reg_out;
wire _guard5367 = ~_guard5366;
wire _guard5368 = _guard5365 & _guard5367;
wire _guard5369 = wrapper_early_reset_static_seq_go_out;
wire _guard5370 = _guard5368 & _guard5369;
wire _guard5371 = _guard5364 | _guard5370;
wire _guard5372 = fsm0_out == 5'd0;
wire _guard5373 = signal_reg_out;
wire _guard5374 = ~_guard5373;
wire _guard5375 = _guard5372 & _guard5374;
wire _guard5376 = wrapper_early_reset_static_seq_go_out;
wire _guard5377 = _guard5375 & _guard5376;
wire _guard5378 = fsm0_out == 5'd0;
wire _guard5379 = signal_reg_out;
wire _guard5380 = _guard5378 & _guard5379;
wire _guard5381 = cond_wire19_out;
wire _guard5382 = early_reset_static_par0_go_out;
wire _guard5383 = _guard5381 & _guard5382;
wire _guard5384 = cond_wire19_out;
wire _guard5385 = early_reset_static_par0_go_out;
wire _guard5386 = _guard5384 & _guard5385;
wire _guard5387 = cond_wire21_out;
wire _guard5388 = early_reset_static_par0_go_out;
wire _guard5389 = _guard5387 & _guard5388;
wire _guard5390 = cond_wire21_out;
wire _guard5391 = early_reset_static_par0_go_out;
wire _guard5392 = _guard5390 & _guard5391;
wire _guard5393 = cond_wire75_out;
wire _guard5394 = early_reset_static_par0_go_out;
wire _guard5395 = _guard5393 & _guard5394;
wire _guard5396 = cond_wire73_out;
wire _guard5397 = early_reset_static_par0_go_out;
wire _guard5398 = _guard5396 & _guard5397;
wire _guard5399 = fsm_out == 1'd0;
wire _guard5400 = cond_wire73_out;
wire _guard5401 = _guard5399 & _guard5400;
wire _guard5402 = fsm_out == 1'd0;
wire _guard5403 = _guard5401 & _guard5402;
wire _guard5404 = fsm_out == 1'd0;
wire _guard5405 = cond_wire75_out;
wire _guard5406 = _guard5404 & _guard5405;
wire _guard5407 = fsm_out == 1'd0;
wire _guard5408 = _guard5406 & _guard5407;
wire _guard5409 = _guard5403 | _guard5408;
wire _guard5410 = early_reset_static_par0_go_out;
wire _guard5411 = _guard5409 & _guard5410;
wire _guard5412 = fsm_out == 1'd0;
wire _guard5413 = cond_wire73_out;
wire _guard5414 = _guard5412 & _guard5413;
wire _guard5415 = fsm_out == 1'd0;
wire _guard5416 = _guard5414 & _guard5415;
wire _guard5417 = fsm_out == 1'd0;
wire _guard5418 = cond_wire75_out;
wire _guard5419 = _guard5417 & _guard5418;
wire _guard5420 = fsm_out == 1'd0;
wire _guard5421 = _guard5419 & _guard5420;
wire _guard5422 = _guard5416 | _guard5421;
wire _guard5423 = early_reset_static_par0_go_out;
wire _guard5424 = _guard5422 & _guard5423;
wire _guard5425 = fsm_out == 1'd0;
wire _guard5426 = cond_wire73_out;
wire _guard5427 = _guard5425 & _guard5426;
wire _guard5428 = fsm_out == 1'd0;
wire _guard5429 = _guard5427 & _guard5428;
wire _guard5430 = fsm_out == 1'd0;
wire _guard5431 = cond_wire75_out;
wire _guard5432 = _guard5430 & _guard5431;
wire _guard5433 = fsm_out == 1'd0;
wire _guard5434 = _guard5432 & _guard5433;
wire _guard5435 = _guard5429 | _guard5434;
wire _guard5436 = early_reset_static_par0_go_out;
wire _guard5437 = _guard5435 & _guard5436;
wire _guard5438 = cond_wire74_out;
wire _guard5439 = early_reset_static_par0_go_out;
wire _guard5440 = _guard5438 & _guard5439;
wire _guard5441 = cond_wire74_out;
wire _guard5442 = early_reset_static_par0_go_out;
wire _guard5443 = _guard5441 & _guard5442;
wire _guard5444 = cond_wire49_out;
wire _guard5445 = early_reset_static_par0_go_out;
wire _guard5446 = _guard5444 & _guard5445;
wire _guard5447 = cond_wire49_out;
wire _guard5448 = early_reset_static_par0_go_out;
wire _guard5449 = _guard5447 & _guard5448;
wire _guard5450 = cond_wire90_out;
wire _guard5451 = early_reset_static_par0_go_out;
wire _guard5452 = _guard5450 & _guard5451;
wire _guard5453 = cond_wire90_out;
wire _guard5454 = early_reset_static_par0_go_out;
wire _guard5455 = _guard5453 & _guard5454;
wire _guard5456 = cond_wire127_out;
wire _guard5457 = early_reset_static_par0_go_out;
wire _guard5458 = _guard5456 & _guard5457;
wire _guard5459 = cond_wire127_out;
wire _guard5460 = early_reset_static_par0_go_out;
wire _guard5461 = _guard5459 & _guard5460;
wire _guard5462 = cond_wire157_out;
wire _guard5463 = early_reset_static_par0_go_out;
wire _guard5464 = _guard5462 & _guard5463;
wire _guard5465 = cond_wire155_out;
wire _guard5466 = early_reset_static_par0_go_out;
wire _guard5467 = _guard5465 & _guard5466;
wire _guard5468 = fsm_out == 1'd0;
wire _guard5469 = cond_wire155_out;
wire _guard5470 = _guard5468 & _guard5469;
wire _guard5471 = fsm_out == 1'd0;
wire _guard5472 = _guard5470 & _guard5471;
wire _guard5473 = fsm_out == 1'd0;
wire _guard5474 = cond_wire157_out;
wire _guard5475 = _guard5473 & _guard5474;
wire _guard5476 = fsm_out == 1'd0;
wire _guard5477 = _guard5475 & _guard5476;
wire _guard5478 = _guard5472 | _guard5477;
wire _guard5479 = early_reset_static_par0_go_out;
wire _guard5480 = _guard5478 & _guard5479;
wire _guard5481 = fsm_out == 1'd0;
wire _guard5482 = cond_wire155_out;
wire _guard5483 = _guard5481 & _guard5482;
wire _guard5484 = fsm_out == 1'd0;
wire _guard5485 = _guard5483 & _guard5484;
wire _guard5486 = fsm_out == 1'd0;
wire _guard5487 = cond_wire157_out;
wire _guard5488 = _guard5486 & _guard5487;
wire _guard5489 = fsm_out == 1'd0;
wire _guard5490 = _guard5488 & _guard5489;
wire _guard5491 = _guard5485 | _guard5490;
wire _guard5492 = early_reset_static_par0_go_out;
wire _guard5493 = _guard5491 & _guard5492;
wire _guard5494 = fsm_out == 1'd0;
wire _guard5495 = cond_wire155_out;
wire _guard5496 = _guard5494 & _guard5495;
wire _guard5497 = fsm_out == 1'd0;
wire _guard5498 = _guard5496 & _guard5497;
wire _guard5499 = fsm_out == 1'd0;
wire _guard5500 = cond_wire157_out;
wire _guard5501 = _guard5499 & _guard5500;
wire _guard5502 = fsm_out == 1'd0;
wire _guard5503 = _guard5501 & _guard5502;
wire _guard5504 = _guard5498 | _guard5503;
wire _guard5505 = early_reset_static_par0_go_out;
wire _guard5506 = _guard5504 & _guard5505;
wire _guard5507 = cond_wire152_out;
wire _guard5508 = early_reset_static_par0_go_out;
wire _guard5509 = _guard5507 & _guard5508;
wire _guard5510 = cond_wire152_out;
wire _guard5511 = early_reset_static_par0_go_out;
wire _guard5512 = _guard5510 & _guard5511;
wire _guard5513 = cond_wire169_out;
wire _guard5514 = early_reset_static_par0_go_out;
wire _guard5515 = _guard5513 & _guard5514;
wire _guard5516 = cond_wire167_out;
wire _guard5517 = early_reset_static_par0_go_out;
wire _guard5518 = _guard5516 & _guard5517;
wire _guard5519 = fsm_out == 1'd0;
wire _guard5520 = cond_wire167_out;
wire _guard5521 = _guard5519 & _guard5520;
wire _guard5522 = fsm_out == 1'd0;
wire _guard5523 = _guard5521 & _guard5522;
wire _guard5524 = fsm_out == 1'd0;
wire _guard5525 = cond_wire169_out;
wire _guard5526 = _guard5524 & _guard5525;
wire _guard5527 = fsm_out == 1'd0;
wire _guard5528 = _guard5526 & _guard5527;
wire _guard5529 = _guard5523 | _guard5528;
wire _guard5530 = early_reset_static_par0_go_out;
wire _guard5531 = _guard5529 & _guard5530;
wire _guard5532 = fsm_out == 1'd0;
wire _guard5533 = cond_wire167_out;
wire _guard5534 = _guard5532 & _guard5533;
wire _guard5535 = fsm_out == 1'd0;
wire _guard5536 = _guard5534 & _guard5535;
wire _guard5537 = fsm_out == 1'd0;
wire _guard5538 = cond_wire169_out;
wire _guard5539 = _guard5537 & _guard5538;
wire _guard5540 = fsm_out == 1'd0;
wire _guard5541 = _guard5539 & _guard5540;
wire _guard5542 = _guard5536 | _guard5541;
wire _guard5543 = early_reset_static_par0_go_out;
wire _guard5544 = _guard5542 & _guard5543;
wire _guard5545 = fsm_out == 1'd0;
wire _guard5546 = cond_wire167_out;
wire _guard5547 = _guard5545 & _guard5546;
wire _guard5548 = fsm_out == 1'd0;
wire _guard5549 = _guard5547 & _guard5548;
wire _guard5550 = fsm_out == 1'd0;
wire _guard5551 = cond_wire169_out;
wire _guard5552 = _guard5550 & _guard5551;
wire _guard5553 = fsm_out == 1'd0;
wire _guard5554 = _guard5552 & _guard5553;
wire _guard5555 = _guard5549 | _guard5554;
wire _guard5556 = early_reset_static_par0_go_out;
wire _guard5557 = _guard5555 & _guard5556;
wire _guard5558 = cond_wire189_out;
wire _guard5559 = early_reset_static_par0_go_out;
wire _guard5560 = _guard5558 & _guard5559;
wire _guard5561 = cond_wire189_out;
wire _guard5562 = early_reset_static_par0_go_out;
wire _guard5563 = _guard5561 & _guard5562;
wire _guard5564 = cond_wire237_out;
wire _guard5565 = early_reset_static_par0_go_out;
wire _guard5566 = _guard5564 & _guard5565;
wire _guard5567 = cond_wire237_out;
wire _guard5568 = early_reset_static_par0_go_out;
wire _guard5569 = _guard5567 & _guard5568;
wire _guard5570 = cond_wire218_out;
wire _guard5571 = early_reset_static_par0_go_out;
wire _guard5572 = _guard5570 & _guard5571;
wire _guard5573 = cond_wire218_out;
wire _guard5574 = early_reset_static_par0_go_out;
wire _guard5575 = _guard5573 & _guard5574;
wire _guard5576 = cond_wire230_out;
wire _guard5577 = early_reset_static_par0_go_out;
wire _guard5578 = _guard5576 & _guard5577;
wire _guard5579 = cond_wire230_out;
wire _guard5580 = early_reset_static_par0_go_out;
wire _guard5581 = _guard5579 & _guard5580;
wire _guard5582 = cond_wire4_out;
wire _guard5583 = early_reset_static_par0_go_out;
wire _guard5584 = _guard5582 & _guard5583;
wire _guard5585 = cond_wire4_out;
wire _guard5586 = early_reset_static_par0_go_out;
wire _guard5587 = _guard5585 & _guard5586;
wire _guard5588 = fsm0_out == 5'd0;
wire _guard5589 = early_reset_static_seq_go_out;
wire _guard5590 = _guard5588 & _guard5589;
wire _guard5591 = cond_wire14_out;
wire _guard5592 = early_reset_static_par0_go_out;
wire _guard5593 = _guard5591 & _guard5592;
wire _guard5594 = _guard5590 | _guard5593;
wire _guard5595 = cond_wire14_out;
wire _guard5596 = early_reset_static_par0_go_out;
wire _guard5597 = _guard5595 & _guard5596;
wire _guard5598 = fsm0_out == 5'd0;
wire _guard5599 = early_reset_static_seq_go_out;
wire _guard5600 = _guard5598 & _guard5599;
wire _guard5601 = cond_wire138_out;
wire _guard5602 = early_reset_static_par0_go_out;
wire _guard5603 = _guard5601 & _guard5602;
wire _guard5604 = cond_wire138_out;
wire _guard5605 = early_reset_static_par0_go_out;
wire _guard5606 = _guard5604 & _guard5605;
wire _guard5607 = fsm0_out == 5'd0;
wire _guard5608 = early_reset_static_seq_go_out;
wire _guard5609 = _guard5607 & _guard5608;
wire _guard5610 = early_reset_static_par0_go_out;
wire _guard5611 = _guard5609 | _guard5610;
wire _guard5612 = early_reset_static_par0_go_out;
wire _guard5613 = fsm0_out == 5'd0;
wire _guard5614 = early_reset_static_seq_go_out;
wire _guard5615 = _guard5613 & _guard5614;
wire _guard5616 = early_reset_static_par0_go_out;
wire _guard5617 = early_reset_static_par0_go_out;
wire _guard5618 = early_reset_static_par0_go_out;
wire _guard5619 = early_reset_static_par0_go_out;
wire _guard5620 = early_reset_static_par0_go_out;
wire _guard5621 = early_reset_static_par0_go_out;
wire _guard5622 = early_reset_static_par0_go_out;
wire _guard5623 = early_reset_static_par0_go_out;
wire _guard5624 = early_reset_static_par0_go_out;
wire _guard5625 = early_reset_static_par0_go_out;
wire _guard5626 = fsm0_out == 5'd0;
wire _guard5627 = early_reset_static_seq_go_out;
wire _guard5628 = _guard5626 & _guard5627;
wire _guard5629 = early_reset_static_par0_go_out;
wire _guard5630 = _guard5628 | _guard5629;
wire _guard5631 = early_reset_static_par0_go_out;
wire _guard5632 = fsm0_out == 5'd0;
wire _guard5633 = early_reset_static_seq_go_out;
wire _guard5634 = _guard5632 & _guard5633;
wire _guard5635 = early_reset_static_par0_go_out;
wire _guard5636 = early_reset_static_par0_go_out;
wire _guard5637 = fsm0_out == 5'd0;
wire _guard5638 = early_reset_static_seq_go_out;
wire _guard5639 = _guard5637 & _guard5638;
wire _guard5640 = early_reset_static_par0_go_out;
wire _guard5641 = _guard5639 | _guard5640;
wire _guard5642 = early_reset_static_par0_go_out;
wire _guard5643 = fsm0_out == 5'd0;
wire _guard5644 = early_reset_static_seq_go_out;
wire _guard5645 = _guard5643 & _guard5644;
wire _guard5646 = early_reset_static_par0_go_out;
wire _guard5647 = early_reset_static_par0_go_out;
wire _guard5648 = early_reset_static_par0_go_out;
wire _guard5649 = early_reset_static_par0_go_out;
wire _guard5650 = early_reset_static_par0_go_out;
wire _guard5651 = early_reset_static_par0_go_out;
wire _guard5652 = ~_guard0;
wire _guard5653 = early_reset_static_par0_go_out;
wire _guard5654 = _guard5652 & _guard5653;
wire _guard5655 = early_reset_static_par0_go_out;
wire _guard5656 = ~_guard0;
wire _guard5657 = early_reset_static_par0_go_out;
wire _guard5658 = _guard5656 & _guard5657;
wire _guard5659 = early_reset_static_par0_go_out;
wire _guard5660 = early_reset_static_par0_go_out;
wire _guard5661 = early_reset_static_par0_go_out;
wire _guard5662 = early_reset_static_par0_go_out;
wire _guard5663 = early_reset_static_par0_go_out;
wire _guard5664 = early_reset_static_par0_go_out;
wire _guard5665 = ~_guard0;
wire _guard5666 = early_reset_static_par0_go_out;
wire _guard5667 = _guard5665 & _guard5666;
wire _guard5668 = early_reset_static_par0_go_out;
wire _guard5669 = ~_guard0;
wire _guard5670 = early_reset_static_par0_go_out;
wire _guard5671 = _guard5669 & _guard5670;
wire _guard5672 = early_reset_static_par0_go_out;
wire _guard5673 = ~_guard0;
wire _guard5674 = early_reset_static_par0_go_out;
wire _guard5675 = _guard5673 & _guard5674;
wire _guard5676 = ~_guard0;
wire _guard5677 = early_reset_static_par0_go_out;
wire _guard5678 = _guard5676 & _guard5677;
wire _guard5679 = early_reset_static_par0_go_out;
wire _guard5680 = early_reset_static_par0_go_out;
wire _guard5681 = ~_guard0;
wire _guard5682 = early_reset_static_par0_go_out;
wire _guard5683 = _guard5681 & _guard5682;
wire _guard5684 = early_reset_static_par0_go_out;
wire _guard5685 = ~_guard0;
wire _guard5686 = early_reset_static_par0_go_out;
wire _guard5687 = _guard5685 & _guard5686;
wire _guard5688 = early_reset_static_par0_go_out;
wire _guard5689 = early_reset_static_par0_go_out;
wire _guard5690 = early_reset_static_par0_go_out;
wire _guard5691 = early_reset_static_par0_go_out;
wire _guard5692 = early_reset_static_par0_go_out;
wire _guard5693 = ~_guard0;
wire _guard5694 = early_reset_static_par0_go_out;
wire _guard5695 = _guard5693 & _guard5694;
wire _guard5696 = early_reset_static_par0_go_out;
wire _guard5697 = ~_guard0;
wire _guard5698 = early_reset_static_par0_go_out;
wire _guard5699 = _guard5697 & _guard5698;
wire _guard5700 = early_reset_static_par0_go_out;
wire _guard5701 = early_reset_static_par0_go_out;
wire _guard5702 = early_reset_static_par0_go_out;
wire _guard5703 = early_reset_static_par0_go_out;
wire _guard5704 = early_reset_static_par0_go_out;
wire _guard5705 = ~_guard0;
wire _guard5706 = early_reset_static_par0_go_out;
wire _guard5707 = _guard5705 & _guard5706;
wire _guard5708 = early_reset_static_par0_go_out;
wire _guard5709 = early_reset_static_par0_go_out;
wire _guard5710 = ~_guard0;
wire _guard5711 = early_reset_static_par0_go_out;
wire _guard5712 = _guard5710 & _guard5711;
wire _guard5713 = early_reset_static_par0_go_out;
wire _guard5714 = early_reset_static_par0_go_out;
wire _guard5715 = early_reset_static_par0_go_out;
wire _guard5716 = early_reset_static_par0_go_out;
wire _guard5717 = early_reset_static_par0_go_out;
wire _guard5718 = early_reset_static_par0_go_out;
wire _guard5719 = early_reset_static_par0_go_out;
wire _guard5720 = early_reset_static_par0_go_out;
wire _guard5721 = early_reset_static_par0_go_out;
wire _guard5722 = early_reset_static_par0_go_out;
wire _guard5723 = ~_guard0;
wire _guard5724 = early_reset_static_par0_go_out;
wire _guard5725 = _guard5723 & _guard5724;
wire _guard5726 = ~_guard0;
wire _guard5727 = early_reset_static_par0_go_out;
wire _guard5728 = _guard5726 & _guard5727;
wire _guard5729 = early_reset_static_par0_go_out;
wire _guard5730 = early_reset_static_par0_go_out;
wire _guard5731 = early_reset_static_par0_go_out;
wire _guard5732 = early_reset_static_par0_go_out;
wire _guard5733 = early_reset_static_par0_go_out;
wire _guard5734 = early_reset_static_par0_go_out;
wire _guard5735 = early_reset_static_par0_go_out;
wire _guard5736 = early_reset_static_par0_go_out;
wire _guard5737 = early_reset_static_par0_go_out;
wire _guard5738 = early_reset_static_par0_go_out;
wire _guard5739 = early_reset_static_par0_go_out;
wire _guard5740 = ~_guard0;
wire _guard5741 = early_reset_static_par0_go_out;
wire _guard5742 = _guard5740 & _guard5741;
wire _guard5743 = early_reset_static_par0_go_out;
wire _guard5744 = ~_guard0;
wire _guard5745 = early_reset_static_par0_go_out;
wire _guard5746 = _guard5744 & _guard5745;
wire _guard5747 = early_reset_static_par0_go_out;
wire _guard5748 = early_reset_static_par0_go_out;
wire _guard5749 = ~_guard0;
wire _guard5750 = early_reset_static_par0_go_out;
wire _guard5751 = _guard5749 & _guard5750;
wire _guard5752 = early_reset_static_par0_go_out;
wire _guard5753 = early_reset_static_par0_go_out;
wire _guard5754 = ~_guard0;
wire _guard5755 = early_reset_static_par0_go_out;
wire _guard5756 = _guard5754 & _guard5755;
wire _guard5757 = early_reset_static_par0_go_out;
wire _guard5758 = early_reset_static_par0_go_out;
wire _guard5759 = early_reset_static_par0_go_out;
wire _guard5760 = cond_wire2_out;
wire _guard5761 = early_reset_static_par0_go_out;
wire _guard5762 = _guard5760 & _guard5761;
wire _guard5763 = cond_wire0_out;
wire _guard5764 = early_reset_static_par0_go_out;
wire _guard5765 = _guard5763 & _guard5764;
wire _guard5766 = fsm_out == 1'd0;
wire _guard5767 = cond_wire0_out;
wire _guard5768 = _guard5766 & _guard5767;
wire _guard5769 = fsm_out == 1'd0;
wire _guard5770 = _guard5768 & _guard5769;
wire _guard5771 = fsm_out == 1'd0;
wire _guard5772 = cond_wire2_out;
wire _guard5773 = _guard5771 & _guard5772;
wire _guard5774 = fsm_out == 1'd0;
wire _guard5775 = _guard5773 & _guard5774;
wire _guard5776 = _guard5770 | _guard5775;
wire _guard5777 = early_reset_static_par0_go_out;
wire _guard5778 = _guard5776 & _guard5777;
wire _guard5779 = fsm_out == 1'd0;
wire _guard5780 = cond_wire0_out;
wire _guard5781 = _guard5779 & _guard5780;
wire _guard5782 = fsm_out == 1'd0;
wire _guard5783 = _guard5781 & _guard5782;
wire _guard5784 = fsm_out == 1'd0;
wire _guard5785 = cond_wire2_out;
wire _guard5786 = _guard5784 & _guard5785;
wire _guard5787 = fsm_out == 1'd0;
wire _guard5788 = _guard5786 & _guard5787;
wire _guard5789 = _guard5783 | _guard5788;
wire _guard5790 = early_reset_static_par0_go_out;
wire _guard5791 = _guard5789 & _guard5790;
wire _guard5792 = fsm_out == 1'd0;
wire _guard5793 = cond_wire0_out;
wire _guard5794 = _guard5792 & _guard5793;
wire _guard5795 = fsm_out == 1'd0;
wire _guard5796 = _guard5794 & _guard5795;
wire _guard5797 = fsm_out == 1'd0;
wire _guard5798 = cond_wire2_out;
wire _guard5799 = _guard5797 & _guard5798;
wire _guard5800 = fsm_out == 1'd0;
wire _guard5801 = _guard5799 & _guard5800;
wire _guard5802 = _guard5796 | _guard5801;
wire _guard5803 = early_reset_static_par0_go_out;
wire _guard5804 = _guard5802 & _guard5803;
wire _guard5805 = cond_wire61_out;
wire _guard5806 = early_reset_static_par0_go_out;
wire _guard5807 = _guard5805 & _guard5806;
wire _guard5808 = cond_wire61_out;
wire _guard5809 = early_reset_static_par0_go_out;
wire _guard5810 = _guard5808 & _guard5809;
wire _guard5811 = cond_wire120_out;
wire _guard5812 = early_reset_static_par0_go_out;
wire _guard5813 = _guard5811 & _guard5812;
wire _guard5814 = cond_wire118_out;
wire _guard5815 = early_reset_static_par0_go_out;
wire _guard5816 = _guard5814 & _guard5815;
wire _guard5817 = fsm_out == 1'd0;
wire _guard5818 = cond_wire118_out;
wire _guard5819 = _guard5817 & _guard5818;
wire _guard5820 = fsm_out == 1'd0;
wire _guard5821 = _guard5819 & _guard5820;
wire _guard5822 = fsm_out == 1'd0;
wire _guard5823 = cond_wire120_out;
wire _guard5824 = _guard5822 & _guard5823;
wire _guard5825 = fsm_out == 1'd0;
wire _guard5826 = _guard5824 & _guard5825;
wire _guard5827 = _guard5821 | _guard5826;
wire _guard5828 = early_reset_static_par0_go_out;
wire _guard5829 = _guard5827 & _guard5828;
wire _guard5830 = fsm_out == 1'd0;
wire _guard5831 = cond_wire118_out;
wire _guard5832 = _guard5830 & _guard5831;
wire _guard5833 = fsm_out == 1'd0;
wire _guard5834 = _guard5832 & _guard5833;
wire _guard5835 = fsm_out == 1'd0;
wire _guard5836 = cond_wire120_out;
wire _guard5837 = _guard5835 & _guard5836;
wire _guard5838 = fsm_out == 1'd0;
wire _guard5839 = _guard5837 & _guard5838;
wire _guard5840 = _guard5834 | _guard5839;
wire _guard5841 = early_reset_static_par0_go_out;
wire _guard5842 = _guard5840 & _guard5841;
wire _guard5843 = fsm_out == 1'd0;
wire _guard5844 = cond_wire118_out;
wire _guard5845 = _guard5843 & _guard5844;
wire _guard5846 = fsm_out == 1'd0;
wire _guard5847 = _guard5845 & _guard5846;
wire _guard5848 = fsm_out == 1'd0;
wire _guard5849 = cond_wire120_out;
wire _guard5850 = _guard5848 & _guard5849;
wire _guard5851 = fsm_out == 1'd0;
wire _guard5852 = _guard5850 & _guard5851;
wire _guard5853 = _guard5847 | _guard5852;
wire _guard5854 = early_reset_static_par0_go_out;
wire _guard5855 = _guard5853 & _guard5854;
wire _guard5856 = cond_wire86_out;
wire _guard5857 = early_reset_static_par0_go_out;
wire _guard5858 = _guard5856 & _guard5857;
wire _guard5859 = cond_wire86_out;
wire _guard5860 = early_reset_static_par0_go_out;
wire _guard5861 = _guard5859 & _guard5860;
wire _guard5862 = cond_wire119_out;
wire _guard5863 = early_reset_static_par0_go_out;
wire _guard5864 = _guard5862 & _guard5863;
wire _guard5865 = cond_wire119_out;
wire _guard5866 = early_reset_static_par0_go_out;
wire _guard5867 = _guard5865 & _guard5866;
wire _guard5868 = cond_wire131_out;
wire _guard5869 = early_reset_static_par0_go_out;
wire _guard5870 = _guard5868 & _guard5869;
wire _guard5871 = cond_wire131_out;
wire _guard5872 = early_reset_static_par0_go_out;
wire _guard5873 = _guard5871 & _guard5872;
wire _guard5874 = cond_wire198_out;
wire _guard5875 = early_reset_static_par0_go_out;
wire _guard5876 = _guard5874 & _guard5875;
wire _guard5877 = cond_wire196_out;
wire _guard5878 = early_reset_static_par0_go_out;
wire _guard5879 = _guard5877 & _guard5878;
wire _guard5880 = fsm_out == 1'd0;
wire _guard5881 = cond_wire196_out;
wire _guard5882 = _guard5880 & _guard5881;
wire _guard5883 = fsm_out == 1'd0;
wire _guard5884 = _guard5882 & _guard5883;
wire _guard5885 = fsm_out == 1'd0;
wire _guard5886 = cond_wire198_out;
wire _guard5887 = _guard5885 & _guard5886;
wire _guard5888 = fsm_out == 1'd0;
wire _guard5889 = _guard5887 & _guard5888;
wire _guard5890 = _guard5884 | _guard5889;
wire _guard5891 = early_reset_static_par0_go_out;
wire _guard5892 = _guard5890 & _guard5891;
wire _guard5893 = fsm_out == 1'd0;
wire _guard5894 = cond_wire196_out;
wire _guard5895 = _guard5893 & _guard5894;
wire _guard5896 = fsm_out == 1'd0;
wire _guard5897 = _guard5895 & _guard5896;
wire _guard5898 = fsm_out == 1'd0;
wire _guard5899 = cond_wire198_out;
wire _guard5900 = _guard5898 & _guard5899;
wire _guard5901 = fsm_out == 1'd0;
wire _guard5902 = _guard5900 & _guard5901;
wire _guard5903 = _guard5897 | _guard5902;
wire _guard5904 = early_reset_static_par0_go_out;
wire _guard5905 = _guard5903 & _guard5904;
wire _guard5906 = fsm_out == 1'd0;
wire _guard5907 = cond_wire196_out;
wire _guard5908 = _guard5906 & _guard5907;
wire _guard5909 = fsm_out == 1'd0;
wire _guard5910 = _guard5908 & _guard5909;
wire _guard5911 = fsm_out == 1'd0;
wire _guard5912 = cond_wire198_out;
wire _guard5913 = _guard5911 & _guard5912;
wire _guard5914 = fsm_out == 1'd0;
wire _guard5915 = _guard5913 & _guard5914;
wire _guard5916 = _guard5910 | _guard5915;
wire _guard5917 = early_reset_static_par0_go_out;
wire _guard5918 = _guard5916 & _guard5917;
wire _guard5919 = cond_wire164_out;
wire _guard5920 = early_reset_static_par0_go_out;
wire _guard5921 = _guard5919 & _guard5920;
wire _guard5922 = cond_wire164_out;
wire _guard5923 = early_reset_static_par0_go_out;
wire _guard5924 = _guard5922 & _guard5923;
wire _guard5925 = cond_wire181_out;
wire _guard5926 = early_reset_static_par0_go_out;
wire _guard5927 = _guard5925 & _guard5926;
wire _guard5928 = cond_wire181_out;
wire _guard5929 = early_reset_static_par0_go_out;
wire _guard5930 = _guard5928 & _guard5929;
wire _guard5931 = cond_wire244_out;
wire _guard5932 = early_reset_static_par0_go_out;
wire _guard5933 = _guard5931 & _guard5932;
wire _guard5934 = cond_wire242_out;
wire _guard5935 = early_reset_static_par0_go_out;
wire _guard5936 = _guard5934 & _guard5935;
wire _guard5937 = fsm_out == 1'd0;
wire _guard5938 = cond_wire242_out;
wire _guard5939 = _guard5937 & _guard5938;
wire _guard5940 = fsm_out == 1'd0;
wire _guard5941 = _guard5939 & _guard5940;
wire _guard5942 = fsm_out == 1'd0;
wire _guard5943 = cond_wire244_out;
wire _guard5944 = _guard5942 & _guard5943;
wire _guard5945 = fsm_out == 1'd0;
wire _guard5946 = _guard5944 & _guard5945;
wire _guard5947 = _guard5941 | _guard5946;
wire _guard5948 = early_reset_static_par0_go_out;
wire _guard5949 = _guard5947 & _guard5948;
wire _guard5950 = fsm_out == 1'd0;
wire _guard5951 = cond_wire242_out;
wire _guard5952 = _guard5950 & _guard5951;
wire _guard5953 = fsm_out == 1'd0;
wire _guard5954 = _guard5952 & _guard5953;
wire _guard5955 = fsm_out == 1'd0;
wire _guard5956 = cond_wire244_out;
wire _guard5957 = _guard5955 & _guard5956;
wire _guard5958 = fsm_out == 1'd0;
wire _guard5959 = _guard5957 & _guard5958;
wire _guard5960 = _guard5954 | _guard5959;
wire _guard5961 = early_reset_static_par0_go_out;
wire _guard5962 = _guard5960 & _guard5961;
wire _guard5963 = fsm_out == 1'd0;
wire _guard5964 = cond_wire242_out;
wire _guard5965 = _guard5963 & _guard5964;
wire _guard5966 = fsm_out == 1'd0;
wire _guard5967 = _guard5965 & _guard5966;
wire _guard5968 = fsm_out == 1'd0;
wire _guard5969 = cond_wire244_out;
wire _guard5970 = _guard5968 & _guard5969;
wire _guard5971 = fsm_out == 1'd0;
wire _guard5972 = _guard5970 & _guard5971;
wire _guard5973 = _guard5967 | _guard5972;
wire _guard5974 = early_reset_static_par0_go_out;
wire _guard5975 = _guard5973 & _guard5974;
wire _guard5976 = cond_wire9_out;
wire _guard5977 = early_reset_static_par0_go_out;
wire _guard5978 = _guard5976 & _guard5977;
wire _guard5979 = cond_wire9_out;
wire _guard5980 = early_reset_static_par0_go_out;
wire _guard5981 = _guard5979 & _guard5980;
wire _guard5982 = cond_wire24_out;
wire _guard5983 = early_reset_static_par0_go_out;
wire _guard5984 = _guard5982 & _guard5983;
wire _guard5985 = cond_wire24_out;
wire _guard5986 = early_reset_static_par0_go_out;
wire _guard5987 = _guard5985 & _guard5986;
wire _guard5988 = early_reset_static_par0_go_out;
wire _guard5989 = early_reset_static_par0_go_out;
wire _guard5990 = early_reset_static_par0_go_out;
wire _guard5991 = early_reset_static_par0_go_out;
wire _guard5992 = early_reset_static_par0_go_out;
wire _guard5993 = early_reset_static_par0_go_out;
wire _guard5994 = early_reset_static_par0_go_out;
wire _guard5995 = early_reset_static_par0_go_out;
wire _guard5996 = early_reset_static_par0_go_out;
wire _guard5997 = early_reset_static_par0_go_out;
wire _guard5998 = fsm0_out == 5'd0;
wire _guard5999 = early_reset_static_seq_go_out;
wire _guard6000 = _guard5998 & _guard5999;
wire _guard6001 = early_reset_static_par0_go_out;
wire _guard6002 = _guard6000 | _guard6001;
wire _guard6003 = early_reset_static_par0_go_out;
wire _guard6004 = fsm0_out == 5'd0;
wire _guard6005 = early_reset_static_seq_go_out;
wire _guard6006 = _guard6004 & _guard6005;
wire _guard6007 = early_reset_static_par0_go_out;
wire _guard6008 = early_reset_static_par0_go_out;
wire _guard6009 = early_reset_static_par0_go_out;
wire _guard6010 = ~_guard0;
wire _guard6011 = early_reset_static_par0_go_out;
wire _guard6012 = _guard6010 & _guard6011;
wire _guard6013 = early_reset_static_par0_go_out;
wire _guard6014 = ~_guard0;
wire _guard6015 = early_reset_static_par0_go_out;
wire _guard6016 = _guard6014 & _guard6015;
wire _guard6017 = early_reset_static_par0_go_out;
wire _guard6018 = ~_guard0;
wire _guard6019 = early_reset_static_par0_go_out;
wire _guard6020 = _guard6018 & _guard6019;
wire _guard6021 = ~_guard0;
wire _guard6022 = early_reset_static_par0_go_out;
wire _guard6023 = _guard6021 & _guard6022;
wire _guard6024 = early_reset_static_par0_go_out;
wire _guard6025 = ~_guard0;
wire _guard6026 = early_reset_static_par0_go_out;
wire _guard6027 = _guard6025 & _guard6026;
wire _guard6028 = early_reset_static_par0_go_out;
wire _guard6029 = early_reset_static_par0_go_out;
wire _guard6030 = ~_guard0;
wire _guard6031 = early_reset_static_par0_go_out;
wire _guard6032 = _guard6030 & _guard6031;
wire _guard6033 = early_reset_static_par0_go_out;
wire _guard6034 = ~_guard0;
wire _guard6035 = early_reset_static_par0_go_out;
wire _guard6036 = _guard6034 & _guard6035;
wire _guard6037 = early_reset_static_par0_go_out;
wire _guard6038 = early_reset_static_par0_go_out;
wire _guard6039 = early_reset_static_par0_go_out;
wire _guard6040 = ~_guard0;
wire _guard6041 = early_reset_static_par0_go_out;
wire _guard6042 = _guard6040 & _guard6041;
wire _guard6043 = early_reset_static_par0_go_out;
wire _guard6044 = early_reset_static_par0_go_out;
wire _guard6045 = early_reset_static_par0_go_out;
wire _guard6046 = early_reset_static_par0_go_out;
wire _guard6047 = early_reset_static_par0_go_out;
wire _guard6048 = early_reset_static_par0_go_out;
wire _guard6049 = ~_guard0;
wire _guard6050 = early_reset_static_par0_go_out;
wire _guard6051 = _guard6049 & _guard6050;
wire _guard6052 = early_reset_static_par0_go_out;
wire _guard6053 = ~_guard0;
wire _guard6054 = early_reset_static_par0_go_out;
wire _guard6055 = _guard6053 & _guard6054;
wire _guard6056 = early_reset_static_par0_go_out;
wire _guard6057 = early_reset_static_par0_go_out;
wire _guard6058 = early_reset_static_par0_go_out;
wire _guard6059 = early_reset_static_par0_go_out;
wire _guard6060 = early_reset_static_par0_go_out;
wire _guard6061 = ~_guard0;
wire _guard6062 = early_reset_static_par0_go_out;
wire _guard6063 = _guard6061 & _guard6062;
wire _guard6064 = early_reset_static_par0_go_out;
wire _guard6065 = early_reset_static_par0_go_out;
wire _guard6066 = early_reset_static_par0_go_out;
wire _guard6067 = early_reset_static_par0_go_out;
wire _guard6068 = ~_guard0;
wire _guard6069 = early_reset_static_par0_go_out;
wire _guard6070 = _guard6068 & _guard6069;
wire _guard6071 = early_reset_static_par0_go_out;
wire _guard6072 = early_reset_static_par0_go_out;
wire _guard6073 = early_reset_static_par0_go_out;
wire _guard6074 = ~_guard0;
wire _guard6075 = early_reset_static_par0_go_out;
wire _guard6076 = _guard6074 & _guard6075;
wire _guard6077 = early_reset_static_par0_go_out;
wire _guard6078 = early_reset_static_par0_go_out;
wire _guard6079 = early_reset_static_par0_go_out;
wire _guard6080 = early_reset_static_par0_go_out;
wire _guard6081 = ~_guard0;
wire _guard6082 = early_reset_static_par0_go_out;
wire _guard6083 = _guard6081 & _guard6082;
wire _guard6084 = early_reset_static_par0_go_out;
wire _guard6085 = early_reset_static_par0_go_out;
wire _guard6086 = ~_guard0;
wire _guard6087 = early_reset_static_par0_go_out;
wire _guard6088 = _guard6086 & _guard6087;
wire _guard6089 = early_reset_static_par0_go_out;
wire _guard6090 = early_reset_static_par0_go_out;
wire _guard6091 = ~_guard0;
wire _guard6092 = early_reset_static_par0_go_out;
wire _guard6093 = _guard6091 & _guard6092;
wire _guard6094 = early_reset_static_par0_go_out;
wire _guard6095 = early_reset_static_par0_go_out;
wire _guard6096 = ~_guard0;
wire _guard6097 = early_reset_static_par0_go_out;
wire _guard6098 = _guard6096 & _guard6097;
wire _guard6099 = early_reset_static_par0_go_out;
wire _guard6100 = ~_guard0;
wire _guard6101 = early_reset_static_par0_go_out;
wire _guard6102 = _guard6100 & _guard6101;
wire _guard6103 = early_reset_static_par0_go_out;
wire _guard6104 = early_reset_static_par0_go_out;
wire _guard6105 = early_reset_static_par0_go_out;
wire _guard6106 = early_reset_static_par0_go_out;
wire _guard6107 = early_reset_static_par0_go_out;
wire _guard6108 = early_reset_static_par0_go_out;
wire _guard6109 = ~_guard0;
wire _guard6110 = early_reset_static_par0_go_out;
wire _guard6111 = _guard6109 & _guard6110;
wire _guard6112 = early_reset_static_par0_go_out;
wire _guard6113 = early_reset_static_par0_go_out;
wire _guard6114 = ~_guard0;
wire _guard6115 = early_reset_static_par0_go_out;
wire _guard6116 = _guard6114 & _guard6115;
wire _guard6117 = cond_wire14_out;
wire _guard6118 = early_reset_static_par0_go_out;
wire _guard6119 = _guard6117 & _guard6118;
wire _guard6120 = cond_wire14_out;
wire _guard6121 = early_reset_static_par0_go_out;
wire _guard6122 = _guard6120 & _guard6121;
wire _guard6123 = cond_wire32_out;
wire _guard6124 = early_reset_static_par0_go_out;
wire _guard6125 = _guard6123 & _guard6124;
wire _guard6126 = cond_wire30_out;
wire _guard6127 = early_reset_static_par0_go_out;
wire _guard6128 = _guard6126 & _guard6127;
wire _guard6129 = fsm_out == 1'd0;
wire _guard6130 = cond_wire30_out;
wire _guard6131 = _guard6129 & _guard6130;
wire _guard6132 = fsm_out == 1'd0;
wire _guard6133 = _guard6131 & _guard6132;
wire _guard6134 = fsm_out == 1'd0;
wire _guard6135 = cond_wire32_out;
wire _guard6136 = _guard6134 & _guard6135;
wire _guard6137 = fsm_out == 1'd0;
wire _guard6138 = _guard6136 & _guard6137;
wire _guard6139 = _guard6133 | _guard6138;
wire _guard6140 = early_reset_static_par0_go_out;
wire _guard6141 = _guard6139 & _guard6140;
wire _guard6142 = fsm_out == 1'd0;
wire _guard6143 = cond_wire30_out;
wire _guard6144 = _guard6142 & _guard6143;
wire _guard6145 = fsm_out == 1'd0;
wire _guard6146 = _guard6144 & _guard6145;
wire _guard6147 = fsm_out == 1'd0;
wire _guard6148 = cond_wire32_out;
wire _guard6149 = _guard6147 & _guard6148;
wire _guard6150 = fsm_out == 1'd0;
wire _guard6151 = _guard6149 & _guard6150;
wire _guard6152 = _guard6146 | _guard6151;
wire _guard6153 = early_reset_static_par0_go_out;
wire _guard6154 = _guard6152 & _guard6153;
wire _guard6155 = fsm_out == 1'd0;
wire _guard6156 = cond_wire30_out;
wire _guard6157 = _guard6155 & _guard6156;
wire _guard6158 = fsm_out == 1'd0;
wire _guard6159 = _guard6157 & _guard6158;
wire _guard6160 = fsm_out == 1'd0;
wire _guard6161 = cond_wire32_out;
wire _guard6162 = _guard6160 & _guard6161;
wire _guard6163 = fsm_out == 1'd0;
wire _guard6164 = _guard6162 & _guard6163;
wire _guard6165 = _guard6159 | _guard6164;
wire _guard6166 = early_reset_static_par0_go_out;
wire _guard6167 = _guard6165 & _guard6166;
wire _guard6168 = cond_wire36_out;
wire _guard6169 = early_reset_static_par0_go_out;
wire _guard6170 = _guard6168 & _guard6169;
wire _guard6171 = cond_wire36_out;
wire _guard6172 = early_reset_static_par0_go_out;
wire _guard6173 = _guard6171 & _guard6172;
wire _guard6174 = cond_wire45_out;
wire _guard6175 = early_reset_static_par0_go_out;
wire _guard6176 = _guard6174 & _guard6175;
wire _guard6177 = cond_wire45_out;
wire _guard6178 = early_reset_static_par0_go_out;
wire _guard6179 = _guard6177 & _guard6178;
wire _guard6180 = cond_wire115_out;
wire _guard6181 = early_reset_static_par0_go_out;
wire _guard6182 = _guard6180 & _guard6181;
wire _guard6183 = cond_wire115_out;
wire _guard6184 = early_reset_static_par0_go_out;
wire _guard6185 = _guard6183 & _guard6184;
wire _guard6186 = cond_wire102_out;
wire _guard6187 = early_reset_static_par0_go_out;
wire _guard6188 = _guard6186 & _guard6187;
wire _guard6189 = cond_wire102_out;
wire _guard6190 = early_reset_static_par0_go_out;
wire _guard6191 = _guard6189 & _guard6190;
wire _guard6192 = cond_wire140_out;
wire _guard6193 = early_reset_static_par0_go_out;
wire _guard6194 = _guard6192 & _guard6193;
wire _guard6195 = cond_wire140_out;
wire _guard6196 = early_reset_static_par0_go_out;
wire _guard6197 = _guard6195 & _guard6196;
wire _guard6198 = cond_wire153_out;
wire _guard6199 = early_reset_static_par0_go_out;
wire _guard6200 = _guard6198 & _guard6199;
wire _guard6201 = cond_wire151_out;
wire _guard6202 = early_reset_static_par0_go_out;
wire _guard6203 = _guard6201 & _guard6202;
wire _guard6204 = fsm_out == 1'd0;
wire _guard6205 = cond_wire151_out;
wire _guard6206 = _guard6204 & _guard6205;
wire _guard6207 = fsm_out == 1'd0;
wire _guard6208 = _guard6206 & _guard6207;
wire _guard6209 = fsm_out == 1'd0;
wire _guard6210 = cond_wire153_out;
wire _guard6211 = _guard6209 & _guard6210;
wire _guard6212 = fsm_out == 1'd0;
wire _guard6213 = _guard6211 & _guard6212;
wire _guard6214 = _guard6208 | _guard6213;
wire _guard6215 = early_reset_static_par0_go_out;
wire _guard6216 = _guard6214 & _guard6215;
wire _guard6217 = fsm_out == 1'd0;
wire _guard6218 = cond_wire151_out;
wire _guard6219 = _guard6217 & _guard6218;
wire _guard6220 = fsm_out == 1'd0;
wire _guard6221 = _guard6219 & _guard6220;
wire _guard6222 = fsm_out == 1'd0;
wire _guard6223 = cond_wire153_out;
wire _guard6224 = _guard6222 & _guard6223;
wire _guard6225 = fsm_out == 1'd0;
wire _guard6226 = _guard6224 & _guard6225;
wire _guard6227 = _guard6221 | _guard6226;
wire _guard6228 = early_reset_static_par0_go_out;
wire _guard6229 = _guard6227 & _guard6228;
wire _guard6230 = fsm_out == 1'd0;
wire _guard6231 = cond_wire151_out;
wire _guard6232 = _guard6230 & _guard6231;
wire _guard6233 = fsm_out == 1'd0;
wire _guard6234 = _guard6232 & _guard6233;
wire _guard6235 = fsm_out == 1'd0;
wire _guard6236 = cond_wire153_out;
wire _guard6237 = _guard6235 & _guard6236;
wire _guard6238 = fsm_out == 1'd0;
wire _guard6239 = _guard6237 & _guard6238;
wire _guard6240 = _guard6234 | _guard6239;
wire _guard6241 = early_reset_static_par0_go_out;
wire _guard6242 = _guard6240 & _guard6241;
wire _guard6243 = cond_wire171_out;
wire _guard6244 = early_reset_static_par0_go_out;
wire _guard6245 = _guard6243 & _guard6244;
wire _guard6246 = cond_wire171_out;
wire _guard6247 = early_reset_static_par0_go_out;
wire _guard6248 = _guard6246 & _guard6247;
wire _guard6249 = cond_wire231_out;
wire _guard6250 = early_reset_static_par0_go_out;
wire _guard6251 = _guard6249 & _guard6250;
wire _guard6252 = cond_wire229_out;
wire _guard6253 = early_reset_static_par0_go_out;
wire _guard6254 = _guard6252 & _guard6253;
wire _guard6255 = fsm_out == 1'd0;
wire _guard6256 = cond_wire229_out;
wire _guard6257 = _guard6255 & _guard6256;
wire _guard6258 = fsm_out == 1'd0;
wire _guard6259 = _guard6257 & _guard6258;
wire _guard6260 = fsm_out == 1'd0;
wire _guard6261 = cond_wire231_out;
wire _guard6262 = _guard6260 & _guard6261;
wire _guard6263 = fsm_out == 1'd0;
wire _guard6264 = _guard6262 & _guard6263;
wire _guard6265 = _guard6259 | _guard6264;
wire _guard6266 = early_reset_static_par0_go_out;
wire _guard6267 = _guard6265 & _guard6266;
wire _guard6268 = fsm_out == 1'd0;
wire _guard6269 = cond_wire229_out;
wire _guard6270 = _guard6268 & _guard6269;
wire _guard6271 = fsm_out == 1'd0;
wire _guard6272 = _guard6270 & _guard6271;
wire _guard6273 = fsm_out == 1'd0;
wire _guard6274 = cond_wire231_out;
wire _guard6275 = _guard6273 & _guard6274;
wire _guard6276 = fsm_out == 1'd0;
wire _guard6277 = _guard6275 & _guard6276;
wire _guard6278 = _guard6272 | _guard6277;
wire _guard6279 = early_reset_static_par0_go_out;
wire _guard6280 = _guard6278 & _guard6279;
wire _guard6281 = fsm_out == 1'd0;
wire _guard6282 = cond_wire229_out;
wire _guard6283 = _guard6281 & _guard6282;
wire _guard6284 = fsm_out == 1'd0;
wire _guard6285 = _guard6283 & _guard6284;
wire _guard6286 = fsm_out == 1'd0;
wire _guard6287 = cond_wire231_out;
wire _guard6288 = _guard6286 & _guard6287;
wire _guard6289 = fsm_out == 1'd0;
wire _guard6290 = _guard6288 & _guard6289;
wire _guard6291 = _guard6285 | _guard6290;
wire _guard6292 = early_reset_static_par0_go_out;
wire _guard6293 = _guard6291 & _guard6292;
wire _guard6294 = cond_wire248_out;
wire _guard6295 = early_reset_static_par0_go_out;
wire _guard6296 = _guard6294 & _guard6295;
wire _guard6297 = cond_wire246_out;
wire _guard6298 = early_reset_static_par0_go_out;
wire _guard6299 = _guard6297 & _guard6298;
wire _guard6300 = fsm_out == 1'd0;
wire _guard6301 = cond_wire246_out;
wire _guard6302 = _guard6300 & _guard6301;
wire _guard6303 = fsm_out == 1'd0;
wire _guard6304 = _guard6302 & _guard6303;
wire _guard6305 = fsm_out == 1'd0;
wire _guard6306 = cond_wire248_out;
wire _guard6307 = _guard6305 & _guard6306;
wire _guard6308 = fsm_out == 1'd0;
wire _guard6309 = _guard6307 & _guard6308;
wire _guard6310 = _guard6304 | _guard6309;
wire _guard6311 = early_reset_static_par0_go_out;
wire _guard6312 = _guard6310 & _guard6311;
wire _guard6313 = fsm_out == 1'd0;
wire _guard6314 = cond_wire246_out;
wire _guard6315 = _guard6313 & _guard6314;
wire _guard6316 = fsm_out == 1'd0;
wire _guard6317 = _guard6315 & _guard6316;
wire _guard6318 = fsm_out == 1'd0;
wire _guard6319 = cond_wire248_out;
wire _guard6320 = _guard6318 & _guard6319;
wire _guard6321 = fsm_out == 1'd0;
wire _guard6322 = _guard6320 & _guard6321;
wire _guard6323 = _guard6317 | _guard6322;
wire _guard6324 = early_reset_static_par0_go_out;
wire _guard6325 = _guard6323 & _guard6324;
wire _guard6326 = fsm_out == 1'd0;
wire _guard6327 = cond_wire246_out;
wire _guard6328 = _guard6326 & _guard6327;
wire _guard6329 = fsm_out == 1'd0;
wire _guard6330 = _guard6328 & _guard6329;
wire _guard6331 = fsm_out == 1'd0;
wire _guard6332 = cond_wire248_out;
wire _guard6333 = _guard6331 & _guard6332;
wire _guard6334 = fsm_out == 1'd0;
wire _guard6335 = _guard6333 & _guard6334;
wire _guard6336 = _guard6330 | _guard6335;
wire _guard6337 = early_reset_static_par0_go_out;
wire _guard6338 = _guard6336 & _guard6337;
wire _guard6339 = cond_wire267_out;
wire _guard6340 = early_reset_static_par0_go_out;
wire _guard6341 = _guard6339 & _guard6340;
wire _guard6342 = cond_wire266_out;
wire _guard6343 = early_reset_static_par0_go_out;
wire _guard6344 = _guard6342 & _guard6343;
wire _guard6345 = fsm_out == 1'd0;
wire _guard6346 = cond_wire266_out;
wire _guard6347 = _guard6345 & _guard6346;
wire _guard6348 = fsm_out == 1'd0;
wire _guard6349 = _guard6347 & _guard6348;
wire _guard6350 = fsm_out == 1'd0;
wire _guard6351 = cond_wire267_out;
wire _guard6352 = _guard6350 & _guard6351;
wire _guard6353 = fsm_out == 1'd0;
wire _guard6354 = _guard6352 & _guard6353;
wire _guard6355 = _guard6349 | _guard6354;
wire _guard6356 = early_reset_static_par0_go_out;
wire _guard6357 = _guard6355 & _guard6356;
wire _guard6358 = fsm_out == 1'd0;
wire _guard6359 = cond_wire266_out;
wire _guard6360 = _guard6358 & _guard6359;
wire _guard6361 = fsm_out == 1'd0;
wire _guard6362 = _guard6360 & _guard6361;
wire _guard6363 = fsm_out == 1'd0;
wire _guard6364 = cond_wire267_out;
wire _guard6365 = _guard6363 & _guard6364;
wire _guard6366 = fsm_out == 1'd0;
wire _guard6367 = _guard6365 & _guard6366;
wire _guard6368 = _guard6362 | _guard6367;
wire _guard6369 = early_reset_static_par0_go_out;
wire _guard6370 = _guard6368 & _guard6369;
wire _guard6371 = fsm_out == 1'd0;
wire _guard6372 = cond_wire266_out;
wire _guard6373 = _guard6371 & _guard6372;
wire _guard6374 = fsm_out == 1'd0;
wire _guard6375 = _guard6373 & _guard6374;
wire _guard6376 = fsm_out == 1'd0;
wire _guard6377 = cond_wire267_out;
wire _guard6378 = _guard6376 & _guard6377;
wire _guard6379 = fsm_out == 1'd0;
wire _guard6380 = _guard6378 & _guard6379;
wire _guard6381 = _guard6375 | _guard6380;
wire _guard6382 = early_reset_static_par0_go_out;
wire _guard6383 = _guard6381 & _guard6382;
wire _guard6384 = fsm0_out == 5'd0;
wire _guard6385 = early_reset_static_seq_go_out;
wire _guard6386 = _guard6384 & _guard6385;
wire _guard6387 = cond_wire9_out;
wire _guard6388 = early_reset_static_par0_go_out;
wire _guard6389 = _guard6387 & _guard6388;
wire _guard6390 = _guard6386 | _guard6389;
wire _guard6391 = fsm0_out == 5'd0;
wire _guard6392 = early_reset_static_seq_go_out;
wire _guard6393 = _guard6391 & _guard6392;
wire _guard6394 = cond_wire9_out;
wire _guard6395 = early_reset_static_par0_go_out;
wire _guard6396 = _guard6394 & _guard6395;
wire _guard6397 = fsm0_out == 5'd0;
wire _guard6398 = early_reset_static_seq_go_out;
wire _guard6399 = _guard6397 & _guard6398;
wire _guard6400 = cond_wire72_out;
wire _guard6401 = early_reset_static_par0_go_out;
wire _guard6402 = _guard6400 & _guard6401;
wire _guard6403 = _guard6399 | _guard6402;
wire _guard6404 = fsm0_out == 5'd0;
wire _guard6405 = early_reset_static_seq_go_out;
wire _guard6406 = _guard6404 & _guard6405;
wire _guard6407 = cond_wire72_out;
wire _guard6408 = early_reset_static_par0_go_out;
wire _guard6409 = _guard6407 & _guard6408;
wire _guard6410 = fsm0_out == 5'd0;
wire _guard6411 = early_reset_static_seq_go_out;
wire _guard6412 = _guard6410 & _guard6411;
wire _guard6413 = cond_wire204_out;
wire _guard6414 = early_reset_static_par0_go_out;
wire _guard6415 = _guard6413 & _guard6414;
wire _guard6416 = _guard6412 | _guard6415;
wire _guard6417 = fsm0_out == 5'd0;
wire _guard6418 = early_reset_static_seq_go_out;
wire _guard6419 = _guard6417 & _guard6418;
wire _guard6420 = cond_wire204_out;
wire _guard6421 = early_reset_static_par0_go_out;
wire _guard6422 = _guard6420 & _guard6421;
wire _guard6423 = early_reset_static_par0_go_out;
wire _guard6424 = early_reset_static_par0_go_out;
wire _guard6425 = early_reset_static_par0_go_out;
wire _guard6426 = early_reset_static_par0_go_out;
wire _guard6427 = fsm0_out == 5'd0;
wire _guard6428 = early_reset_static_seq_go_out;
wire _guard6429 = _guard6427 & _guard6428;
wire _guard6430 = early_reset_static_par0_go_out;
wire _guard6431 = _guard6429 | _guard6430;
wire _guard6432 = early_reset_static_par0_go_out;
wire _guard6433 = fsm0_out == 5'd0;
wire _guard6434 = early_reset_static_seq_go_out;
wire _guard6435 = _guard6433 & _guard6434;
wire _guard6436 = early_reset_static_par0_go_out;
wire _guard6437 = early_reset_static_par0_go_out;
wire _guard6438 = early_reset_static_par0_go_out;
wire _guard6439 = early_reset_static_par0_go_out;
wire _guard6440 = early_reset_static_par0_go_out;
wire _guard6441 = early_reset_static_par0_go_out;
wire _guard6442 = fsm0_out == 5'd0;
wire _guard6443 = early_reset_static_seq_go_out;
wire _guard6444 = _guard6442 & _guard6443;
wire _guard6445 = early_reset_static_par0_go_out;
wire _guard6446 = _guard6444 | _guard6445;
wire _guard6447 = fsm0_out == 5'd0;
wire _guard6448 = early_reset_static_seq_go_out;
wire _guard6449 = _guard6447 & _guard6448;
wire _guard6450 = early_reset_static_par0_go_out;
wire _guard6451 = early_reset_static_par0_go_out;
wire _guard6452 = early_reset_static_par0_go_out;
wire _guard6453 = early_reset_static_par0_go_out;
wire _guard6454 = early_reset_static_par0_go_out;
wire _guard6455 = fsm0_out == 5'd0;
wire _guard6456 = early_reset_static_seq_go_out;
wire _guard6457 = _guard6455 & _guard6456;
wire _guard6458 = early_reset_static_par0_go_out;
wire _guard6459 = _guard6457 | _guard6458;
wire _guard6460 = fsm0_out == 5'd0;
wire _guard6461 = early_reset_static_seq_go_out;
wire _guard6462 = _guard6460 & _guard6461;
wire _guard6463 = early_reset_static_par0_go_out;
wire _guard6464 = fsm0_out == 5'd0;
wire _guard6465 = early_reset_static_seq_go_out;
wire _guard6466 = _guard6464 & _guard6465;
wire _guard6467 = early_reset_static_par0_go_out;
wire _guard6468 = _guard6466 | _guard6467;
wire _guard6469 = early_reset_static_par0_go_out;
wire _guard6470 = fsm0_out == 5'd0;
wire _guard6471 = early_reset_static_seq_go_out;
wire _guard6472 = _guard6470 & _guard6471;
wire _guard6473 = early_reset_static_par0_go_out;
wire _guard6474 = early_reset_static_par0_go_out;
wire _guard6475 = early_reset_static_par0_go_out;
wire _guard6476 = early_reset_static_par0_go_out;
wire _guard6477 = ~_guard0;
wire _guard6478 = early_reset_static_par0_go_out;
wire _guard6479 = _guard6477 & _guard6478;
wire _guard6480 = early_reset_static_par0_go_out;
wire _guard6481 = early_reset_static_par0_go_out;
wire _guard6482 = early_reset_static_par0_go_out;
wire _guard6483 = early_reset_static_par0_go_out;
wire _guard6484 = early_reset_static_par0_go_out;
wire _guard6485 = early_reset_static_par0_go_out;
wire _guard6486 = ~_guard0;
wire _guard6487 = early_reset_static_par0_go_out;
wire _guard6488 = _guard6486 & _guard6487;
wire _guard6489 = early_reset_static_par0_go_out;
wire _guard6490 = early_reset_static_par0_go_out;
wire _guard6491 = early_reset_static_par0_go_out;
wire _guard6492 = early_reset_static_par0_go_out;
wire _guard6493 = ~_guard0;
wire _guard6494 = early_reset_static_par0_go_out;
wire _guard6495 = _guard6493 & _guard6494;
wire _guard6496 = early_reset_static_par0_go_out;
wire _guard6497 = ~_guard0;
wire _guard6498 = early_reset_static_par0_go_out;
wire _guard6499 = _guard6497 & _guard6498;
wire _guard6500 = early_reset_static_par0_go_out;
wire _guard6501 = ~_guard0;
wire _guard6502 = early_reset_static_par0_go_out;
wire _guard6503 = _guard6501 & _guard6502;
wire _guard6504 = early_reset_static_par0_go_out;
wire _guard6505 = ~_guard0;
wire _guard6506 = early_reset_static_par0_go_out;
wire _guard6507 = _guard6505 & _guard6506;
wire _guard6508 = early_reset_static_par0_go_out;
wire _guard6509 = early_reset_static_par0_go_out;
wire _guard6510 = early_reset_static_par0_go_out;
wire _guard6511 = early_reset_static_par0_go_out;
wire _guard6512 = early_reset_static_par0_go_out;
wire _guard6513 = ~_guard0;
wire _guard6514 = early_reset_static_par0_go_out;
wire _guard6515 = _guard6513 & _guard6514;
wire _guard6516 = early_reset_static_par0_go_out;
wire _guard6517 = early_reset_static_par0_go_out;
wire _guard6518 = early_reset_static_par0_go_out;
wire _guard6519 = early_reset_static_par0_go_out;
wire _guard6520 = early_reset_static_par0_go_out;
wire _guard6521 = early_reset_static_par0_go_out;
wire _guard6522 = early_reset_static_par0_go_out;
wire _guard6523 = early_reset_static_par0_go_out;
wire _guard6524 = early_reset_static_par0_go_out;
wire _guard6525 = early_reset_static_par0_go_out;
wire _guard6526 = early_reset_static_par0_go_out;
wire _guard6527 = early_reset_static_par0_go_out;
wire _guard6528 = early_reset_static_par0_go_out;
wire _guard6529 = early_reset_static_par0_go_out;
wire _guard6530 = ~_guard0;
wire _guard6531 = early_reset_static_par0_go_out;
wire _guard6532 = _guard6530 & _guard6531;
wire _guard6533 = early_reset_static_par0_go_out;
wire _guard6534 = early_reset_static_par0_go_out;
wire _guard6535 = early_reset_static_par0_go_out;
wire _guard6536 = early_reset_static_par0_go_out;
wire _guard6537 = ~_guard0;
wire _guard6538 = early_reset_static_par0_go_out;
wire _guard6539 = _guard6537 & _guard6538;
wire _guard6540 = early_reset_static_par0_go_out;
wire _guard6541 = early_reset_static_par0_go_out;
wire _guard6542 = early_reset_static_par0_go_out;
wire _guard6543 = early_reset_static_par0_go_out;
wire _guard6544 = early_reset_static_par0_go_out;
wire _guard6545 = early_reset_static_par0_go_out;
wire _guard6546 = early_reset_static_par0_go_out;
wire _guard6547 = early_reset_static_par0_go_out;
wire _guard6548 = ~_guard0;
wire _guard6549 = early_reset_static_par0_go_out;
wire _guard6550 = _guard6548 & _guard6549;
wire _guard6551 = ~_guard0;
wire _guard6552 = early_reset_static_par0_go_out;
wire _guard6553 = _guard6551 & _guard6552;
wire _guard6554 = early_reset_static_par0_go_out;
wire _guard6555 = early_reset_static_par0_go_out;
wire _guard6556 = early_reset_static_par0_go_out;
wire _guard6557 = early_reset_static_par0_go_out;
wire _guard6558 = ~_guard0;
wire _guard6559 = early_reset_static_par0_go_out;
wire _guard6560 = _guard6558 & _guard6559;
wire _guard6561 = early_reset_static_par0_go_out;
wire _guard6562 = early_reset_static_par0_go_out;
wire _guard6563 = early_reset_static_par0_go_out;
wire _guard6564 = ~_guard0;
wire _guard6565 = early_reset_static_par0_go_out;
wire _guard6566 = _guard6564 & _guard6565;
wire _guard6567 = early_reset_static_par0_go_out;
wire _guard6568 = ~_guard0;
wire _guard6569 = early_reset_static_par0_go_out;
wire _guard6570 = _guard6568 & _guard6569;
wire _guard6571 = ~_guard0;
wire _guard6572 = early_reset_static_par0_go_out;
wire _guard6573 = _guard6571 & _guard6572;
wire _guard6574 = early_reset_static_par0_go_out;
wire _guard6575 = early_reset_static_par0_go_out;
wire _guard6576 = early_reset_static_par0_go_out;
wire _guard6577 = early_reset_static_par0_go_out;
wire _guard6578 = ~_guard0;
wire _guard6579 = early_reset_static_par0_go_out;
wire _guard6580 = _guard6578 & _guard6579;
wire _guard6581 = early_reset_static_par0_go_out;
wire _guard6582 = early_reset_static_par0_go_out;
wire _guard6583 = cond_wire_out;
wire _guard6584 = early_reset_static_par0_go_out;
wire _guard6585 = _guard6583 & _guard6584;
wire _guard6586 = cond_wire_out;
wire _guard6587 = early_reset_static_par0_go_out;
wire _guard6588 = _guard6586 & _guard6587;
wire _guard6589 = cond_wire24_out;
wire _guard6590 = early_reset_static_par0_go_out;
wire _guard6591 = _guard6589 & _guard6590;
wire _guard6592 = cond_wire24_out;
wire _guard6593 = early_reset_static_par0_go_out;
wire _guard6594 = _guard6592 & _guard6593;
wire _guard6595 = cond_wire46_out;
wire _guard6596 = early_reset_static_par0_go_out;
wire _guard6597 = _guard6595 & _guard6596;
wire _guard6598 = cond_wire44_out;
wire _guard6599 = early_reset_static_par0_go_out;
wire _guard6600 = _guard6598 & _guard6599;
wire _guard6601 = fsm_out == 1'd0;
wire _guard6602 = cond_wire44_out;
wire _guard6603 = _guard6601 & _guard6602;
wire _guard6604 = fsm_out == 1'd0;
wire _guard6605 = _guard6603 & _guard6604;
wire _guard6606 = fsm_out == 1'd0;
wire _guard6607 = cond_wire46_out;
wire _guard6608 = _guard6606 & _guard6607;
wire _guard6609 = fsm_out == 1'd0;
wire _guard6610 = _guard6608 & _guard6609;
wire _guard6611 = _guard6605 | _guard6610;
wire _guard6612 = early_reset_static_par0_go_out;
wire _guard6613 = _guard6611 & _guard6612;
wire _guard6614 = fsm_out == 1'd0;
wire _guard6615 = cond_wire44_out;
wire _guard6616 = _guard6614 & _guard6615;
wire _guard6617 = fsm_out == 1'd0;
wire _guard6618 = _guard6616 & _guard6617;
wire _guard6619 = fsm_out == 1'd0;
wire _guard6620 = cond_wire46_out;
wire _guard6621 = _guard6619 & _guard6620;
wire _guard6622 = fsm_out == 1'd0;
wire _guard6623 = _guard6621 & _guard6622;
wire _guard6624 = _guard6618 | _guard6623;
wire _guard6625 = early_reset_static_par0_go_out;
wire _guard6626 = _guard6624 & _guard6625;
wire _guard6627 = fsm_out == 1'd0;
wire _guard6628 = cond_wire44_out;
wire _guard6629 = _guard6627 & _guard6628;
wire _guard6630 = fsm_out == 1'd0;
wire _guard6631 = _guard6629 & _guard6630;
wire _guard6632 = fsm_out == 1'd0;
wire _guard6633 = cond_wire46_out;
wire _guard6634 = _guard6632 & _guard6633;
wire _guard6635 = fsm_out == 1'd0;
wire _guard6636 = _guard6634 & _guard6635;
wire _guard6637 = _guard6631 | _guard6636;
wire _guard6638 = early_reset_static_par0_go_out;
wire _guard6639 = _guard6637 & _guard6638;
wire _guard6640 = cond_wire69_out;
wire _guard6641 = early_reset_static_par0_go_out;
wire _guard6642 = _guard6640 & _guard6641;
wire _guard6643 = cond_wire69_out;
wire _guard6644 = early_reset_static_par0_go_out;
wire _guard6645 = _guard6643 & _guard6644;
wire _guard6646 = cond_wire177_out;
wire _guard6647 = early_reset_static_par0_go_out;
wire _guard6648 = _guard6646 & _guard6647;
wire _guard6649 = cond_wire177_out;
wire _guard6650 = early_reset_static_par0_go_out;
wire _guard6651 = _guard6649 & _guard6650;
wire _guard6652 = cond_wire168_out;
wire _guard6653 = early_reset_static_par0_go_out;
wire _guard6654 = _guard6652 & _guard6653;
wire _guard6655 = cond_wire168_out;
wire _guard6656 = early_reset_static_par0_go_out;
wire _guard6657 = _guard6655 & _guard6656;
wire _guard6658 = cond_wire197_out;
wire _guard6659 = early_reset_static_par0_go_out;
wire _guard6660 = _guard6658 & _guard6659;
wire _guard6661 = cond_wire197_out;
wire _guard6662 = early_reset_static_par0_go_out;
wire _guard6663 = _guard6661 & _guard6662;
wire _guard6664 = cond_wire204_out;
wire _guard6665 = early_reset_static_par0_go_out;
wire _guard6666 = _guard6664 & _guard6665;
wire _guard6667 = cond_wire204_out;
wire _guard6668 = early_reset_static_par0_go_out;
wire _guard6669 = _guard6667 & _guard6668;
wire _guard6670 = cond_wire210_out;
wire _guard6671 = early_reset_static_par0_go_out;
wire _guard6672 = _guard6670 & _guard6671;
wire _guard6673 = cond_wire210_out;
wire _guard6674 = early_reset_static_par0_go_out;
wire _guard6675 = _guard6673 & _guard6674;
wire _guard6676 = early_reset_static_par0_go_out;
wire _guard6677 = early_reset_static_par0_go_out;
wire _guard6678 = fsm0_out == 5'd0;
wire _guard6679 = early_reset_static_seq_go_out;
wire _guard6680 = _guard6678 & _guard6679;
wire _guard6681 = early_reset_static_par0_go_out;
wire _guard6682 = _guard6680 | _guard6681;
wire _guard6683 = early_reset_static_par0_go_out;
wire _guard6684 = fsm0_out == 5'd0;
wire _guard6685 = early_reset_static_seq_go_out;
wire _guard6686 = _guard6684 & _guard6685;
wire _guard6687 = early_reset_static_par0_go_out;
wire _guard6688 = early_reset_static_par0_go_out;
wire _guard6689 = early_reset_static_par0_go_out;
wire _guard6690 = early_reset_static_par0_go_out;
wire _guard6691 = early_reset_static_par0_go_out;
wire _guard6692 = early_reset_static_par0_go_out;
wire _guard6693 = fsm0_out == 5'd0;
wire _guard6694 = early_reset_static_seq_go_out;
wire _guard6695 = _guard6693 & _guard6694;
wire _guard6696 = early_reset_static_par0_go_out;
wire _guard6697 = _guard6695 | _guard6696;
wire _guard6698 = early_reset_static_par0_go_out;
wire _guard6699 = fsm0_out == 5'd0;
wire _guard6700 = early_reset_static_seq_go_out;
wire _guard6701 = _guard6699 & _guard6700;
wire _guard6702 = early_reset_static_par0_go_out;
wire _guard6703 = early_reset_static_par0_go_out;
wire _guard6704 = fsm0_out == 5'd0;
wire _guard6705 = early_reset_static_seq_go_out;
wire _guard6706 = _guard6704 & _guard6705;
wire _guard6707 = early_reset_static_par0_go_out;
wire _guard6708 = _guard6706 | _guard6707;
wire _guard6709 = early_reset_static_par0_go_out;
wire _guard6710 = fsm0_out == 5'd0;
wire _guard6711 = early_reset_static_seq_go_out;
wire _guard6712 = _guard6710 & _guard6711;
wire _guard6713 = fsm0_out == 5'd0;
wire _guard6714 = early_reset_static_seq_go_out;
wire _guard6715 = _guard6713 & _guard6714;
wire _guard6716 = early_reset_static_par0_go_out;
wire _guard6717 = _guard6715 | _guard6716;
wire _guard6718 = early_reset_static_par0_go_out;
wire _guard6719 = fsm0_out == 5'd0;
wire _guard6720 = early_reset_static_seq_go_out;
wire _guard6721 = _guard6719 & _guard6720;
wire _guard6722 = fsm0_out == 5'd0;
wire _guard6723 = early_reset_static_seq_go_out;
wire _guard6724 = _guard6722 & _guard6723;
wire _guard6725 = early_reset_static_par0_go_out;
wire _guard6726 = _guard6724 | _guard6725;
wire _guard6727 = fsm0_out == 5'd0;
wire _guard6728 = early_reset_static_seq_go_out;
wire _guard6729 = _guard6727 & _guard6728;
wire _guard6730 = early_reset_static_par0_go_out;
wire _guard6731 = ~_guard0;
wire _guard6732 = early_reset_static_par0_go_out;
wire _guard6733 = _guard6731 & _guard6732;
wire _guard6734 = early_reset_static_par0_go_out;
wire _guard6735 = early_reset_static_par0_go_out;
wire _guard6736 = early_reset_static_par0_go_out;
wire _guard6737 = early_reset_static_par0_go_out;
wire _guard6738 = early_reset_static_par0_go_out;
wire _guard6739 = early_reset_static_par0_go_out;
wire _guard6740 = early_reset_static_par0_go_out;
wire _guard6741 = early_reset_static_par0_go_out;
wire _guard6742 = ~_guard0;
wire _guard6743 = early_reset_static_par0_go_out;
wire _guard6744 = _guard6742 & _guard6743;
wire _guard6745 = ~_guard0;
wire _guard6746 = early_reset_static_par0_go_out;
wire _guard6747 = _guard6745 & _guard6746;
wire _guard6748 = early_reset_static_par0_go_out;
wire _guard6749 = early_reset_static_par0_go_out;
wire _guard6750 = early_reset_static_par0_go_out;
wire _guard6751 = ~_guard0;
wire _guard6752 = early_reset_static_par0_go_out;
wire _guard6753 = _guard6751 & _guard6752;
wire _guard6754 = early_reset_static_par0_go_out;
wire _guard6755 = early_reset_static_par0_go_out;
wire _guard6756 = early_reset_static_par0_go_out;
wire _guard6757 = early_reset_static_par0_go_out;
wire _guard6758 = ~_guard0;
wire _guard6759 = early_reset_static_par0_go_out;
wire _guard6760 = _guard6758 & _guard6759;
wire _guard6761 = ~_guard0;
wire _guard6762 = early_reset_static_par0_go_out;
wire _guard6763 = _guard6761 & _guard6762;
wire _guard6764 = early_reset_static_par0_go_out;
wire _guard6765 = early_reset_static_par0_go_out;
wire _guard6766 = ~_guard0;
wire _guard6767 = early_reset_static_par0_go_out;
wire _guard6768 = _guard6766 & _guard6767;
wire _guard6769 = early_reset_static_par0_go_out;
wire _guard6770 = ~_guard0;
wire _guard6771 = early_reset_static_par0_go_out;
wire _guard6772 = _guard6770 & _guard6771;
wire _guard6773 = ~_guard0;
wire _guard6774 = early_reset_static_par0_go_out;
wire _guard6775 = _guard6773 & _guard6774;
wire _guard6776 = early_reset_static_par0_go_out;
wire _guard6777 = early_reset_static_par0_go_out;
wire _guard6778 = early_reset_static_par0_go_out;
wire _guard6779 = early_reset_static_par0_go_out;
wire _guard6780 = ~_guard0;
wire _guard6781 = early_reset_static_par0_go_out;
wire _guard6782 = _guard6780 & _guard6781;
wire _guard6783 = early_reset_static_par0_go_out;
wire _guard6784 = early_reset_static_par0_go_out;
wire _guard6785 = early_reset_static_par0_go_out;
wire _guard6786 = early_reset_static_par0_go_out;
wire _guard6787 = ~_guard0;
wire _guard6788 = early_reset_static_par0_go_out;
wire _guard6789 = _guard6787 & _guard6788;
wire _guard6790 = early_reset_static_par0_go_out;
wire _guard6791 = early_reset_static_par0_go_out;
wire _guard6792 = early_reset_static_par0_go_out;
wire _guard6793 = early_reset_static_par0_go_out;
wire _guard6794 = ~_guard0;
wire _guard6795 = early_reset_static_par0_go_out;
wire _guard6796 = _guard6794 & _guard6795;
wire _guard6797 = ~_guard0;
wire _guard6798 = early_reset_static_par0_go_out;
wire _guard6799 = _guard6797 & _guard6798;
wire _guard6800 = early_reset_static_par0_go_out;
wire _guard6801 = ~_guard0;
wire _guard6802 = early_reset_static_par0_go_out;
wire _guard6803 = _guard6801 & _guard6802;
wire _guard6804 = early_reset_static_par0_go_out;
wire _guard6805 = early_reset_static_par0_go_out;
wire _guard6806 = early_reset_static_par0_go_out;
wire _guard6807 = early_reset_static_par0_go_out;
wire _guard6808 = early_reset_static_par0_go_out;
wire _guard6809 = early_reset_static_par0_go_out;
wire _guard6810 = ~_guard0;
wire _guard6811 = early_reset_static_par0_go_out;
wire _guard6812 = _guard6810 & _guard6811;
wire _guard6813 = ~_guard0;
wire _guard6814 = early_reset_static_par0_go_out;
wire _guard6815 = _guard6813 & _guard6814;
wire _guard6816 = early_reset_static_par0_go_out;
wire _guard6817 = early_reset_static_par0_go_out;
wire _guard6818 = early_reset_static_par0_go_out;
wire _guard6819 = early_reset_static_par0_go_out;
wire _guard6820 = early_reset_static_par0_go_out;
wire _guard6821 = early_reset_static_par0_go_out;
wire _guard6822 = ~_guard0;
wire _guard6823 = early_reset_static_par0_go_out;
wire _guard6824 = _guard6822 & _guard6823;
wire _guard6825 = early_reset_static_par0_go_out;
wire _guard6826 = early_reset_static_par0_go_out;
wire _guard6827 = ~_guard0;
wire _guard6828 = early_reset_static_par0_go_out;
wire _guard6829 = _guard6827 & _guard6828;
wire _guard6830 = early_reset_static_par0_go_out;
wire _guard6831 = early_reset_static_par0_go_out;
wire _guard6832 = early_reset_static_par0_go_out;
wire _guard6833 = cond_wire1_out;
wire _guard6834 = early_reset_static_par0_go_out;
wire _guard6835 = _guard6833 & _guard6834;
wire _guard6836 = cond_wire1_out;
wire _guard6837 = early_reset_static_par0_go_out;
wire _guard6838 = _guard6836 & _guard6837;
wire _guard6839 = cond_wire34_out;
wire _guard6840 = early_reset_static_par0_go_out;
wire _guard6841 = _guard6839 & _guard6840;
wire _guard6842 = cond_wire34_out;
wire _guard6843 = early_reset_static_par0_go_out;
wire _guard6844 = _guard6842 & _guard6843;
wire _guard6845 = cond_wire65_out;
wire _guard6846 = early_reset_static_par0_go_out;
wire _guard6847 = _guard6845 & _guard6846;
wire _guard6848 = cond_wire65_out;
wire _guard6849 = early_reset_static_par0_go_out;
wire _guard6850 = _guard6848 & _guard6849;
wire _guard6851 = cond_wire83_out;
wire _guard6852 = early_reset_static_par0_go_out;
wire _guard6853 = _guard6851 & _guard6852;
wire _guard6854 = cond_wire81_out;
wire _guard6855 = early_reset_static_par0_go_out;
wire _guard6856 = _guard6854 & _guard6855;
wire _guard6857 = fsm_out == 1'd0;
wire _guard6858 = cond_wire81_out;
wire _guard6859 = _guard6857 & _guard6858;
wire _guard6860 = fsm_out == 1'd0;
wire _guard6861 = _guard6859 & _guard6860;
wire _guard6862 = fsm_out == 1'd0;
wire _guard6863 = cond_wire83_out;
wire _guard6864 = _guard6862 & _guard6863;
wire _guard6865 = fsm_out == 1'd0;
wire _guard6866 = _guard6864 & _guard6865;
wire _guard6867 = _guard6861 | _guard6866;
wire _guard6868 = early_reset_static_par0_go_out;
wire _guard6869 = _guard6867 & _guard6868;
wire _guard6870 = fsm_out == 1'd0;
wire _guard6871 = cond_wire81_out;
wire _guard6872 = _guard6870 & _guard6871;
wire _guard6873 = fsm_out == 1'd0;
wire _guard6874 = _guard6872 & _guard6873;
wire _guard6875 = fsm_out == 1'd0;
wire _guard6876 = cond_wire83_out;
wire _guard6877 = _guard6875 & _guard6876;
wire _guard6878 = fsm_out == 1'd0;
wire _guard6879 = _guard6877 & _guard6878;
wire _guard6880 = _guard6874 | _guard6879;
wire _guard6881 = early_reset_static_par0_go_out;
wire _guard6882 = _guard6880 & _guard6881;
wire _guard6883 = fsm_out == 1'd0;
wire _guard6884 = cond_wire81_out;
wire _guard6885 = _guard6883 & _guard6884;
wire _guard6886 = fsm_out == 1'd0;
wire _guard6887 = _guard6885 & _guard6886;
wire _guard6888 = fsm_out == 1'd0;
wire _guard6889 = cond_wire83_out;
wire _guard6890 = _guard6888 & _guard6889;
wire _guard6891 = fsm_out == 1'd0;
wire _guard6892 = _guard6890 & _guard6891;
wire _guard6893 = _guard6887 | _guard6892;
wire _guard6894 = early_reset_static_par0_go_out;
wire _guard6895 = _guard6893 & _guard6894;
wire _guard6896 = cond_wire145_out;
wire _guard6897 = early_reset_static_par0_go_out;
wire _guard6898 = _guard6896 & _guard6897;
wire _guard6899 = cond_wire143_out;
wire _guard6900 = early_reset_static_par0_go_out;
wire _guard6901 = _guard6899 & _guard6900;
wire _guard6902 = fsm_out == 1'd0;
wire _guard6903 = cond_wire143_out;
wire _guard6904 = _guard6902 & _guard6903;
wire _guard6905 = fsm_out == 1'd0;
wire _guard6906 = _guard6904 & _guard6905;
wire _guard6907 = fsm_out == 1'd0;
wire _guard6908 = cond_wire145_out;
wire _guard6909 = _guard6907 & _guard6908;
wire _guard6910 = fsm_out == 1'd0;
wire _guard6911 = _guard6909 & _guard6910;
wire _guard6912 = _guard6906 | _guard6911;
wire _guard6913 = early_reset_static_par0_go_out;
wire _guard6914 = _guard6912 & _guard6913;
wire _guard6915 = fsm_out == 1'd0;
wire _guard6916 = cond_wire143_out;
wire _guard6917 = _guard6915 & _guard6916;
wire _guard6918 = fsm_out == 1'd0;
wire _guard6919 = _guard6917 & _guard6918;
wire _guard6920 = fsm_out == 1'd0;
wire _guard6921 = cond_wire145_out;
wire _guard6922 = _guard6920 & _guard6921;
wire _guard6923 = fsm_out == 1'd0;
wire _guard6924 = _guard6922 & _guard6923;
wire _guard6925 = _guard6919 | _guard6924;
wire _guard6926 = early_reset_static_par0_go_out;
wire _guard6927 = _guard6925 & _guard6926;
wire _guard6928 = fsm_out == 1'd0;
wire _guard6929 = cond_wire143_out;
wire _guard6930 = _guard6928 & _guard6929;
wire _guard6931 = fsm_out == 1'd0;
wire _guard6932 = _guard6930 & _guard6931;
wire _guard6933 = fsm_out == 1'd0;
wire _guard6934 = cond_wire145_out;
wire _guard6935 = _guard6933 & _guard6934;
wire _guard6936 = fsm_out == 1'd0;
wire _guard6937 = _guard6935 & _guard6936;
wire _guard6938 = _guard6932 | _guard6937;
wire _guard6939 = early_reset_static_par0_go_out;
wire _guard6940 = _guard6938 & _guard6939;
wire _guard6941 = cond_wire148_out;
wire _guard6942 = early_reset_static_par0_go_out;
wire _guard6943 = _guard6941 & _guard6942;
wire _guard6944 = cond_wire148_out;
wire _guard6945 = early_reset_static_par0_go_out;
wire _guard6946 = _guard6944 & _guard6945;
wire _guard6947 = cond_wire214_out;
wire _guard6948 = early_reset_static_par0_go_out;
wire _guard6949 = _guard6947 & _guard6948;
wire _guard6950 = cond_wire214_out;
wire _guard6951 = early_reset_static_par0_go_out;
wire _guard6952 = _guard6950 & _guard6951;
wire _guard6953 = cond_wire72_out;
wire _guard6954 = early_reset_static_par0_go_out;
wire _guard6955 = _guard6953 & _guard6954;
wire _guard6956 = cond_wire72_out;
wire _guard6957 = early_reset_static_par0_go_out;
wire _guard6958 = _guard6956 & _guard6957;
wire _guard6959 = fsm0_out == 5'd0;
wire _guard6960 = early_reset_static_seq_go_out;
wire _guard6961 = _guard6959 & _guard6960;
wire _guard6962 = cond_wire171_out;
wire _guard6963 = early_reset_static_par0_go_out;
wire _guard6964 = _guard6962 & _guard6963;
wire _guard6965 = _guard6961 | _guard6964;
wire _guard6966 = fsm0_out == 5'd0;
wire _guard6967 = early_reset_static_seq_go_out;
wire _guard6968 = _guard6966 & _guard6967;
wire _guard6969 = cond_wire171_out;
wire _guard6970 = early_reset_static_par0_go_out;
wire _guard6971 = _guard6969 & _guard6970;
wire _guard6972 = cond_wire204_out;
wire _guard6973 = early_reset_static_par0_go_out;
wire _guard6974 = _guard6972 & _guard6973;
wire _guard6975 = cond_wire204_out;
wire _guard6976 = early_reset_static_par0_go_out;
wire _guard6977 = _guard6975 & _guard6976;
wire _guard6978 = early_reset_static_par0_go_out;
wire _guard6979 = early_reset_static_par0_go_out;
wire _guard6980 = early_reset_static_par0_go_out;
wire _guard6981 = early_reset_static_par0_go_out;
wire _guard6982 = fsm0_out == 5'd0;
wire _guard6983 = early_reset_static_seq_go_out;
wire _guard6984 = _guard6982 & _guard6983;
wire _guard6985 = early_reset_static_par0_go_out;
wire _guard6986 = _guard6984 | _guard6985;
wire _guard6987 = early_reset_static_par0_go_out;
wire _guard6988 = fsm0_out == 5'd0;
wire _guard6989 = early_reset_static_seq_go_out;
wire _guard6990 = _guard6988 & _guard6989;
wire _guard6991 = early_reset_static_par0_go_out;
wire _guard6992 = early_reset_static_par0_go_out;
wire _guard6993 = early_reset_static_par0_go_out;
wire _guard6994 = early_reset_static_par0_go_out;
wire _guard6995 = early_reset_static_par0_go_out;
wire _guard6996 = early_reset_static_par0_go_out;
wire _guard6997 = fsm0_out == 5'd0;
wire _guard6998 = early_reset_static_seq_go_out;
wire _guard6999 = _guard6997 & _guard6998;
wire _guard7000 = early_reset_static_par0_go_out;
wire _guard7001 = _guard6999 | _guard7000;
wire _guard7002 = early_reset_static_par0_go_out;
wire _guard7003 = fsm0_out == 5'd0;
wire _guard7004 = early_reset_static_seq_go_out;
wire _guard7005 = _guard7003 & _guard7004;
wire _guard7006 = fsm0_out == 5'd0;
wire _guard7007 = early_reset_static_seq_go_out;
wire _guard7008 = _guard7006 & _guard7007;
wire _guard7009 = early_reset_static_par0_go_out;
wire _guard7010 = _guard7008 | _guard7009;
wire _guard7011 = fsm0_out == 5'd0;
wire _guard7012 = early_reset_static_seq_go_out;
wire _guard7013 = _guard7011 & _guard7012;
wire _guard7014 = early_reset_static_par0_go_out;
wire _guard7015 = early_reset_static_par0_go_out;
wire _guard7016 = early_reset_static_par0_go_out;
wire _guard7017 = ~_guard0;
wire _guard7018 = early_reset_static_par0_go_out;
wire _guard7019 = _guard7017 & _guard7018;
wire _guard7020 = early_reset_static_par0_go_out;
wire _guard7021 = early_reset_static_par0_go_out;
wire _guard7022 = ~_guard0;
wire _guard7023 = early_reset_static_par0_go_out;
wire _guard7024 = _guard7022 & _guard7023;
wire _guard7025 = early_reset_static_par0_go_out;
wire _guard7026 = early_reset_static_par0_go_out;
wire _guard7027 = early_reset_static_par0_go_out;
wire _guard7028 = early_reset_static_par0_go_out;
wire _guard7029 = early_reset_static_par0_go_out;
wire _guard7030 = ~_guard0;
wire _guard7031 = early_reset_static_par0_go_out;
wire _guard7032 = _guard7030 & _guard7031;
wire _guard7033 = early_reset_static_par0_go_out;
wire _guard7034 = early_reset_static_par0_go_out;
wire _guard7035 = early_reset_static_par0_go_out;
wire _guard7036 = ~_guard0;
wire _guard7037 = early_reset_static_par0_go_out;
wire _guard7038 = _guard7036 & _guard7037;
wire _guard7039 = early_reset_static_par0_go_out;
wire _guard7040 = ~_guard0;
wire _guard7041 = early_reset_static_par0_go_out;
wire _guard7042 = _guard7040 & _guard7041;
wire _guard7043 = early_reset_static_par0_go_out;
wire _guard7044 = early_reset_static_par0_go_out;
wire _guard7045 = early_reset_static_par0_go_out;
wire _guard7046 = ~_guard0;
wire _guard7047 = early_reset_static_par0_go_out;
wire _guard7048 = _guard7046 & _guard7047;
wire _guard7049 = early_reset_static_par0_go_out;
wire _guard7050 = early_reset_static_par0_go_out;
wire _guard7051 = ~_guard0;
wire _guard7052 = early_reset_static_par0_go_out;
wire _guard7053 = _guard7051 & _guard7052;
wire _guard7054 = early_reset_static_par0_go_out;
wire _guard7055 = early_reset_static_par0_go_out;
wire _guard7056 = early_reset_static_par0_go_out;
wire _guard7057 = early_reset_static_par0_go_out;
wire _guard7058 = early_reset_static_par0_go_out;
wire _guard7059 = early_reset_static_par0_go_out;
wire _guard7060 = ~_guard0;
wire _guard7061 = early_reset_static_par0_go_out;
wire _guard7062 = _guard7060 & _guard7061;
wire _guard7063 = ~_guard0;
wire _guard7064 = early_reset_static_par0_go_out;
wire _guard7065 = _guard7063 & _guard7064;
wire _guard7066 = early_reset_static_par0_go_out;
wire _guard7067 = early_reset_static_par0_go_out;
wire _guard7068 = ~_guard0;
wire _guard7069 = early_reset_static_par0_go_out;
wire _guard7070 = _guard7068 & _guard7069;
wire _guard7071 = ~_guard0;
wire _guard7072 = early_reset_static_par0_go_out;
wire _guard7073 = _guard7071 & _guard7072;
wire _guard7074 = early_reset_static_par0_go_out;
wire _guard7075 = early_reset_static_par0_go_out;
wire _guard7076 = early_reset_static_par0_go_out;
wire _guard7077 = ~_guard0;
wire _guard7078 = early_reset_static_par0_go_out;
wire _guard7079 = _guard7077 & _guard7078;
wire _guard7080 = early_reset_static_par0_go_out;
wire _guard7081 = ~_guard0;
wire _guard7082 = early_reset_static_par0_go_out;
wire _guard7083 = _guard7081 & _guard7082;
wire _guard7084 = early_reset_static_par0_go_out;
wire _guard7085 = ~_guard0;
wire _guard7086 = early_reset_static_par0_go_out;
wire _guard7087 = _guard7085 & _guard7086;
wire _guard7088 = early_reset_static_par0_go_out;
wire _guard7089 = ~_guard0;
wire _guard7090 = early_reset_static_par0_go_out;
wire _guard7091 = _guard7089 & _guard7090;
wire _guard7092 = early_reset_static_par0_go_out;
wire _guard7093 = ~_guard0;
wire _guard7094 = early_reset_static_par0_go_out;
wire _guard7095 = _guard7093 & _guard7094;
wire _guard7096 = early_reset_static_par0_go_out;
wire _guard7097 = early_reset_static_par0_go_out;
wire _guard7098 = early_reset_static_par0_go_out;
wire _guard7099 = early_reset_static_par0_go_out;
wire _guard7100 = early_reset_static_par0_go_out;
wire _guard7101 = early_reset_static_par0_go_out;
wire _guard7102 = ~_guard0;
wire _guard7103 = early_reset_static_par0_go_out;
wire _guard7104 = _guard7102 & _guard7103;
assign pe_1_4_mul_ready =
  _guard3 ? 1'd1 :
  _guard6 ? 1'd0 :
  1'd0;
assign pe_1_4_clk = clk;
assign pe_1_4_top =
  _guard19 ? top_1_4_out :
  32'd0;
assign pe_1_4_left =
  _guard32 ? left_1_4_out :
  32'd0;
assign pe_1_4_reset = reset;
assign pe_1_4_go = _guard45;
assign pe_1_7_mul_ready =
  _guard48 ? 1'd1 :
  _guard51 ? 1'd0 :
  1'd0;
assign pe_1_7_clk = clk;
assign pe_1_7_top =
  _guard64 ? top_1_7_out :
  32'd0;
assign pe_1_7_left =
  _guard77 ? left_1_7_out :
  32'd0;
assign pe_1_7_reset = reset;
assign pe_1_7_go = _guard90;
assign top_2_4_write_en = _guard93;
assign top_2_4_clk = clk;
assign top_2_4_reset = reset;
assign top_2_4_in = top_1_4_out;
assign left_2_4_write_en = _guard99;
assign left_2_4_clk = clk;
assign left_2_4_reset = reset;
assign left_2_4_in = left_2_3_out;
assign top_3_5_write_en = _guard105;
assign top_3_5_clk = clk;
assign top_3_5_reset = reset;
assign top_3_5_in = top_2_5_out;
assign top_3_6_write_en = _guard111;
assign top_3_6_clk = clk;
assign top_3_6_reset = reset;
assign top_3_6_in = top_2_6_out;
assign left_4_0_write_en = _guard117;
assign left_4_0_clk = clk;
assign left_4_0_reset = reset;
assign left_4_0_in = l4_read_data;
assign top_4_4_write_en = _guard123;
assign top_4_4_clk = clk;
assign top_4_4_reset = reset;
assign top_4_4_in = top_3_4_out;
assign pe_5_2_mul_ready =
  _guard129 ? 1'd1 :
  _guard132 ? 1'd0 :
  1'd0;
assign pe_5_2_clk = clk;
assign pe_5_2_top =
  _guard145 ? top_5_2_out :
  32'd0;
assign pe_5_2_left =
  _guard158 ? left_5_2_out :
  32'd0;
assign pe_5_2_reset = reset;
assign pe_5_2_go = _guard171;
assign top_6_1_write_en = _guard174;
assign top_6_1_clk = clk;
assign top_6_1_reset = reset;
assign top_6_1_in = top_5_1_out;
assign left_6_2_write_en = _guard180;
assign left_6_2_clk = clk;
assign left_6_2_reset = reset;
assign left_6_2_in = left_6_1_out;
assign top_6_3_write_en = _guard186;
assign top_6_3_clk = clk;
assign top_6_3_reset = reset;
assign top_6_3_in = top_5_3_out;
assign left_6_4_write_en = _guard192;
assign left_6_4_clk = clk;
assign left_6_4_reset = reset;
assign left_6_4_in = left_6_3_out;
assign top_7_0_write_en = _guard198;
assign top_7_0_clk = clk;
assign top_7_0_reset = reset;
assign top_7_0_in = top_6_0_out;
assign t3_add_left = 4'd1;
assign t3_add_right = t3_idx_out;
assign l1_add_left = 4'd1;
assign l1_add_right = l1_idx_out;
assign idx_between_18_26_comb_left = index_ge_18_out;
assign idx_between_18_26_comb_right = index_lt_26_out;
assign idx_between_3_7_reg_write_en = _guard220;
assign idx_between_3_7_reg_clk = clk;
assign idx_between_3_7_reg_reset = reset;
assign idx_between_3_7_reg_in =
  _guard221 ? idx_between_3_7_comb_out :
  _guard224 ? 1'd0 :
  'x;
assign index_ge_15_left = idx_add_out;
assign index_ge_15_right = 5'd15;
assign index_lt_5_left = idx_add_out;
assign index_lt_5_right = 5'd5;
assign idx_between_11_19_reg_write_en = _guard233;
assign idx_between_11_19_reg_clk = clk;
assign idx_between_11_19_reg_reset = reset;
assign idx_between_11_19_reg_in =
  _guard236 ? 1'd0 :
  _guard237 ? idx_between_11_19_comb_out :
  'x;
assign idx_between_24_25_comb_left = index_ge_24_out;
assign idx_between_24_25_comb_right = index_lt_25_out;
assign idx_between_15_19_reg_write_en = _guard244;
assign idx_between_15_19_reg_clk = clk;
assign idx_between_15_19_reg_reset = reset;
assign idx_between_15_19_reg_in =
  _guard245 ? idx_between_15_19_comb_out :
  _guard248 ? 1'd0 :
  'x;
assign idx_between_8_16_comb_left = index_ge_8_out;
assign idx_between_8_16_comb_right = index_lt_16_out;
assign idx_between_17_25_comb_left = index_ge_17_out;
assign idx_between_17_25_comb_right = index_lt_25_out;
assign cond_wire3_in =
  _guard253 ? idx_between_13_14_reg_out :
  _guard256 ? cond3_out :
  1'd0;
assign cond_wire30_in =
  _guard259 ? cond30_out :
  _guard260 ? idx_between_7_11_reg_out :
  1'd0;
assign cond_wire38_in =
  _guard261 ? idx_between_20_21_reg_out :
  _guard264 ? cond38_out :
  1'd0;
assign cond_wire39_in =
  _guard267 ? cond39_out :
  _guard268 ? idx_between_1_9_reg_out :
  1'd0;
assign cond_wire47_in =
  _guard269 ? idx_between_15_16_reg_out :
  _guard272 ? cond47_out :
  1'd0;
assign cond53_write_en = _guard273;
assign cond53_clk = clk;
assign cond53_reset = reset;
assign cond53_in =
  _guard274 ? idx_between_5_13_reg_out :
  1'd0;
assign cond_wire54_in =
  _guard277 ? cond54_out :
  _guard278 ? idx_between_9_17_reg_out :
  1'd0;
assign cond65_write_en = _guard279;
assign cond65_clk = clk;
assign cond65_reset = reset;
assign cond65_in =
  _guard280 ? idx_between_8_16_reg_out :
  1'd0;
assign cond70_write_en = _guard281;
assign cond70_clk = clk;
assign cond70_reset = reset;
assign cond70_in =
  _guard282 ? idx_between_13_21_reg_out :
  1'd0;
assign cond71_write_en = _guard283;
assign cond71_clk = clk;
assign cond71_reset = reset;
assign cond71_in =
  _guard284 ? idx_between_21_22_reg_out :
  1'd0;
assign cond_wire89_in =
  _guard285 ? idx_between_7_11_reg_out :
  _guard288 ? cond89_out :
  1'd0;
assign cond_wire90_in =
  _guard289 ? idx_between_7_15_reg_out :
  _guard292 ? cond90_out :
  1'd0;
assign cond_wire103_in =
  _guard295 ? cond103_out :
  _guard296 ? idx_between_14_22_reg_out :
  1'd0;
assign cond_wire131_in =
  _guard299 ? cond131_out :
  _guard300 ? idx_between_10_18_reg_out :
  1'd0;
assign cond_wire164_in =
  _guard301 ? idx_between_11_19_reg_out :
  _guard304 ? cond164_out :
  1'd0;
assign cond167_write_en = _guard305;
assign cond167_clk = clk;
assign cond167_reset = reset;
assign cond167_in =
  _guard306 ? idx_between_12_16_reg_out :
  1'd0;
assign cond181_write_en = _guard307;
assign cond181_clk = clk;
assign cond181_reset = reset;
assign cond181_in =
  _guard308 ? idx_between_8_16_reg_out :
  1'd0;
assign cond_wire185_in =
  _guard311 ? cond185_out :
  _guard312 ? idx_between_9_17_reg_out :
  1'd0;
assign cond_wire193_in =
  _guard313 ? idx_between_11_19_reg_out :
  _guard316 ? cond193_out :
  1'd0;
assign cond202_write_en = _guard317;
assign cond202_clk = clk;
assign cond202_reset = reset;
assign cond202_in =
  _guard318 ? idx_between_17_25_reg_out :
  1'd0;
assign cond_wire204_in =
  _guard319 ? idx_between_6_14_reg_out :
  _guard322 ? cond204_out :
  1'd0;
assign cond_wire224_in =
  _guard323 ? idx_between_23_24_reg_out :
  _guard326 ? cond224_out :
  1'd0;
assign cond227_write_en = _guard327;
assign cond227_clk = clk;
assign cond227_reset = reset;
assign cond227_in =
  _guard328 ? idx_between_16_24_reg_out :
  1'd0;
assign cond230_write_en = _guard329;
assign cond230_clk = clk;
assign cond230_reset = reset;
assign cond230_in =
  _guard330 ? idx_between_13_21_reg_out :
  1'd0;
assign cond_wire234_in =
  _guard331 ? idx_between_14_22_reg_out :
  _guard334 ? cond234_out :
  1'd0;
assign cond239_write_en = _guard335;
assign cond239_clk = clk;
assign cond239_reset = reset;
assign cond239_in =
  _guard336 ? idx_between_8_16_reg_out :
  1'd0;
assign cond_wire240_in =
  _guard339 ? cond240_out :
  _guard340 ? idx_between_12_20_reg_out :
  1'd0;
assign cond263_write_en = _guard341;
assign cond263_clk = clk;
assign cond263_reset = reset;
assign cond263_in =
  _guard342 ? idx_between_14_22_reg_out :
  1'd0;
assign left_0_3_write_en = _guard345;
assign left_0_3_clk = clk;
assign left_0_3_reset = reset;
assign left_0_3_in = left_0_2_out;
assign left_0_4_write_en = _guard351;
assign left_0_4_clk = clk;
assign left_0_4_reset = reset;
assign left_0_4_in = left_0_3_out;
assign top_1_0_write_en = _guard357;
assign top_1_0_clk = clk;
assign top_1_0_reset = reset;
assign top_1_0_in = top_0_0_out;
assign pe_1_2_mul_ready =
  _guard363 ? 1'd1 :
  _guard366 ? 1'd0 :
  1'd0;
assign pe_1_2_clk = clk;
assign pe_1_2_top =
  _guard379 ? top_1_2_out :
  32'd0;
assign pe_1_2_left =
  _guard392 ? left_1_2_out :
  32'd0;
assign pe_1_2_reset = reset;
assign pe_1_2_go = _guard405;
assign pe_1_3_mul_ready =
  _guard408 ? 1'd1 :
  _guard411 ? 1'd0 :
  1'd0;
assign pe_1_3_clk = clk;
assign pe_1_3_top =
  _guard424 ? top_1_3_out :
  32'd0;
assign pe_1_3_left =
  _guard437 ? left_1_3_out :
  32'd0;
assign pe_1_3_reset = reset;
assign pe_1_3_go = _guard450;
assign left_1_3_write_en = _guard453;
assign left_1_3_clk = clk;
assign left_1_3_reset = reset;
assign left_1_3_in = left_1_2_out;
assign left_2_6_write_en = _guard459;
assign left_2_6_clk = clk;
assign left_2_6_reset = reset;
assign left_2_6_in = left_2_5_out;
assign top_4_7_write_en = _guard465;
assign top_4_7_clk = clk;
assign top_4_7_reset = reset;
assign top_4_7_in = top_3_7_out;
assign left_5_1_write_en = _guard471;
assign left_5_1_clk = clk;
assign left_5_1_reset = reset;
assign left_5_1_in = left_5_0_out;
assign left_5_3_write_en = _guard477;
assign left_5_3_clk = clk;
assign left_5_3_reset = reset;
assign left_5_3_in = left_5_2_out;
assign pe_6_4_mul_ready =
  _guard483 ? 1'd1 :
  _guard486 ? 1'd0 :
  1'd0;
assign pe_6_4_clk = clk;
assign pe_6_4_top =
  _guard499 ? top_6_4_out :
  32'd0;
assign pe_6_4_left =
  _guard512 ? left_6_4_out :
  32'd0;
assign pe_6_4_reset = reset;
assign pe_6_4_go = _guard525;
assign top_6_7_write_en = _guard528;
assign top_6_7_clk = clk;
assign top_6_7_reset = reset;
assign top_6_7_in = top_5_7_out;
assign pe_7_3_mul_ready =
  _guard534 ? 1'd1 :
  _guard537 ? 1'd0 :
  1'd0;
assign pe_7_3_clk = clk;
assign pe_7_3_top =
  _guard550 ? top_7_3_out :
  32'd0;
assign pe_7_3_left =
  _guard563 ? left_7_3_out :
  32'd0;
assign pe_7_3_reset = reset;
assign pe_7_3_go = _guard576;
assign left_7_4_write_en = _guard579;
assign left_7_4_clk = clk;
assign left_7_4_reset = reset;
assign left_7_4_in = left_7_3_out;
assign left_7_6_write_en = _guard585;
assign left_7_6_clk = clk;
assign left_7_6_reset = reset;
assign left_7_6_in = left_7_5_out;
assign top_7_7_write_en = _guard591;
assign top_7_7_clk = clk;
assign top_7_7_reset = reset;
assign top_7_7_in = top_6_7_out;
assign l3_idx_write_en = _guard601;
assign l3_idx_clk = clk;
assign l3_idx_reset = reset;
assign l3_idx_in =
  _guard604 ? l3_add_out :
  _guard607 ? 4'd0 :
  'x;
assign l7_idx_write_en = _guard614;
assign l7_idx_clk = clk;
assign l7_idx_reset = reset;
assign l7_idx_in =
  _guard617 ? 4'd0 :
  _guard620 ? l7_add_out :
  'x;
assign idx_between_26_27_reg_write_en = _guard625;
assign idx_between_26_27_reg_clk = clk;
assign idx_between_26_27_reg_reset = reset;
assign idx_between_26_27_reg_in =
  _guard626 ? idx_between_26_27_comb_out :
  _guard629 ? 1'd0 :
  'x;
assign index_lt_13_left = idx_add_out;
assign index_lt_13_right = 5'd13;
assign index_ge_14_left = idx_add_out;
assign index_ge_14_right = 5'd14;
assign index_ge_8_left = idx_add_out;
assign index_ge_8_right = 5'd8;
assign index_lt_17_left = idx_add_out;
assign index_lt_17_right = 5'd17;
assign idx_between_25_26_reg_write_en = _guard642;
assign idx_between_25_26_reg_clk = clk;
assign idx_between_25_26_reg_reset = reset;
assign idx_between_25_26_reg_in =
  _guard645 ? 1'd0 :
  _guard646 ? idx_between_25_26_comb_out :
  'x;
assign idx_between_15_16_reg_write_en = _guard651;
assign idx_between_15_16_reg_clk = clk;
assign idx_between_15_16_reg_reset = reset;
assign idx_between_15_16_reg_in =
  _guard652 ? idx_between_15_16_comb_out :
  _guard655 ? 1'd0 :
  'x;
assign idx_between_6_10_reg_write_en = _guard660;
assign idx_between_6_10_reg_clk = clk;
assign idx_between_6_10_reg_reset = reset;
assign idx_between_6_10_reg_in =
  _guard661 ? idx_between_6_10_comb_out :
  _guard664 ? 1'd0 :
  'x;
assign idx_between_20_21_reg_write_en = _guard669;
assign idx_between_20_21_reg_clk = clk;
assign idx_between_20_21_reg_reset = reset;
assign idx_between_20_21_reg_in =
  _guard672 ? 1'd0 :
  _guard673 ? idx_between_20_21_comb_out :
  'x;
assign done = _guard674;
assign t2_addr0 =
  _guard677 ? t2_idx_out :
  4'd0;
assign t3_reset = reset;
assign out_mem_4_write_data =
  _guard680 ? pe_4_0_out :
  _guard683 ? pe_4_5_out :
  _guard686 ? pe_4_6_out :
  _guard689 ? pe_4_2_out :
  _guard692 ? pe_4_4_out :
  _guard695 ? pe_4_7_out :
  _guard698 ? pe_4_3_out :
  _guard701 ? pe_4_1_out :
  32'd0;
assign t0_reset = reset;
assign t6_reset = reset;
assign l5_addr0 =
  _guard704 ? l5_idx_out :
  4'd0;
assign l5_clk = clk;
assign out_mem_2_reset = reset;
assign t2_clk = clk;
assign l0_addr0 =
  _guard707 ? l0_idx_out :
  4'd0;
assign l3_clk = clk;
assign out_mem_1_addr0 =
  _guard710 ? 4'd3 :
  _guard713 ? 4'd5 :
  _guard716 ? 4'd4 :
  _guard719 ? 4'd0 :
  _guard722 ? 4'd7 :
  _guard725 ? 4'd2 :
  _guard728 ? 4'd6 :
  _guard731 ? 4'd1 :
  4'd0;
assign out_mem_1_clk = clk;
assign out_mem_3_reset = reset;
assign out_mem_5_addr0 =
  _guard734 ? 4'd3 :
  _guard737 ? 4'd5 :
  _guard740 ? 4'd4 :
  _guard743 ? 4'd0 :
  _guard746 ? 4'd7 :
  _guard749 ? 4'd2 :
  _guard752 ? 4'd6 :
  _guard755 ? 4'd1 :
  4'd0;
assign out_mem_5_write_data =
  _guard758 ? pe_5_2_out :
  _guard761 ? pe_5_0_out :
  _guard764 ? pe_5_4_out :
  _guard767 ? pe_5_1_out :
  _guard770 ? pe_5_7_out :
  _guard773 ? pe_5_3_out :
  _guard776 ? pe_5_5_out :
  _guard779 ? pe_5_6_out :
  32'd0;
assign l6_addr0 =
  _guard782 ? l6_idx_out :
  4'd0;
assign out_mem_0_write_data =
  _guard785 ? pe_0_1_out :
  _guard788 ? pe_0_7_out :
  _guard791 ? pe_0_3_out :
  _guard794 ? pe_0_5_out :
  _guard797 ? pe_0_2_out :
  _guard800 ? pe_0_4_out :
  _guard803 ? pe_0_0_out :
  _guard806 ? pe_0_6_out :
  32'd0;
assign out_mem_5_clk = clk;
assign t5_reset = reset;
assign l7_reset = reset;
assign out_mem_6_addr0 =
  _guard809 ? 4'd3 :
  _guard812 ? 4'd5 :
  _guard815 ? 4'd4 :
  _guard818 ? 4'd0 :
  _guard821 ? 4'd7 :
  _guard824 ? 4'd2 :
  _guard827 ? 4'd6 :
  _guard830 ? 4'd1 :
  4'd0;
assign t0_clk = clk;
assign l5_reset = reset;
assign out_mem_1_reset = reset;
assign out_mem_3_write_data =
  _guard833 ? pe_3_4_out :
  _guard836 ? pe_3_7_out :
  _guard839 ? pe_3_2_out :
  _guard842 ? pe_3_5_out :
  _guard845 ? pe_3_6_out :
  _guard848 ? pe_3_0_out :
  _guard851 ? pe_3_1_out :
  _guard854 ? pe_3_3_out :
  32'd0;
assign t4_reset = reset;
assign t5_addr0 =
  _guard857 ? t5_idx_out :
  4'd0;
assign t5_clk = clk;
assign t6_clk = clk;
assign l0_reset = reset;
assign l1_addr0 =
  _guard860 ? l1_idx_out :
  4'd0;
assign l7_clk = clk;
assign out_mem_5_write_en = _guard909;
assign out_mem_5_reset = reset;
assign out_mem_7_addr0 =
  _guard912 ? 4'd3 :
  _guard915 ? 4'd5 :
  _guard918 ? 4'd4 :
  _guard921 ? 4'd0 :
  _guard924 ? 4'd7 :
  _guard927 ? 4'd2 :
  _guard930 ? 4'd6 :
  _guard933 ? 4'd1 :
  4'd0;
assign t4_clk = clk;
assign t4_addr0 =
  _guard936 ? t4_idx_out :
  4'd0;
assign t6_addr0 =
  _guard939 ? t6_idx_out :
  4'd0;
assign out_mem_0_clk = clk;
assign out_mem_7_write_en = _guard988;
assign out_mem_7_clk = clk;
assign out_mem_7_reset = reset;
assign t1_reset = reset;
assign l6_clk = clk;
assign out_mem_3_clk = clk;
assign out_mem_4_addr0 =
  _guard991 ? 4'd3 :
  _guard994 ? 4'd5 :
  _guard997 ? 4'd4 :
  _guard1000 ? 4'd0 :
  _guard1003 ? 4'd7 :
  _guard1006 ? 4'd2 :
  _guard1009 ? 4'd6 :
  _guard1012 ? 4'd1 :
  4'd0;
assign out_mem_4_clk = clk;
assign out_mem_4_reset = reset;
assign out_mem_6_reset = reset;
assign t7_clk = clk;
assign l3_addr0 =
  _guard1015 ? l3_idx_out :
  4'd0;
assign l4_reset = reset;
assign out_mem_2_write_data =
  _guard1018 ? pe_2_7_out :
  _guard1021 ? pe_2_4_out :
  _guard1024 ? pe_2_1_out :
  _guard1027 ? pe_2_3_out :
  _guard1030 ? pe_2_5_out :
  _guard1033 ? pe_2_6_out :
  _guard1036 ? pe_2_0_out :
  _guard1039 ? pe_2_2_out :
  32'd0;
assign l4_addr0 =
  _guard1042 ? l4_idx_out :
  4'd0;
assign l7_addr0 =
  _guard1045 ? l7_idx_out :
  4'd0;
assign out_mem_0_reset = reset;
assign out_mem_1_write_data =
  _guard1048 ? pe_1_4_out :
  _guard1051 ? pe_1_7_out :
  _guard1054 ? pe_1_2_out :
  _guard1057 ? pe_1_3_out :
  _guard1060 ? pe_1_0_out :
  _guard1063 ? pe_1_6_out :
  _guard1066 ? pe_1_5_out :
  _guard1069 ? pe_1_1_out :
  32'd0;
assign out_mem_1_write_en = _guard1118;
assign out_mem_4_write_en = _guard1167;
assign out_mem_6_clk = clk;
assign t0_addr0 =
  _guard1170 ? t0_idx_out :
  4'd0;
assign t1_addr0 =
  _guard1173 ? t1_idx_out :
  4'd0;
assign t1_clk = clk;
assign l1_reset = reset;
assign l2_clk = clk;
assign l2_reset = reset;
assign out_mem_0_write_en = _guard1222;
assign out_mem_2_write_en = _guard1271;
assign out_mem_2_clk = clk;
assign t3_clk = clk;
assign t7_reset = reset;
assign out_mem_3_write_en = _guard1320;
assign out_mem_6_write_data =
  _guard1323 ? pe_6_4_out :
  _guard1326 ? pe_6_0_out :
  _guard1329 ? pe_6_1_out :
  _guard1332 ? pe_6_5_out :
  _guard1335 ? pe_6_2_out :
  _guard1338 ? pe_6_3_out :
  _guard1341 ? pe_6_7_out :
  _guard1344 ? pe_6_6_out :
  32'd0;
assign out_mem_6_write_en = _guard1393;
assign out_mem_7_write_data =
  _guard1396 ? pe_7_3_out :
  _guard1399 ? pe_7_4_out :
  _guard1402 ? pe_7_0_out :
  _guard1405 ? pe_7_5_out :
  _guard1408 ? pe_7_6_out :
  _guard1411 ? pe_7_1_out :
  _guard1414 ? pe_7_2_out :
  _guard1417 ? pe_7_7_out :
  32'd0;
assign l0_clk = clk;
assign l1_clk = clk;
assign l2_addr0 =
  _guard1420 ? l2_idx_out :
  4'd0;
assign l3_reset = reset;
assign l4_clk = clk;
assign l6_reset = reset;
assign out_mem_0_addr0 =
  _guard1423 ? 4'd3 :
  _guard1426 ? 4'd5 :
  _guard1429 ? 4'd4 :
  _guard1432 ? 4'd0 :
  _guard1435 ? 4'd7 :
  _guard1438 ? 4'd2 :
  _guard1441 ? 4'd6 :
  _guard1444 ? 4'd1 :
  4'd0;
assign out_mem_3_addr0 =
  _guard1447 ? 4'd3 :
  _guard1450 ? 4'd5 :
  _guard1453 ? 4'd4 :
  _guard1456 ? 4'd0 :
  _guard1459 ? 4'd7 :
  _guard1462 ? 4'd2 :
  _guard1465 ? 4'd6 :
  _guard1468 ? 4'd1 :
  4'd0;
assign t2_reset = reset;
assign t3_addr0 =
  _guard1471 ? t3_idx_out :
  4'd0;
assign t7_addr0 =
  _guard1474 ? t7_idx_out :
  4'd0;
assign out_mem_2_addr0 =
  _guard1477 ? 4'd3 :
  _guard1480 ? 4'd5 :
  _guard1483 ? 4'd4 :
  _guard1486 ? 4'd0 :
  _guard1489 ? 4'd7 :
  _guard1492 ? 4'd2 :
  _guard1495 ? 4'd6 :
  _guard1498 ? 4'd1 :
  4'd0;
assign cond_wire0_in =
  _guard1499 ? idx_between_1_5_reg_out :
  _guard1502 ? cond0_out :
  1'd0;
assign cond_wire4_in =
  _guard1505 ? cond4_out :
  _guard1506 ? idx_between_1_9_reg_out :
  1'd0;
assign cond6_write_en = _guard1507;
assign cond6_clk = clk;
assign cond6_reset = reset;
assign cond6_in =
  _guard1508 ? idx_between_2_10_reg_out :
  1'd0;
assign cond_wire13_in =
  _guard1509 ? idx_between_15_16_reg_out :
  _guard1512 ? cond13_out :
  1'd0;
assign cond_wire16_in =
  _guard1513 ? idx_between_4_12_reg_out :
  _guard1516 ? cond16_out :
  1'd0;
assign cond30_write_en = _guard1517;
assign cond30_clk = clk;
assign cond30_reset = reset;
assign cond30_in =
  _guard1518 ? idx_between_7_11_reg_out :
  1'd0;
assign cond_wire32_in =
  _guard1519 ? idx_between_11_19_reg_out :
  _guard1522 ? cond32_out :
  1'd0;
assign cond_wire40_in =
  _guard1525 ? cond40_out :
  _guard1526 ? idx_between_2_6_reg_out :
  1'd0;
assign cond44_write_en = _guard1527;
assign cond44_clk = clk;
assign cond44_reset = reset;
assign cond44_in =
  _guard1528 ? idx_between_3_7_reg_out :
  1'd0;
assign cond45_write_en = _guard1529;
assign cond45_clk = clk;
assign cond45_reset = reset;
assign cond45_in =
  _guard1530 ? idx_between_3_11_reg_out :
  1'd0;
assign cond_wire73_in =
  _guard1531 ? idx_between_3_7_reg_out :
  _guard1534 ? cond73_out :
  1'd0;
assign cond81_write_en = _guard1535;
assign cond81_clk = clk;
assign cond81_reset = reset;
assign cond81_in =
  _guard1536 ? idx_between_5_9_reg_out :
  1'd0;
assign cond98_write_en = _guard1537;
assign cond98_clk = clk;
assign cond98_reset = reset;
assign cond98_in =
  _guard1538 ? idx_between_9_17_reg_out :
  1'd0;
assign cond100_write_en = _guard1539;
assign cond100_clk = clk;
assign cond100_reset = reset;
assign cond100_in =
  _guard1540 ? idx_between_21_22_reg_out :
  1'd0;
assign cond_wire101_in =
  _guard1543 ? cond101_out :
  _guard1544 ? idx_between_10_14_reg_out :
  1'd0;
assign cond107_write_en = _guard1545;
assign cond107_clk = clk;
assign cond107_reset = reset;
assign cond107_in =
  _guard1546 ? idx_between_4_12_reg_out :
  1'd0;
assign cond_wire107_in =
  _guard1549 ? cond107_out :
  _guard1550 ? idx_between_4_12_reg_out :
  1'd0;
assign cond115_write_en = _guard1551;
assign cond115_clk = clk;
assign cond115_reset = reset;
assign cond115_in =
  _guard1552 ? idx_between_6_14_reg_out :
  1'd0;
assign cond_wire121_in =
  _guard1555 ? cond121_out :
  _guard1556 ? idx_between_19_20_reg_out :
  1'd0;
assign cond_wire127_in =
  _guard1559 ? cond127_out :
  _guard1560 ? idx_between_9_17_reg_out :
  1'd0;
assign cond_wire144_in =
  _guard1561 ? idx_between_6_14_reg_out :
  _guard1564 ? cond144_out :
  1'd0;
assign cond149_write_en = _guard1565;
assign cond149_clk = clk;
assign cond149_reset = reset;
assign cond149_in =
  _guard1566 ? idx_between_11_19_reg_out :
  1'd0;
assign cond150_write_en = _guard1567;
assign cond150_clk = clk;
assign cond150_reset = reset;
assign cond150_in =
  _guard1568 ? idx_between_19_20_reg_out :
  1'd0;
assign cond_wire160_in =
  _guard1569 ? idx_between_10_18_reg_out :
  _guard1572 ? cond160_out :
  1'd0;
assign cond169_write_en = _guard1573;
assign cond169_clk = clk;
assign cond169_reset = reset;
assign cond169_in =
  _guard1574 ? idx_between_16_24_reg_out :
  1'd0;
assign cond179_write_en = _guard1575;
assign cond179_clk = clk;
assign cond179_reset = reset;
assign cond179_in =
  _guard1576 ? idx_between_19_20_reg_out :
  1'd0;
assign cond193_write_en = _guard1577;
assign cond193_clk = clk;
assign cond193_reset = reset;
assign cond193_in =
  _guard1578 ? idx_between_11_19_reg_out :
  1'd0;
assign cond_wire208_in =
  _guard1579 ? idx_between_19_20_reg_out :
  _guard1582 ? cond208_out :
  1'd0;
assign cond214_write_en = _guard1583;
assign cond214_clk = clk;
assign cond214_reset = reset;
assign cond214_in =
  _guard1584 ? idx_between_9_17_reg_out :
  1'd0;
assign cond_wire230_in =
  _guard1587 ? cond230_out :
  _guard1588 ? idx_between_13_21_reg_out :
  1'd0;
assign cond236_write_en = _guard1589;
assign cond236_clk = clk;
assign cond236_reset = reset;
assign cond236_in =
  _guard1590 ? idx_between_26_27_reg_out :
  1'd0;
assign cond_wire239_in =
  _guard1593 ? cond239_out :
  _guard1594 ? idx_between_8_16_reg_out :
  1'd0;
assign cond245_write_en = _guard1595;
assign cond245_clk = clk;
assign cond245_reset = reset;
assign cond245_in =
  _guard1596 ? idx_between_21_22_reg_out :
  1'd0;
assign cond255_write_en = _guard1597;
assign cond255_clk = clk;
assign cond255_reset = reset;
assign cond255_in =
  _guard1598 ? idx_between_12_20_reg_out :
  1'd0;
assign cond_wire261_in =
  _guard1599 ? idx_between_25_26_reg_out :
  _guard1602 ? cond261_out :
  1'd0;
assign fsm_write_en = _guard1603;
assign fsm_clk = clk;
assign fsm_reset = reset;
assign fsm_in =
  _guard1606 ? 1'd0 :
  _guard1609 ? adder0_out :
  1'd0;
assign adder_left =
  _guard1610 ? fsm0_out :
  5'd0;
assign adder_right =
  _guard1611 ? 5'd1 :
  5'd0;
assign early_reset_static_par0_go_in = _guard1616;
assign top_0_6_write_en = _guard1619;
assign top_0_6_clk = clk;
assign top_0_6_reset = reset;
assign top_0_6_in = t6_read_data;
assign left_1_4_write_en = _guard1625;
assign left_1_4_clk = clk;
assign left_1_4_reset = reset;
assign left_1_4_in = left_1_3_out;
assign top_1_5_write_en = _guard1631;
assign top_1_5_clk = clk;
assign top_1_5_reset = reset;
assign top_1_5_in = top_0_5_out;
assign left_1_5_write_en = _guard1637;
assign left_1_5_clk = clk;
assign left_1_5_reset = reset;
assign left_1_5_in = left_1_4_out;
assign pe_3_4_mul_ready =
  _guard1643 ? 1'd1 :
  _guard1646 ? 1'd0 :
  1'd0;
assign pe_3_4_clk = clk;
assign pe_3_4_top =
  _guard1659 ? top_3_4_out :
  32'd0;
assign pe_3_4_left =
  _guard1672 ? left_3_4_out :
  32'd0;
assign pe_3_4_reset = reset;
assign pe_3_4_go = _guard1685;
assign pe_3_7_mul_ready =
  _guard1688 ? 1'd1 :
  _guard1691 ? 1'd0 :
  1'd0;
assign pe_3_7_clk = clk;
assign pe_3_7_top =
  _guard1704 ? top_3_7_out :
  32'd0;
assign pe_3_7_left =
  _guard1717 ? left_3_7_out :
  32'd0;
assign pe_3_7_reset = reset;
assign pe_3_7_go = _guard1730;
assign pe_4_0_mul_ready =
  _guard1733 ? 1'd1 :
  _guard1736 ? 1'd0 :
  1'd0;
assign pe_4_0_clk = clk;
assign pe_4_0_top =
  _guard1749 ? top_4_0_out :
  32'd0;
assign pe_4_0_left =
  _guard1762 ? left_4_0_out :
  32'd0;
assign pe_4_0_reset = reset;
assign pe_4_0_go = _guard1775;
assign left_4_2_write_en = _guard1778;
assign left_4_2_clk = clk;
assign left_4_2_reset = reset;
assign left_4_2_in = left_4_1_out;
assign pe_5_0_mul_ready =
  _guard1784 ? 1'd1 :
  _guard1787 ? 1'd0 :
  1'd0;
assign pe_5_0_clk = clk;
assign pe_5_0_top =
  _guard1800 ? top_5_0_out :
  32'd0;
assign pe_5_0_left =
  _guard1813 ? left_5_0_out :
  32'd0;
assign pe_5_0_reset = reset;
assign pe_5_0_go = _guard1826;
assign left_5_6_write_en = _guard1829;
assign left_5_6_clk = clk;
assign left_5_6_reset = reset;
assign left_5_6_in = left_5_5_out;
assign left_6_5_write_en = _guard1835;
assign left_6_5_clk = clk;
assign left_6_5_reset = reset;
assign left_6_5_in = left_6_4_out;
assign top_6_6_write_en = _guard1841;
assign top_6_6_clk = clk;
assign top_6_6_reset = reset;
assign top_6_6_in = top_5_6_out;
assign l0_idx_write_en = _guard1851;
assign l0_idx_clk = clk;
assign l0_idx_reset = reset;
assign l0_idx_in =
  _guard1854 ? 4'd0 :
  _guard1857 ? l0_add_out :
  'x;
assign idx_between_5_13_reg_write_en = _guard1862;
assign idx_between_5_13_reg_clk = clk;
assign idx_between_5_13_reg_reset = reset;
assign idx_between_5_13_reg_in =
  _guard1865 ? 1'd0 :
  _guard1866 ? idx_between_5_13_comb_out :
  'x;
assign idx_between_9_17_comb_left = index_ge_9_out;
assign idx_between_9_17_comb_right = index_lt_17_out;
assign idx_between_17_18_reg_write_en = _guard1873;
assign idx_between_17_18_reg_clk = clk;
assign idx_between_17_18_reg_reset = reset;
assign idx_between_17_18_reg_in =
  _guard1874 ? idx_between_17_18_comb_out :
  _guard1877 ? 1'd0 :
  'x;
assign idx_between_17_18_comb_left = index_ge_17_out;
assign idx_between_17_18_comb_right = index_lt_18_out;
assign idx_between_13_14_reg_write_en = _guard1884;
assign idx_between_13_14_reg_clk = clk;
assign idx_between_13_14_reg_reset = reset;
assign idx_between_13_14_reg_in =
  _guard1885 ? idx_between_13_14_comb_out :
  _guard1888 ? 1'd0 :
  'x;
assign idx_between_15_23_comb_left = index_ge_15_out;
assign idx_between_15_23_comb_right = index_lt_23_out;
assign idx_between_23_24_reg_write_en = _guard1895;
assign idx_between_23_24_reg_clk = clk;
assign idx_between_23_24_reg_reset = reset;
assign idx_between_23_24_reg_in =
  _guard1896 ? idx_between_23_24_comb_out :
  _guard1899 ? 1'd0 :
  'x;
assign idx_between_15_16_comb_left = index_ge_15_out;
assign idx_between_15_16_comb_right = index_lt_16_out;
assign index_ge_24_left = idx_add_out;
assign index_ge_24_right = 5'd24;
assign index_lt_11_left = idx_add_out;
assign index_lt_11_right = 5'd11;
assign idx_between_7_11_reg_write_en = _guard1910;
assign idx_between_7_11_reg_clk = clk;
assign idx_between_7_11_reg_reset = reset;
assign idx_between_7_11_reg_in =
  _guard1913 ? 1'd0 :
  _guard1914 ? idx_between_7_11_comb_out :
  'x;
assign cond11_write_en = _guard1915;
assign cond11_clk = clk;
assign cond11_reset = reset;
assign cond11_in =
  _guard1916 ? idx_between_3_11_reg_out :
  1'd0;
assign cond15_write_en = _guard1917;
assign cond15_clk = clk;
assign cond15_reset = reset;
assign cond15_in =
  _guard1918 ? idx_between_4_8_reg_out :
  1'd0;
assign cond_wire27_in =
  _guard1919 ? idx_between_10_18_reg_out :
  _guard1922 ? cond27_out :
  1'd0;
assign cond43_write_en = _guard1923;
assign cond43_clk = clk;
assign cond43_reset = reset;
assign cond43_in =
  _guard1924 ? idx_between_14_15_reg_out :
  1'd0;
assign cond_wire43_in =
  _guard1927 ? cond43_out :
  _guard1928 ? idx_between_14_15_reg_out :
  1'd0;
assign cond_wire44_in =
  _guard1929 ? idx_between_3_7_reg_out :
  _guard1932 ? cond44_out :
  1'd0;
assign cond62_write_en = _guard1933;
assign cond62_clk = clk;
assign cond62_reset = reset;
assign cond62_in =
  _guard1934 ? idx_between_11_19_reg_out :
  1'd0;
assign cond_wire63_in =
  _guard1935 ? idx_between_19_20_reg_out :
  _guard1938 ? cond63_out :
  1'd0;
assign cond_wire67_in =
  _guard1939 ? idx_between_20_21_reg_out :
  _guard1942 ? cond67_out :
  1'd0;
assign cond73_write_en = _guard1943;
assign cond73_clk = clk;
assign cond73_reset = reset;
assign cond73_in =
  _guard1944 ? idx_between_3_7_reg_out :
  1'd0;
assign cond_wire77_in =
  _guard1945 ? idx_between_4_8_reg_out :
  _guard1948 ? cond77_out :
  1'd0;
assign cond103_write_en = _guard1949;
assign cond103_clk = clk;
assign cond103_reset = reset;
assign cond103_in =
  _guard1950 ? idx_between_14_22_reg_out :
  1'd0;
assign cond114_write_en = _guard1951;
assign cond114_clk = clk;
assign cond114_reset = reset;
assign cond114_in =
  _guard1952 ? idx_between_6_10_reg_out :
  1'd0;
assign cond118_write_en = _guard1953;
assign cond118_clk = clk;
assign cond118_reset = reset;
assign cond118_in =
  _guard1954 ? idx_between_7_11_reg_out :
  1'd0;
assign cond121_write_en = _guard1955;
assign cond121_clk = clk;
assign cond121_reset = reset;
assign cond121_in =
  _guard1956 ? idx_between_19_20_reg_out :
  1'd0;
assign cond123_write_en = _guard1957;
assign cond123_clk = clk;
assign cond123_reset = reset;
assign cond123_in =
  _guard1958 ? idx_between_8_16_reg_out :
  1'd0;
assign cond_wire126_in =
  _guard1959 ? idx_between_9_13_reg_out :
  _guard1962 ? cond126_out :
  1'd0;
assign cond_wire154_in =
  _guard1963 ? idx_between_20_21_reg_out :
  _guard1966 ? cond154_out :
  1'd0;
assign cond_wire195_in =
  _guard1967 ? idx_between_23_24_reg_out :
  _guard1970 ? cond195_out :
  1'd0;
assign cond206_write_en = _guard1971;
assign cond206_clk = clk;
assign cond206_reset = reset;
assign cond206_in =
  _guard1972 ? idx_between_7_15_reg_out :
  1'd0;
assign cond216_write_en = _guard1973;
assign cond216_clk = clk;
assign cond216_reset = reset;
assign cond216_in =
  _guard1974 ? idx_between_21_22_reg_out :
  1'd0;
assign cond_wire218_in =
  _guard1975 ? idx_between_10_18_reg_out :
  _guard1978 ? cond218_out :
  1'd0;
assign cond_wire238_in =
  _guard1979 ? idx_between_8_12_reg_out :
  _guard1982 ? cond238_out :
  1'd0;
assign cond240_write_en = _guard1983;
assign cond240_clk = clk;
assign cond240_reset = reset;
assign cond240_in =
  _guard1984 ? idx_between_12_20_reg_out :
  1'd0;
assign cond251_write_en = _guard1985;
assign cond251_clk = clk;
assign cond251_reset = reset;
assign cond251_in =
  _guard1986 ? idx_between_11_19_reg_out :
  1'd0;
assign cond264_write_en = _guard1987;
assign cond264_clk = clk;
assign cond264_reset = reset;
assign cond264_in =
  _guard1988 ? idx_between_18_26_reg_out :
  1'd0;
assign cond_wire265_in =
  _guard1989 ? idx_between_26_27_reg_out :
  _guard1992 ? cond265_out :
  1'd0;
assign pe_0_1_mul_ready =
  _guard1995 ? 1'd1 :
  _guard1998 ? 1'd0 :
  1'd0;
assign pe_0_1_clk = clk;
assign pe_0_1_top =
  _guard2011 ? top_0_1_out :
  32'd0;
assign pe_0_1_left =
  _guard2024 ? left_0_1_out :
  32'd0;
assign pe_0_1_reset = reset;
assign pe_0_1_go = _guard2037;
assign left_0_6_write_en = _guard2040;
assign left_0_6_clk = clk;
assign left_0_6_reset = reset;
assign left_0_6_in = left_0_5_out;
assign pe_0_7_mul_ready =
  _guard2046 ? 1'd1 :
  _guard2049 ? 1'd0 :
  1'd0;
assign pe_0_7_clk = clk;
assign pe_0_7_top =
  _guard2062 ? top_0_7_out :
  32'd0;
assign pe_0_7_left =
  _guard2075 ? left_0_7_out :
  32'd0;
assign pe_0_7_reset = reset;
assign pe_0_7_go = _guard2088;
assign left_1_2_write_en = _guard2091;
assign left_1_2_clk = clk;
assign left_1_2_reset = reset;
assign left_1_2_in = left_1_1_out;
assign left_2_2_write_en = _guard2097;
assign left_2_2_clk = clk;
assign left_2_2_reset = reset;
assign left_2_2_in = left_2_1_out;
assign top_2_5_write_en = _guard2103;
assign top_2_5_clk = clk;
assign top_2_5_reset = reset;
assign top_2_5_in = top_1_5_out;
assign pe_2_7_mul_ready =
  _guard2109 ? 1'd1 :
  _guard2112 ? 1'd0 :
  1'd0;
assign pe_2_7_clk = clk;
assign pe_2_7_top =
  _guard2125 ? top_2_7_out :
  32'd0;
assign pe_2_7_left =
  _guard2138 ? left_2_7_out :
  32'd0;
assign pe_2_7_reset = reset;
assign pe_2_7_go = _guard2151;
assign left_2_7_write_en = _guard2154;
assign left_2_7_clk = clk;
assign left_2_7_reset = reset;
assign left_2_7_in = left_2_6_out;
assign pe_4_5_mul_ready =
  _guard2160 ? 1'd1 :
  _guard2163 ? 1'd0 :
  1'd0;
assign pe_4_5_clk = clk;
assign pe_4_5_top =
  _guard2176 ? top_4_5_out :
  32'd0;
assign pe_4_5_left =
  _guard2189 ? left_4_5_out :
  32'd0;
assign pe_4_5_reset = reset;
assign pe_4_5_go = _guard2202;
assign left_4_5_write_en = _guard2205;
assign left_4_5_clk = clk;
assign left_4_5_reset = reset;
assign left_4_5_in = left_4_4_out;
assign top_5_0_write_en = _guard2211;
assign top_5_0_clk = clk;
assign top_5_0_reset = reset;
assign top_5_0_in = top_4_0_out;
assign top_5_3_write_en = _guard2217;
assign top_5_3_clk = clk;
assign top_5_3_reset = reset;
assign top_5_3_in = top_4_3_out;
assign l3_add_left = 4'd1;
assign l3_add_right = l3_idx_out;
assign index_ge_3_left = idx_add_out;
assign index_ge_3_right = 5'd3;
assign index_ge_12_left = idx_add_out;
assign index_ge_12_right = 5'd12;
assign idx_between_6_14_reg_write_en = _guard2235;
assign idx_between_6_14_reg_clk = clk;
assign idx_between_6_14_reg_reset = reset;
assign idx_between_6_14_reg_in =
  _guard2238 ? 1'd0 :
  _guard2239 ? idx_between_6_14_comb_out :
  'x;
assign index_lt_19_left = idx_add_out;
assign index_lt_19_right = 5'd19;
assign idx_between_4_8_reg_write_en = _guard2246;
assign idx_between_4_8_reg_clk = clk;
assign idx_between_4_8_reg_reset = reset;
assign idx_between_4_8_reg_in =
  _guard2249 ? 1'd0 :
  _guard2250 ? idx_between_4_8_comb_out :
  'x;
assign idx_between_5_9_comb_left = index_ge_5_out;
assign idx_between_5_9_comb_right = index_lt_9_out;
assign idx_between_9_13_comb_left = index_ge_9_out;
assign idx_between_9_13_comb_right = index_lt_13_out;
assign idx_between_10_14_comb_left = index_ge_10_out;
assign idx_between_10_14_comb_right = index_lt_14_out;
assign idx_between_2_10_comb_left = index_ge_2_out;
assign idx_between_2_10_comb_right = index_lt_10_out;
assign idx_between_6_10_comb_left = index_ge_6_out;
assign idx_between_6_10_comb_right = index_lt_10_out;
assign idx_between_16_24_comb_left = index_ge_16_out;
assign idx_between_16_24_comb_right = index_lt_24_out;
assign cond_write_en = _guard2263;
assign cond_clk = clk;
assign cond_reset = reset;
assign cond_in =
  _guard2264 ? idx_between_0_8_reg_out :
  1'd0;
assign cond_wire26_in =
  _guard2265 ? idx_between_6_14_reg_out :
  _guard2268 ? cond26_out :
  1'd0;
assign cond35_write_en = _guard2269;
assign cond35_clk = clk;
assign cond35_reset = reset;
assign cond35_in =
  _guard2270 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire35_in =
  _guard2273 ? cond35_out :
  _guard2274 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire50_in =
  _guard2277 ? cond50_out :
  _guard2278 ? idx_between_8_16_reg_out :
  1'd0;
assign cond_wire56_in =
  _guard2279 ? idx_between_6_10_reg_out :
  _guard2282 ? cond56_out :
  1'd0;
assign cond60_write_en = _guard2283;
assign cond60_clk = clk;
assign cond60_reset = reset;
assign cond60_in =
  _guard2284 ? idx_between_7_11_reg_out :
  1'd0;
assign cond69_write_en = _guard2285;
assign cond69_clk = clk;
assign cond69_reset = reset;
assign cond69_in =
  _guard2286 ? idx_between_9_17_reg_out :
  1'd0;
assign cond72_write_en = _guard2287;
assign cond72_clk = clk;
assign cond72_reset = reset;
assign cond72_in =
  _guard2288 ? idx_between_2_10_reg_out :
  1'd0;
assign cond76_write_en = _guard2289;
assign cond76_clk = clk;
assign cond76_reset = reset;
assign cond76_in =
  _guard2290 ? idx_between_15_16_reg_out :
  1'd0;
assign cond_wire85_in =
  _guard2291 ? idx_between_6_10_reg_out :
  _guard2294 ? cond85_out :
  1'd0;
assign cond92_write_en = _guard2295;
assign cond92_clk = clk;
assign cond92_reset = reset;
assign cond92_in =
  _guard2296 ? idx_between_19_20_reg_out :
  1'd0;
assign cond_wire116_in =
  _guard2297 ? idx_between_10_18_reg_out :
  _guard2300 ? cond116_out :
  1'd0;
assign cond_wire149_in =
  _guard2301 ? idx_between_11_19_reg_out :
  _guard2304 ? cond149_out :
  1'd0;
assign cond_wire163_in =
  _guard2307 ? cond163_out :
  _guard2308 ? idx_between_11_15_reg_out :
  1'd0;
assign cond_wire182_in =
  _guard2309 ? idx_between_12_20_reg_out :
  _guard2312 ? cond182_out :
  1'd0;
assign cond189_write_en = _guard2313;
assign cond189_clk = clk;
assign cond189_reset = reset;
assign cond189_in =
  _guard2314 ? idx_between_10_18_reg_out :
  1'd0;
assign cond_wire192_in =
  _guard2317 ? cond192_out :
  _guard2318 ? idx_between_11_15_reg_out :
  1'd0;
assign cond_wire200_in =
  _guard2319 ? idx_between_13_17_reg_out :
  _guard2322 ? cond200_out :
  1'd0;
assign cond_wire205_in =
  _guard2323 ? idx_between_7_11_reg_out :
  _guard2326 ? cond205_out :
  1'd0;
assign cond226_write_en = _guard2327;
assign cond226_clk = clk;
assign cond226_reset = reset;
assign cond226_in =
  _guard2328 ? idx_between_12_20_reg_out :
  1'd0;
assign cond233_write_en = _guard2329;
assign cond233_clk = clk;
assign cond233_reset = reset;
assign cond233_in =
  _guard2330 ? idx_between_14_18_reg_out :
  1'd0;
assign cond241_write_en = _guard2331;
assign cond241_clk = clk;
assign cond241_reset = reset;
assign cond241_in =
  _guard2332 ? idx_between_20_21_reg_out :
  1'd0;
assign cond_wire243_in =
  _guard2335 ? cond243_out :
  _guard2336 ? idx_between_9_17_reg_out :
  1'd0;
assign cond_wire245_in =
  _guard2339 ? cond245_out :
  _guard2340 ? idx_between_21_22_reg_out :
  1'd0;
assign cond248_write_en = _guard2341;
assign cond248_clk = clk;
assign cond248_reset = reset;
assign cond248_in =
  _guard2342 ? idx_between_14_22_reg_out :
  1'd0;
assign cond257_write_en = _guard2343;
assign cond257_clk = clk;
assign cond257_reset = reset;
assign cond257_in =
  _guard2344 ? idx_between_24_25_reg_out :
  1'd0;
assign cond_wire263_in =
  _guard2347 ? cond263_out :
  _guard2348 ? idx_between_14_22_reg_out :
  1'd0;
assign cond266_write_en = _guard2349;
assign cond266_clk = clk;
assign cond266_reset = reset;
assign cond266_in =
  _guard2350 ? idx_between_15_19_reg_out :
  1'd0;
assign pe_1_0_mul_ready =
  _guard2353 ? 1'd1 :
  _guard2356 ? 1'd0 :
  1'd0;
assign pe_1_0_clk = clk;
assign pe_1_0_top =
  _guard2369 ? top_1_0_out :
  32'd0;
assign pe_1_0_left =
  _guard2382 ? left_1_0_out :
  32'd0;
assign pe_1_0_reset = reset;
assign pe_1_0_go = _guard2395;
assign left_1_0_write_en = _guard2398;
assign left_1_0_clk = clk;
assign left_1_0_reset = reset;
assign left_1_0_in = l1_read_data;
assign left_1_1_write_en = _guard2404;
assign left_1_1_clk = clk;
assign left_1_1_reset = reset;
assign left_1_1_in = left_1_0_out;
assign top_1_2_write_en = _guard2410;
assign top_1_2_clk = clk;
assign top_1_2_reset = reset;
assign top_1_2_in = top_0_2_out;
assign left_2_0_write_en = _guard2416;
assign left_2_0_clk = clk;
assign left_2_0_reset = reset;
assign left_2_0_in = l2_read_data;
assign left_3_1_write_en = _guard2422;
assign left_3_1_clk = clk;
assign left_3_1_reset = reset;
assign left_3_1_in = left_3_0_out;
assign pe_3_2_mul_ready =
  _guard2428 ? 1'd1 :
  _guard2431 ? 1'd0 :
  1'd0;
assign pe_3_2_clk = clk;
assign pe_3_2_top =
  _guard2444 ? top_3_2_out :
  32'd0;
assign pe_3_2_left =
  _guard2457 ? left_3_2_out :
  32'd0;
assign pe_3_2_reset = reset;
assign pe_3_2_go = _guard2470;
assign pe_3_5_mul_ready =
  _guard2473 ? 1'd1 :
  _guard2476 ? 1'd0 :
  1'd0;
assign pe_3_5_clk = clk;
assign pe_3_5_top =
  _guard2489 ? top_3_5_out :
  32'd0;
assign pe_3_5_left =
  _guard2502 ? left_3_5_out :
  32'd0;
assign pe_3_5_reset = reset;
assign pe_3_5_go = _guard2515;
assign pe_3_6_mul_ready =
  _guard2518 ? 1'd1 :
  _guard2521 ? 1'd0 :
  1'd0;
assign pe_3_6_clk = clk;
assign pe_3_6_top =
  _guard2534 ? top_3_6_out :
  32'd0;
assign pe_3_6_left =
  _guard2547 ? left_3_6_out :
  32'd0;
assign pe_3_6_reset = reset;
assign pe_3_6_go = _guard2560;
assign left_3_7_write_en = _guard2563;
assign left_3_7_clk = clk;
assign left_3_7_reset = reset;
assign left_3_7_in = left_3_6_out;
assign top_4_5_write_en = _guard2569;
assign top_4_5_clk = clk;
assign top_4_5_reset = reset;
assign top_4_5_in = top_3_5_out;
assign pe_5_4_mul_ready =
  _guard2575 ? 1'd1 :
  _guard2578 ? 1'd0 :
  1'd0;
assign pe_5_4_clk = clk;
assign pe_5_4_top =
  _guard2591 ? top_5_4_out :
  32'd0;
assign pe_5_4_left =
  _guard2604 ? left_5_4_out :
  32'd0;
assign pe_5_4_reset = reset;
assign pe_5_4_go = _guard2617;
assign top_7_2_write_en = _guard2620;
assign top_7_2_clk = clk;
assign top_7_2_reset = reset;
assign top_7_2_in = top_6_2_out;
assign pe_7_4_mul_ready =
  _guard2626 ? 1'd1 :
  _guard2629 ? 1'd0 :
  1'd0;
assign pe_7_4_clk = clk;
assign pe_7_4_top =
  _guard2642 ? top_7_4_out :
  32'd0;
assign pe_7_4_left =
  _guard2655 ? left_7_4_out :
  32'd0;
assign pe_7_4_reset = reset;
assign pe_7_4_go = _guard2668;
assign t1_idx_write_en = _guard2675;
assign t1_idx_clk = clk;
assign t1_idx_reset = reset;
assign t1_idx_in =
  _guard2678 ? 4'd0 :
  _guard2681 ? t1_add_out :
  'x;
assign t7_idx_write_en = _guard2688;
assign t7_idx_clk = clk;
assign t7_idx_reset = reset;
assign t7_idx_in =
  _guard2691 ? 4'd0 :
  _guard2694 ? t7_add_out :
  'x;
assign index_ge_18_left = idx_add_out;
assign index_ge_18_right = 5'd18;
assign idx_between_26_27_comb_left = index_ge_26_out;
assign idx_between_26_27_comb_right = index_lt_27_out;
assign idx_between_19_27_reg_write_en = _guard2703;
assign idx_between_19_27_reg_clk = clk;
assign idx_between_19_27_reg_reset = reset;
assign idx_between_19_27_reg_in =
  _guard2706 ? 1'd0 :
  _guard2707 ? idx_between_19_27_comb_out :
  'x;
assign idx_between_15_23_reg_write_en = _guard2712;
assign idx_between_15_23_reg_clk = clk;
assign idx_between_15_23_reg_reset = reset;
assign idx_between_15_23_reg_in =
  _guard2713 ? idx_between_15_23_comb_out :
  _guard2716 ? 1'd0 :
  'x;
assign idx_between_23_24_comb_left = index_ge_23_out;
assign idx_between_23_24_comb_right = index_lt_24_out;
assign idx_between_13_21_comb_left = index_ge_13_out;
assign idx_between_13_21_comb_right = index_lt_21_out;
assign cond18_write_en = _guard2721;
assign cond18_clk = clk;
assign cond18_reset = reset;
assign cond18_in =
  _guard2722 ? idx_between_16_17_reg_out :
  1'd0;
assign cond_wire24_in =
  _guard2723 ? idx_between_5_13_reg_out :
  _guard2726 ? cond24_out :
  1'd0;
assign cond_wire31_in =
  _guard2727 ? idx_between_7_15_reg_out :
  _guard2730 ? cond31_out :
  1'd0;
assign cond_wire46_in =
  _guard2731 ? idx_between_7_15_reg_out :
  _guard2734 ? cond46_out :
  1'd0;
assign cond_wire48_in =
  _guard2735 ? idx_between_4_8_reg_out :
  _guard2738 ? cond48_out :
  1'd0;
assign cond_wire72_in =
  _guard2741 ? cond72_out :
  _guard2742 ? idx_between_2_10_reg_out :
  1'd0;
assign cond_wire76_in =
  _guard2743 ? idx_between_15_16_reg_out :
  _guard2746 ? cond76_out :
  1'd0;
assign cond_wire100_in =
  _guard2749 ? cond100_out :
  _guard2750 ? idx_between_21_22_reg_out :
  1'd0;
assign cond105_write_en = _guard2751;
assign cond105_clk = clk;
assign cond105_reset = reset;
assign cond105_in =
  _guard2752 ? idx_between_3_11_reg_out :
  1'd0;
assign cond_wire134_in =
  _guard2755 ? cond134_out :
  _guard2756 ? idx_between_11_15_reg_out :
  1'd0;
assign cond146_write_en = _guard2757;
assign cond146_clk = clk;
assign cond146_reset = reset;
assign cond146_in =
  _guard2758 ? idx_between_18_19_reg_out :
  1'd0;
assign cond_wire146_in =
  _guard2761 ? cond146_out :
  _guard2762 ? idx_between_18_19_reg_out :
  1'd0;
assign cond151_write_en = _guard2763;
assign cond151_clk = clk;
assign cond151_reset = reset;
assign cond151_in =
  _guard2764 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire157_in =
  _guard2765 ? idx_between_13_21_reg_out :
  _guard2768 ? cond157_out :
  1'd0;
assign cond_wire167_in =
  _guard2771 ? cond167_out :
  _guard2772 ? idx_between_12_16_reg_out :
  1'd0;
assign cond_wire174_in =
  _guard2773 ? idx_between_10_18_reg_out :
  _guard2776 ? cond174_out :
  1'd0;
assign cond177_write_en = _guard2777;
assign cond177_clk = clk;
assign cond177_reset = reset;
assign cond177_in =
  _guard2778 ? idx_between_7_15_reg_out :
  1'd0;
assign cond178_write_en = _guard2779;
assign cond178_clk = clk;
assign cond178_reset = reset;
assign cond178_in =
  _guard2780 ? idx_between_11_19_reg_out :
  1'd0;
assign cond_wire191_in =
  _guard2781 ? idx_between_22_23_reg_out :
  _guard2784 ? cond191_out :
  1'd0;
assign cond_wire198_in =
  _guard2787 ? cond198_out :
  _guard2788 ? idx_between_16_24_reg_out :
  1'd0;
assign cond204_write_en = _guard2789;
assign cond204_clk = clk;
assign cond204_reset = reset;
assign cond204_in =
  _guard2790 ? idx_between_6_14_reg_out :
  1'd0;
assign cond215_write_en = _guard2791;
assign cond215_clk = clk;
assign cond215_reset = reset;
assign cond215_in =
  _guard2792 ? idx_between_13_21_reg_out :
  1'd0;
assign cond_wire216_in =
  _guard2795 ? cond216_out :
  _guard2796 ? idx_between_21_22_reg_out :
  1'd0;
assign cond_wire228_in =
  _guard2799 ? cond228_out :
  _guard2800 ? idx_between_24_25_reg_out :
  1'd0;
assign cond231_write_en = _guard2801;
assign cond231_clk = clk;
assign cond231_reset = reset;
assign cond231_in =
  _guard2802 ? idx_between_17_25_reg_out :
  1'd0;
assign cond_wire231_in =
  _guard2805 ? cond231_out :
  _guard2806 ? idx_between_17_25_reg_out :
  1'd0;
assign cond237_write_en = _guard2807;
assign cond237_clk = clk;
assign cond237_reset = reset;
assign cond237_in =
  _guard2808 ? idx_between_7_15_reg_out :
  1'd0;
assign left_0_0_write_en = _guard2811;
assign left_0_0_clk = clk;
assign left_0_0_reset = reset;
assign left_0_0_in = l0_read_data;
assign pe_0_3_mul_ready =
  _guard2817 ? 1'd1 :
  _guard2820 ? 1'd0 :
  1'd0;
assign pe_0_3_clk = clk;
assign pe_0_3_top =
  _guard2833 ? top_0_3_out :
  32'd0;
assign pe_0_3_left =
  _guard2846 ? left_0_3_out :
  32'd0;
assign pe_0_3_reset = reset;
assign pe_0_3_go = _guard2859;
assign pe_0_5_mul_ready =
  _guard2862 ? 1'd1 :
  _guard2865 ? 1'd0 :
  1'd0;
assign pe_0_5_clk = clk;
assign pe_0_5_top =
  _guard2878 ? top_0_5_out :
  32'd0;
assign pe_0_5_left =
  _guard2891 ? left_0_5_out :
  32'd0;
assign pe_0_5_reset = reset;
assign pe_0_5_go = _guard2904;
assign top_1_3_write_en = _guard2907;
assign top_1_3_clk = clk;
assign top_1_3_reset = reset;
assign top_1_3_in = top_0_3_out;
assign top_1_4_write_en = _guard2913;
assign top_1_4_clk = clk;
assign top_1_4_reset = reset;
assign top_1_4_in = top_0_4_out;
assign left_2_3_write_en = _guard2919;
assign left_2_3_clk = clk;
assign left_2_3_reset = reset;
assign left_2_3_in = left_2_2_out;
assign pe_2_4_mul_ready =
  _guard2925 ? 1'd1 :
  _guard2928 ? 1'd0 :
  1'd0;
assign pe_2_4_clk = clk;
assign pe_2_4_top =
  _guard2941 ? top_2_4_out :
  32'd0;
assign pe_2_4_left =
  _guard2954 ? left_2_4_out :
  32'd0;
assign pe_2_4_reset = reset;
assign pe_2_4_go = _guard2967;
assign top_2_6_write_en = _guard2970;
assign top_2_6_clk = clk;
assign top_2_6_reset = reset;
assign top_2_6_in = top_1_6_out;
assign pe_3_0_mul_ready =
  _guard2976 ? 1'd1 :
  _guard2979 ? 1'd0 :
  1'd0;
assign pe_3_0_clk = clk;
assign pe_3_0_top =
  _guard2992 ? top_3_0_out :
  32'd0;
assign pe_3_0_left =
  _guard3005 ? left_3_0_out :
  32'd0;
assign pe_3_0_reset = reset;
assign pe_3_0_go = _guard3018;
assign top_3_2_write_en = _guard3021;
assign top_3_2_clk = clk;
assign top_3_2_reset = reset;
assign top_3_2_in = top_2_2_out;
assign top_4_0_write_en = _guard3027;
assign top_4_0_clk = clk;
assign top_4_0_reset = reset;
assign top_4_0_in = top_3_0_out;
assign left_4_6_write_en = _guard3033;
assign left_4_6_clk = clk;
assign left_4_6_reset = reset;
assign left_4_6_in = left_4_5_out;
assign left_4_7_write_en = _guard3039;
assign left_4_7_clk = clk;
assign left_4_7_reset = reset;
assign left_4_7_in = left_4_6_out;
assign pe_5_1_mul_ready =
  _guard3045 ? 1'd1 :
  _guard3048 ? 1'd0 :
  1'd0;
assign pe_5_1_clk = clk;
assign pe_5_1_top =
  _guard3061 ? top_5_1_out :
  32'd0;
assign pe_5_1_left =
  _guard3074 ? left_5_1_out :
  32'd0;
assign pe_5_1_reset = reset;
assign pe_5_1_go = _guard3087;
assign pe_5_7_mul_ready =
  _guard3090 ? 1'd1 :
  _guard3093 ? 1'd0 :
  1'd0;
assign pe_5_7_clk = clk;
assign pe_5_7_top =
  _guard3106 ? top_5_7_out :
  32'd0;
assign pe_5_7_left =
  _guard3119 ? left_5_7_out :
  32'd0;
assign pe_5_7_reset = reset;
assign pe_5_7_go = _guard3132;
assign pe_6_0_mul_ready =
  _guard3135 ? 1'd1 :
  _guard3138 ? 1'd0 :
  1'd0;
assign pe_6_0_clk = clk;
assign pe_6_0_top =
  _guard3151 ? top_6_0_out :
  32'd0;
assign pe_6_0_left =
  _guard3164 ? left_6_0_out :
  32'd0;
assign pe_6_0_reset = reset;
assign pe_6_0_go = _guard3177;
assign top_6_0_write_en = _guard3180;
assign top_6_0_clk = clk;
assign top_6_0_reset = reset;
assign top_6_0_in = top_5_0_out;
assign pe_6_1_mul_ready =
  _guard3186 ? 1'd1 :
  _guard3189 ? 1'd0 :
  1'd0;
assign pe_6_1_clk = clk;
assign pe_6_1_top =
  _guard3202 ? top_6_1_out :
  32'd0;
assign pe_6_1_left =
  _guard3215 ? left_6_1_out :
  32'd0;
assign pe_6_1_reset = reset;
assign pe_6_1_go = _guard3228;
assign left_7_5_write_en = _guard3231;
assign left_7_5_clk = clk;
assign left_7_5_reset = reset;
assign left_7_5_in = left_7_4_out;
assign index_lt_27_left = idx_add_out;
assign index_lt_27_right = 5'd27;
assign idx_between_21_22_reg_write_en = _guard3241;
assign idx_between_21_22_reg_clk = clk;
assign idx_between_21_22_reg_reset = reset;
assign idx_between_21_22_reg_in =
  _guard3242 ? idx_between_21_22_comb_out :
  _guard3245 ? 1'd0 :
  'x;
assign idx_between_22_23_reg_write_en = _guard3250;
assign idx_between_22_23_reg_clk = clk;
assign idx_between_22_23_reg_reset = reset;
assign idx_between_22_23_reg_in =
  _guard3253 ? 1'd0 :
  _guard3254 ? idx_between_22_23_comb_out :
  'x;
assign idx_between_1_9_comb_left = index_ge_1_out;
assign idx_between_1_9_comb_right = index_lt_9_out;
assign index_ge_25_left = idx_add_out;
assign index_ge_25_right = 5'd25;
assign idx_between_14_18_comb_left = index_ge_14_out;
assign idx_between_14_18_comb_right = index_lt_18_out;
assign idx_between_14_15_comb_left = index_ge_14_out;
assign idx_between_14_15_comb_right = index_lt_15_out;
assign idx_between_15_19_comb_left = index_ge_15_out;
assign idx_between_15_19_comb_right = index_lt_19_out;
assign idx_between_7_15_reg_write_en = _guard3269;
assign idx_between_7_15_reg_clk = clk;
assign idx_between_7_15_reg_reset = reset;
assign idx_between_7_15_reg_in =
  _guard3270 ? idx_between_7_15_comb_out :
  _guard3273 ? 1'd0 :
  'x;
assign index_ge_20_left = idx_add_out;
assign index_ge_20_right = 5'd20;
assign idx_between_16_17_reg_write_en = _guard3280;
assign idx_between_16_17_reg_clk = clk;
assign idx_between_16_17_reg_reset = reset;
assign idx_between_16_17_reg_in =
  _guard3283 ? 1'd0 :
  _guard3284 ? idx_between_16_17_comb_out :
  'x;
assign cond_wire18_in =
  _guard3287 ? cond18_out :
  _guard3288 ? idx_between_16_17_reg_out :
  1'd0;
assign cond19_write_en = _guard3289;
assign cond19_clk = clk;
assign cond19_reset = reset;
assign cond19_in =
  _guard3290 ? idx_between_4_12_reg_out :
  1'd0;
assign cond_wire29_in =
  _guard3291 ? idx_between_6_14_reg_out :
  _guard3294 ? cond29_out :
  1'd0;
assign cond34_write_en = _guard3295;
assign cond34_clk = clk;
assign cond34_reset = reset;
assign cond34_in =
  _guard3296 ? idx_between_7_15_reg_out :
  1'd0;
assign cond40_write_en = _guard3297;
assign cond40_clk = clk;
assign cond40_reset = reset;
assign cond40_in =
  _guard3298 ? idx_between_2_6_reg_out :
  1'd0;
assign cond57_write_en = _guard3299;
assign cond57_clk = clk;
assign cond57_reset = reset;
assign cond57_in =
  _guard3300 ? idx_between_6_14_reg_out :
  1'd0;
assign cond_wire59_in =
  _guard3301 ? idx_between_18_19_reg_out :
  _guard3304 ? cond59_out :
  1'd0;
assign cond_wire61_in =
  _guard3305 ? idx_between_7_15_reg_out :
  _guard3308 ? cond61_out :
  1'd0;
assign cond74_write_en = _guard3309;
assign cond74_clk = clk;
assign cond74_reset = reset;
assign cond74_in =
  _guard3310 ? idx_between_3_11_reg_out :
  1'd0;
assign cond95_write_en = _guard3311;
assign cond95_clk = clk;
assign cond95_reset = reset;
assign cond95_in =
  _guard3312 ? idx_between_12_20_reg_out :
  1'd0;
assign cond109_write_en = _guard3313;
assign cond109_clk = clk;
assign cond109_reset = reset;
assign cond109_in =
  _guard3314 ? idx_between_16_17_reg_out :
  1'd0;
assign cond_wire111_in =
  _guard3315 ? idx_between_5_13_reg_out :
  _guard3318 ? cond111_out :
  1'd0;
assign cond_wire112_in =
  _guard3321 ? cond112_out :
  _guard3322 ? idx_between_9_17_reg_out :
  1'd0;
assign cond_wire118_in =
  _guard3323 ? idx_between_7_11_reg_out :
  _guard3326 ? cond118_out :
  1'd0;
assign cond_wire137_in =
  _guard3327 ? idx_between_23_24_reg_out :
  _guard3330 ? cond137_out :
  1'd0;
assign cond158_write_en = _guard3331;
assign cond158_clk = clk;
assign cond158_reset = reset;
assign cond158_in =
  _guard3332 ? idx_between_21_22_reg_out :
  1'd0;
assign cond159_write_en = _guard3333;
assign cond159_clk = clk;
assign cond159_reset = reset;
assign cond159_in =
  _guard3334 ? idx_between_10_14_reg_out :
  1'd0;
assign cond162_write_en = _guard3335;
assign cond162_clk = clk;
assign cond162_reset = reset;
assign cond162_in =
  _guard3336 ? idx_between_22_23_reg_out :
  1'd0;
assign cond164_write_en = _guard3337;
assign cond164_clk = clk;
assign cond164_reset = reset;
assign cond164_in =
  _guard3338 ? idx_between_11_19_reg_out :
  1'd0;
assign cond166_write_en = _guard3339;
assign cond166_clk = clk;
assign cond166_reset = reset;
assign cond166_in =
  _guard3340 ? idx_between_23_24_reg_out :
  1'd0;
assign cond_wire170_in =
  _guard3341 ? idx_between_24_25_reg_out :
  _guard3344 ? cond170_out :
  1'd0;
assign cond_wire175_in =
  _guard3345 ? idx_between_18_19_reg_out :
  _guard3348 ? cond175_out :
  1'd0;
assign cond180_write_en = _guard3349;
assign cond180_clk = clk;
assign cond180_reset = reset;
assign cond180_in =
  _guard3350 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire197_in =
  _guard3353 ? cond197_out :
  _guard3354 ? idx_between_12_20_reg_out :
  1'd0;
assign cond198_write_en = _guard3355;
assign cond198_clk = clk;
assign cond198_reset = reset;
assign cond198_in =
  _guard3356 ? idx_between_16_24_reg_out :
  1'd0;
assign cond217_write_en = _guard3357;
assign cond217_clk = clk;
assign cond217_reset = reset;
assign cond217_in =
  _guard3358 ? idx_between_10_14_reg_out :
  1'd0;
assign cond222_write_en = _guard3359;
assign cond222_clk = clk;
assign cond222_reset = reset;
assign cond222_in =
  _guard3360 ? idx_between_11_19_reg_out :
  1'd0;
assign cond_wire222_in =
  _guard3361 ? idx_between_11_19_reg_out :
  _guard3364 ? cond222_out :
  1'd0;
assign cond_wire223_in =
  _guard3365 ? idx_between_15_23_reg_out :
  _guard3368 ? cond223_out :
  1'd0;
assign cond_wire225_in =
  _guard3371 ? cond225_out :
  _guard3372 ? idx_between_12_16_reg_out :
  1'd0;
assign cond_wire237_in =
  _guard3375 ? cond237_out :
  _guard3376 ? idx_between_7_15_reg_out :
  1'd0;
assign cond247_write_en = _guard3377;
assign cond247_clk = clk;
assign cond247_reset = reset;
assign cond247_in =
  _guard3378 ? idx_between_10_18_reg_out :
  1'd0;
assign cond_wire260_in =
  _guard3379 ? idx_between_17_25_reg_out :
  _guard3382 ? cond260_out :
  1'd0;
assign pe_0_2_mul_ready =
  _guard3385 ? 1'd1 :
  _guard3388 ? 1'd0 :
  1'd0;
assign pe_0_2_clk = clk;
assign pe_0_2_top =
  _guard3401 ? top_0_2_out :
  32'd0;
assign pe_0_2_left =
  _guard3414 ? left_0_2_out :
  32'd0;
assign pe_0_2_reset = reset;
assign pe_0_2_go = _guard3427;
assign pe_1_6_mul_ready =
  _guard3430 ? 1'd1 :
  _guard3433 ? 1'd0 :
  1'd0;
assign pe_1_6_clk = clk;
assign pe_1_6_top =
  _guard3446 ? top_1_6_out :
  32'd0;
assign pe_1_6_left =
  _guard3459 ? left_1_6_out :
  32'd0;
assign pe_1_6_reset = reset;
assign pe_1_6_go = _guard3472;
assign left_3_5_write_en = _guard3475;
assign left_3_5_clk = clk;
assign left_3_5_reset = reset;
assign left_3_5_in = left_3_4_out;
assign top_5_5_write_en = _guard3481;
assign top_5_5_clk = clk;
assign top_5_5_reset = reset;
assign top_5_5_in = top_4_5_out;
assign left_6_1_write_en = _guard3487;
assign left_6_1_clk = clk;
assign left_6_1_reset = reset;
assign left_6_1_in = left_6_0_out;
assign pe_6_5_mul_ready =
  _guard3493 ? 1'd1 :
  _guard3496 ? 1'd0 :
  1'd0;
assign pe_6_5_clk = clk;
assign pe_6_5_top =
  _guard3509 ? top_6_5_out :
  32'd0;
assign pe_6_5_left =
  _guard3522 ? left_6_5_out :
  32'd0;
assign pe_6_5_reset = reset;
assign pe_6_5_go = _guard3535;
assign left_6_7_write_en = _guard3538;
assign left_6_7_clk = clk;
assign left_6_7_reset = reset;
assign left_6_7_in = left_6_6_out;
assign pe_7_0_mul_ready =
  _guard3544 ? 1'd1 :
  _guard3547 ? 1'd0 :
  1'd0;
assign pe_7_0_clk = clk;
assign pe_7_0_top =
  _guard3560 ? top_7_0_out :
  32'd0;
assign pe_7_0_left =
  _guard3573 ? left_7_0_out :
  32'd0;
assign pe_7_0_reset = reset;
assign pe_7_0_go = _guard3586;
assign top_7_4_write_en = _guard3589;
assign top_7_4_clk = clk;
assign top_7_4_reset = reset;
assign top_7_4_in = top_6_4_out;
assign t0_idx_write_en = _guard3599;
assign t0_idx_clk = clk;
assign t0_idx_reset = reset;
assign t0_idx_in =
  _guard3602 ? 4'd0 :
  _guard3605 ? t0_add_out :
  'x;
assign t4_idx_write_en = _guard3612;
assign t4_idx_clk = clk;
assign t4_idx_reset = reset;
assign t4_idx_in =
  _guard3615 ? 4'd0 :
  _guard3618 ? t4_add_out :
  'x;
assign t6_idx_write_en = _guard3625;
assign t6_idx_clk = clk;
assign t6_idx_reset = reset;
assign t6_idx_in =
  _guard3628 ? 4'd0 :
  _guard3631 ? t6_add_out :
  'x;
assign l1_idx_write_en = _guard3638;
assign l1_idx_clk = clk;
assign l1_idx_reset = reset;
assign l1_idx_in =
  _guard3641 ? l1_add_out :
  _guard3644 ? 4'd0 :
  'x;
assign l5_add_left = 4'd1;
assign l5_add_right = l5_idx_out;
assign idx_add_left = idx_out;
assign idx_add_right = 5'd1;
assign index_lt_16_left = idx_add_out;
assign index_lt_16_right = 5'd16;
assign idx_between_12_16_comb_left = index_ge_12_out;
assign idx_between_12_16_comb_right = index_lt_16_out;
assign idx_between_4_12_reg_write_en = _guard3661;
assign idx_between_4_12_reg_clk = clk;
assign idx_between_4_12_reg_reset = reset;
assign idx_between_4_12_reg_in =
  _guard3662 ? idx_between_4_12_comb_out :
  _guard3665 ? 1'd0 :
  'x;
assign idx_between_21_22_comb_left = index_ge_21_out;
assign idx_between_21_22_comb_right = index_lt_22_out;
assign idx_between_8_12_reg_write_en = _guard3672;
assign idx_between_8_12_reg_clk = clk;
assign idx_between_8_12_reg_reset = reset;
assign idx_between_8_12_reg_in =
  _guard3675 ? 1'd0 :
  _guard3676 ? idx_between_8_12_comb_out :
  'x;
assign index_ge_7_left = idx_add_out;
assign index_ge_7_right = 5'd7;
assign idx_between_3_11_comb_left = index_ge_3_out;
assign idx_between_3_11_comb_right = index_lt_11_out;
assign cond3_write_en = _guard3681;
assign cond3_clk = clk;
assign cond3_reset = reset;
assign cond3_in =
  _guard3682 ? idx_between_13_14_reg_out :
  1'd0;
assign cond13_write_en = _guard3683;
assign cond13_clk = clk;
assign cond13_reset = reset;
assign cond13_in =
  _guard3684 ? idx_between_15_16_reg_out :
  1'd0;
assign cond29_write_en = _guard3685;
assign cond29_clk = clk;
assign cond29_reset = reset;
assign cond29_in =
  _guard3686 ? idx_between_6_14_reg_out :
  1'd0;
assign cond41_write_en = _guard3687;
assign cond41_clk = clk;
assign cond41_reset = reset;
assign cond41_in =
  _guard3688 ? idx_between_2_10_reg_out :
  1'd0;
assign cond54_write_en = _guard3689;
assign cond54_clk = clk;
assign cond54_reset = reset;
assign cond54_in =
  _guard3690 ? idx_between_9_17_reg_out :
  1'd0;
assign cond64_write_en = _guard3691;
assign cond64_clk = clk;
assign cond64_reset = reset;
assign cond64_in =
  _guard3692 ? idx_between_8_12_reg_out :
  1'd0;
assign cond67_write_en = _guard3693;
assign cond67_clk = clk;
assign cond67_reset = reset;
assign cond67_in =
  _guard3694 ? idx_between_20_21_reg_out :
  1'd0;
assign cond68_write_en = _guard3695;
assign cond68_clk = clk;
assign cond68_reset = reset;
assign cond68_in =
  _guard3696 ? idx_between_9_13_reg_out :
  1'd0;
assign cond77_write_en = _guard3697;
assign cond77_clk = clk;
assign cond77_reset = reset;
assign cond77_in =
  _guard3698 ? idx_between_4_8_reg_out :
  1'd0;
assign cond89_write_en = _guard3699;
assign cond89_clk = clk;
assign cond89_reset = reset;
assign cond89_in =
  _guard3700 ? idx_between_7_11_reg_out :
  1'd0;
assign cond94_write_en = _guard3701;
assign cond94_clk = clk;
assign cond94_reset = reset;
assign cond94_in =
  _guard3702 ? idx_between_8_16_reg_out :
  1'd0;
assign cond_wire125_in =
  _guard3703 ? idx_between_20_21_reg_out :
  _guard3706 ? cond125_out :
  1'd0;
assign cond128_write_en = _guard3707;
assign cond128_clk = clk;
assign cond128_reset = reset;
assign cond128_in =
  _guard3708 ? idx_between_13_21_reg_out :
  1'd0;
assign cond131_write_en = _guard3709;
assign cond131_clk = clk;
assign cond131_reset = reset;
assign cond131_in =
  _guard3710 ? idx_between_10_18_reg_out :
  1'd0;
assign cond132_write_en = _guard3711;
assign cond132_clk = clk;
assign cond132_reset = reset;
assign cond132_in =
  _guard3712 ? idx_between_14_22_reg_out :
  1'd0;
assign cond_wire132_in =
  _guard3715 ? cond132_out :
  _guard3716 ? idx_between_14_22_reg_out :
  1'd0;
assign cond134_write_en = _guard3717;
assign cond134_clk = clk;
assign cond134_reset = reset;
assign cond134_in =
  _guard3718 ? idx_between_11_15_reg_out :
  1'd0;
assign cond136_write_en = _guard3719;
assign cond136_clk = clk;
assign cond136_reset = reset;
assign cond136_in =
  _guard3720 ? idx_between_15_23_reg_out :
  1'd0;
assign cond139_write_en = _guard3721;
assign cond139_clk = clk;
assign cond139_reset = reset;
assign cond139_in =
  _guard3722 ? idx_between_5_9_reg_out :
  1'd0;
assign cond140_write_en = _guard3723;
assign cond140_clk = clk;
assign cond140_reset = reset;
assign cond140_in =
  _guard3724 ? idx_between_5_13_reg_out :
  1'd0;
assign cond_wire142_in =
  _guard3725 ? idx_between_17_18_reg_out :
  _guard3728 ? cond142_out :
  1'd0;
assign cond_wire148_in =
  _guard3729 ? idx_between_7_15_reg_out :
  _guard3732 ? cond148_out :
  1'd0;
assign cond_wire151_in =
  _guard3735 ? cond151_out :
  _guard3736 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire161_in =
  _guard3739 ? cond161_out :
  _guard3740 ? idx_between_14_22_reg_out :
  1'd0;
assign cond_wire162_in =
  _guard3741 ? idx_between_22_23_reg_out :
  _guard3744 ? cond162_out :
  1'd0;
assign cond_wire165_in =
  _guard3745 ? idx_between_15_23_reg_out :
  _guard3748 ? cond165_out :
  1'd0;
assign cond_wire171_in =
  _guard3749 ? idx_between_5_13_reg_out :
  _guard3752 ? cond171_out :
  1'd0;
assign cond172_write_en = _guard3753;
assign cond172_clk = clk;
assign cond172_reset = reset;
assign cond172_in =
  _guard3754 ? idx_between_6_10_reg_out :
  1'd0;
assign cond_wire177_in =
  _guard3757 ? cond177_out :
  _guard3758 ? idx_between_7_15_reg_out :
  1'd0;
assign cond183_write_en = _guard3759;
assign cond183_clk = clk;
assign cond183_reset = reset;
assign cond183_in =
  _guard3760 ? idx_between_20_21_reg_out :
  1'd0;
assign cond187_write_en = _guard3761;
assign cond187_clk = clk;
assign cond187_reset = reset;
assign cond187_in =
  _guard3762 ? idx_between_21_22_reg_out :
  1'd0;
assign cond190_write_en = _guard3763;
assign cond190_clk = clk;
assign cond190_reset = reset;
assign cond190_in =
  _guard3764 ? idx_between_14_22_reg_out :
  1'd0;
assign cond191_write_en = _guard3765;
assign cond191_clk = clk;
assign cond191_reset = reset;
assign cond191_in =
  _guard3766 ? idx_between_22_23_reg_out :
  1'd0;
assign cond223_write_en = _guard3767;
assign cond223_clk = clk;
assign cond223_reset = reset;
assign cond223_in =
  _guard3768 ? idx_between_15_23_reg_out :
  1'd0;
assign cond238_write_en = _guard3769;
assign cond238_clk = clk;
assign cond238_reset = reset;
assign cond238_in =
  _guard3770 ? idx_between_8_12_reg_out :
  1'd0;
assign cond244_write_en = _guard3771;
assign cond244_clk = clk;
assign cond244_reset = reset;
assign cond244_in =
  _guard3772 ? idx_between_13_21_reg_out :
  1'd0;
assign cond_wire252_in =
  _guard3773 ? idx_between_15_23_reg_out :
  _guard3776 ? cond252_out :
  1'd0;
assign cond_wire262_in =
  _guard3777 ? idx_between_14_18_reg_out :
  _guard3780 ? cond262_out :
  1'd0;
assign cond_wire264_in =
  _guard3783 ? cond264_out :
  _guard3784 ? idx_between_18_26_reg_out :
  1'd0;
assign cond265_write_en = _guard3785;
assign cond265_clk = clk;
assign cond265_reset = reset;
assign cond265_in =
  _guard3786 ? idx_between_26_27_reg_out :
  1'd0;
assign cond_wire267_in =
  _guard3787 ? idx_between_19_27_reg_out :
  _guard3790 ? cond267_out :
  1'd0;
assign early_reset_static_par0_done_in = ud0_out;
assign left_0_7_write_en = _guard3793;
assign left_0_7_clk = clk;
assign left_0_7_reset = reset;
assign left_0_7_in = left_0_6_out;
assign pe_2_1_mul_ready =
  _guard3799 ? 1'd1 :
  _guard3802 ? 1'd0 :
  1'd0;
assign pe_2_1_clk = clk;
assign pe_2_1_top =
  _guard3815 ? top_2_1_out :
  32'd0;
assign pe_2_1_left =
  _guard3828 ? left_2_1_out :
  32'd0;
assign pe_2_1_reset = reset;
assign pe_2_1_go = _guard3841;
assign pe_2_3_mul_ready =
  _guard3844 ? 1'd1 :
  _guard3847 ? 1'd0 :
  1'd0;
assign pe_2_3_clk = clk;
assign pe_2_3_top =
  _guard3860 ? top_2_3_out :
  32'd0;
assign pe_2_3_left =
  _guard3873 ? left_2_3_out :
  32'd0;
assign pe_2_3_reset = reset;
assign pe_2_3_go = _guard3886;
assign pe_2_5_mul_ready =
  _guard3889 ? 1'd1 :
  _guard3892 ? 1'd0 :
  1'd0;
assign pe_2_5_clk = clk;
assign pe_2_5_top =
  _guard3905 ? top_2_5_out :
  32'd0;
assign pe_2_5_left =
  _guard3918 ? left_2_5_out :
  32'd0;
assign pe_2_5_reset = reset;
assign pe_2_5_go = _guard3931;
assign pe_3_1_mul_ready =
  _guard3934 ? 1'd1 :
  _guard3937 ? 1'd0 :
  1'd0;
assign pe_3_1_clk = clk;
assign pe_3_1_top =
  _guard3950 ? top_3_1_out :
  32'd0;
assign pe_3_1_left =
  _guard3963 ? left_3_1_out :
  32'd0;
assign pe_3_1_reset = reset;
assign pe_3_1_go = _guard3976;
assign top_3_4_write_en = _guard3979;
assign top_3_4_clk = clk;
assign top_3_4_reset = reset;
assign top_3_4_in = top_2_4_out;
assign pe_5_3_mul_ready =
  _guard3985 ? 1'd1 :
  _guard3988 ? 1'd0 :
  1'd0;
assign pe_5_3_clk = clk;
assign pe_5_3_top =
  _guard4001 ? top_5_3_out :
  32'd0;
assign pe_5_3_left =
  _guard4014 ? left_5_3_out :
  32'd0;
assign pe_5_3_reset = reset;
assign pe_5_3_go = _guard4027;
assign pe_5_5_mul_ready =
  _guard4030 ? 1'd1 :
  _guard4033 ? 1'd0 :
  1'd0;
assign pe_5_5_clk = clk;
assign pe_5_5_top =
  _guard4046 ? top_5_5_out :
  32'd0;
assign pe_5_5_left =
  _guard4059 ? left_5_5_out :
  32'd0;
assign pe_5_5_reset = reset;
assign pe_5_5_go = _guard4072;
assign pe_6_2_mul_ready =
  _guard4075 ? 1'd1 :
  _guard4078 ? 1'd0 :
  1'd0;
assign pe_6_2_clk = clk;
assign pe_6_2_top =
  _guard4091 ? top_6_2_out :
  32'd0;
assign pe_6_2_left =
  _guard4104 ? left_6_2_out :
  32'd0;
assign pe_6_2_reset = reset;
assign pe_6_2_go = _guard4117;
assign pe_6_3_mul_ready =
  _guard4120 ? 1'd1 :
  _guard4123 ? 1'd0 :
  1'd0;
assign pe_6_3_clk = clk;
assign pe_6_3_top =
  _guard4136 ? top_6_3_out :
  32'd0;
assign pe_6_3_left =
  _guard4149 ? left_6_3_out :
  32'd0;
assign pe_6_3_reset = reset;
assign pe_6_3_go = _guard4162;
assign left_7_1_write_en = _guard4165;
assign left_7_1_clk = clk;
assign left_7_1_reset = reset;
assign left_7_1_in = left_7_0_out;
assign left_7_3_write_en = _guard4171;
assign left_7_3_clk = clk;
assign left_7_3_reset = reset;
assign left_7_3_in = left_7_2_out;
assign top_7_5_write_en = _guard4177;
assign top_7_5_clk = clk;
assign top_7_5_reset = reset;
assign top_7_5_in = top_6_5_out;
assign t4_add_left = 4'd1;
assign t4_add_right = t4_idx_out;
assign t5_idx_write_en = _guard4193;
assign t5_idx_clk = clk;
assign t5_idx_reset = reset;
assign t5_idx_in =
  _guard4196 ? 4'd0 :
  _guard4199 ? t5_add_out :
  'x;
assign t6_add_left = 4'd1;
assign t6_add_right = t6_idx_out;
assign idx_between_4_12_comb_left = index_ge_4_out;
assign idx_between_4_12_comb_right = index_lt_12_out;
assign index_ge_17_left = idx_add_out;
assign index_ge_17_right = 5'd17;
assign idx_between_27_28_reg_write_en = _guard4214;
assign idx_between_27_28_reg_clk = clk;
assign idx_between_27_28_reg_reset = reset;
assign idx_between_27_28_reg_in =
  _guard4217 ? 1'd0 :
  _guard4218 ? idx_between_27_28_comb_out :
  'x;
assign idx_between_13_17_comb_left = index_ge_13_out;
assign idx_between_13_17_comb_right = index_lt_17_out;
assign idx_between_14_18_reg_write_en = _guard4225;
assign idx_between_14_18_reg_clk = clk;
assign idx_between_14_18_reg_reset = reset;
assign idx_between_14_18_reg_in =
  _guard4226 ? idx_between_14_18_comb_out :
  _guard4229 ? 1'd0 :
  'x;
assign index_lt_24_left = idx_add_out;
assign index_lt_24_right = 5'd24;
assign idx_between_19_20_reg_write_en = _guard4236;
assign idx_between_19_20_reg_clk = clk;
assign idx_between_19_20_reg_reset = reset;
assign idx_between_19_20_reg_in =
  _guard4239 ? 1'd0 :
  _guard4240 ? idx_between_19_20_comb_out :
  'x;
assign cond17_write_en = _guard4241;
assign cond17_clk = clk;
assign cond17_reset = reset;
assign cond17_in =
  _guard4242 ? idx_between_8_16_reg_out :
  1'd0;
assign cond_wire22_in =
  _guard4245 ? cond22_out :
  _guard4246 ? idx_between_9_17_reg_out :
  1'd0;
assign cond23_write_en = _guard4247;
assign cond23_clk = clk;
assign cond23_reset = reset;
assign cond23_in =
  _guard4248 ? idx_between_17_18_reg_out :
  1'd0;
assign cond25_write_en = _guard4249;
assign cond25_clk = clk;
assign cond25_reset = reset;
assign cond25_in =
  _guard4250 ? idx_between_6_10_reg_out :
  1'd0;
assign cond_wire33_in =
  _guard4251 ? idx_between_19_20_reg_out :
  _guard4254 ? cond33_out :
  1'd0;
assign cond52_write_en = _guard4255;
assign cond52_clk = clk;
assign cond52_reset = reset;
assign cond52_in =
  _guard4256 ? idx_between_5_9_reg_out :
  1'd0;
assign cond56_write_en = _guard4257;
assign cond56_clk = clk;
assign cond56_reset = reset;
assign cond56_in =
  _guard4258 ? idx_between_6_10_reg_out :
  1'd0;
assign cond58_write_en = _guard4259;
assign cond58_clk = clk;
assign cond58_reset = reset;
assign cond58_in =
  _guard4260 ? idx_between_10_18_reg_out :
  1'd0;
assign cond75_write_en = _guard4261;
assign cond75_clk = clk;
assign cond75_reset = reset;
assign cond75_in =
  _guard4262 ? idx_between_7_15_reg_out :
  1'd0;
assign cond88_write_en = _guard4263;
assign cond88_clk = clk;
assign cond88_reset = reset;
assign cond88_in =
  _guard4264 ? idx_between_18_19_reg_out :
  1'd0;
assign cond93_write_en = _guard4265;
assign cond93_clk = clk;
assign cond93_reset = reset;
assign cond93_in =
  _guard4266 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire98_in =
  _guard4269 ? cond98_out :
  _guard4270 ? idx_between_9_17_reg_out :
  1'd0;
assign cond_wire106_in =
  _guard4271 ? idx_between_4_8_reg_out :
  _guard4274 ? cond106_out :
  1'd0;
assign cond_wire120_in =
  _guard4275 ? idx_between_11_19_reg_out :
  _guard4278 ? cond120_out :
  1'd0;
assign cond124_write_en = _guard4279;
assign cond124_clk = clk;
assign cond124_reset = reset;
assign cond124_in =
  _guard4280 ? idx_between_12_20_reg_out :
  1'd0;
assign cond137_write_en = _guard4281;
assign cond137_clk = clk;
assign cond137_reset = reset;
assign cond137_in =
  _guard4282 ? idx_between_23_24_reg_out :
  1'd0;
assign cond155_write_en = _guard4283;
assign cond155_clk = clk;
assign cond155_reset = reset;
assign cond155_in =
  _guard4284 ? idx_between_9_13_reg_out :
  1'd0;
assign cond_wire176_in =
  _guard4285 ? idx_between_7_11_reg_out :
  _guard4288 ? cond176_out :
  1'd0;
assign cond188_write_en = _guard4289;
assign cond188_clk = clk;
assign cond188_reset = reset;
assign cond188_in =
  _guard4290 ? idx_between_10_14_reg_out :
  1'd0;
assign cond209_write_en = _guard4291;
assign cond209_clk = clk;
assign cond209_reset = reset;
assign cond209_in =
  _guard4292 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire213_in =
  _guard4293 ? idx_between_9_13_reg_out :
  _guard4296 ? cond213_out :
  1'd0;
assign cond220_write_en = _guard4297;
assign cond220_clk = clk;
assign cond220_reset = reset;
assign cond220_in =
  _guard4298 ? idx_between_22_23_reg_out :
  1'd0;
assign cond_wire221_in =
  _guard4301 ? cond221_out :
  _guard4302 ? idx_between_11_15_reg_out :
  1'd0;
assign cond228_write_en = _guard4303;
assign cond228_clk = clk;
assign cond228_reset = reset;
assign cond228_in =
  _guard4304 ? idx_between_24_25_reg_out :
  1'd0;
assign cond232_write_en = _guard4305;
assign cond232_clk = clk;
assign cond232_reset = reset;
assign cond232_in =
  _guard4306 ? idx_between_25_26_reg_out :
  1'd0;
assign cond_wire236_in =
  _guard4307 ? idx_between_26_27_reg_out :
  _guard4310 ? cond236_out :
  1'd0;
assign cond258_write_en = _guard4311;
assign cond258_clk = clk;
assign cond258_reset = reset;
assign cond258_in =
  _guard4312 ? idx_between_13_17_reg_out :
  1'd0;
assign cond262_write_en = _guard4313;
assign cond262_clk = clk;
assign cond262_reset = reset;
assign cond262_in =
  _guard4314 ? idx_between_14_18_reg_out :
  1'd0;
assign fsm0_write_en = _guard4315;
assign fsm0_clk = clk;
assign fsm0_reset = reset;
assign fsm0_in =
  _guard4318 ? adder_out :
  _guard4321 ? 5'd0 :
  5'd0;
assign pe_1_5_mul_ready =
  _guard4324 ? 1'd1 :
  _guard4327 ? 1'd0 :
  1'd0;
assign pe_1_5_clk = clk;
assign pe_1_5_top =
  _guard4340 ? top_1_5_out :
  32'd0;
assign pe_1_5_left =
  _guard4353 ? left_1_5_out :
  32'd0;
assign pe_1_5_reset = reset;
assign pe_1_5_go = _guard4366;
assign top_1_6_write_en = _guard4369;
assign top_1_6_clk = clk;
assign top_1_6_reset = reset;
assign top_1_6_in = top_0_6_out;
assign top_2_0_write_en = _guard4375;
assign top_2_0_clk = clk;
assign top_2_0_reset = reset;
assign top_2_0_in = top_1_0_out;
assign top_3_0_write_en = _guard4381;
assign top_3_0_clk = clk;
assign top_3_0_reset = reset;
assign top_3_0_in = top_2_0_out;
assign top_3_1_write_en = _guard4387;
assign top_3_1_clk = clk;
assign top_3_1_reset = reset;
assign top_3_1_in = top_2_1_out;
assign pe_4_6_mul_ready =
  _guard4393 ? 1'd1 :
  _guard4396 ? 1'd0 :
  1'd0;
assign pe_4_6_clk = clk;
assign pe_4_6_top =
  _guard4409 ? top_4_6_out :
  32'd0;
assign pe_4_6_left =
  _guard4422 ? left_4_6_out :
  32'd0;
assign pe_4_6_reset = reset;
assign pe_4_6_go = _guard4435;
assign top_5_2_write_en = _guard4438;
assign top_5_2_clk = clk;
assign top_5_2_reset = reset;
assign top_5_2_in = top_4_2_out;
assign top_5_4_write_en = _guard4444;
assign top_5_4_clk = clk;
assign top_5_4_reset = reset;
assign top_5_4_in = top_4_4_out;
assign left_7_7_write_en = _guard4450;
assign left_7_7_clk = clk;
assign left_7_7_reset = reset;
assign left_7_7_in = left_7_6_out;
assign t7_add_left = 4'd1;
assign t7_add_right = t7_idx_out;
assign l4_idx_write_en = _guard4466;
assign l4_idx_clk = clk;
assign l4_idx_reset = reset;
assign l4_idx_in =
  _guard4469 ? 4'd0 :
  _guard4472 ? l4_add_out :
  'x;
assign idx_write_en = _guard4477;
assign idx_clk = clk;
assign idx_reset = reset;
assign idx_in =
  _guard4480 ? 5'd0 :
  _guard4481 ? idx_add_out :
  'x;
assign index_ge_21_left = idx_add_out;
assign index_ge_21_right = 5'd21;
assign idx_between_14_22_comb_left = index_ge_14_out;
assign idx_between_14_22_comb_right = index_lt_22_out;
assign idx_between_10_18_reg_write_en = _guard4490;
assign idx_between_10_18_reg_clk = clk;
assign idx_between_10_18_reg_reset = reset;
assign idx_between_10_18_reg_in =
  _guard4493 ? 1'd0 :
  _guard4494 ? idx_between_10_18_comb_out :
  'x;
assign idx_between_5_9_reg_write_en = _guard4499;
assign idx_between_5_9_reg_clk = clk;
assign idx_between_5_9_reg_reset = reset;
assign idx_between_5_9_reg_in =
  _guard4500 ? idx_between_5_9_comb_out :
  _guard4503 ? 1'd0 :
  'x;
assign index_lt_15_left = idx_add_out;
assign index_lt_15_right = 5'd15;
assign cond7_write_en = _guard4506;
assign cond7_clk = clk;
assign cond7_reset = reset;
assign cond7_in =
  _guard4507 ? idx_between_6_14_reg_out :
  1'd0;
assign cond_wire8_in =
  _guard4508 ? idx_between_14_15_reg_out :
  _guard4511 ? cond8_out :
  1'd0;
assign cond9_write_en = _guard4512;
assign cond9_clk = clk;
assign cond9_reset = reset;
assign cond9_in =
  _guard4513 ? idx_between_2_10_reg_out :
  1'd0;
assign cond14_write_en = _guard4514;
assign cond14_clk = clk;
assign cond14_reset = reset;
assign cond14_in =
  _guard4515 ? idx_between_3_11_reg_out :
  1'd0;
assign cond_wire20_in =
  _guard4516 ? idx_between_5_9_reg_out :
  _guard4519 ? cond20_out :
  1'd0;
assign cond27_write_en = _guard4520;
assign cond27_clk = clk;
assign cond27_reset = reset;
assign cond27_in =
  _guard4521 ? idx_between_10_18_reg_out :
  1'd0;
assign cond32_write_en = _guard4522;
assign cond32_clk = clk;
assign cond32_reset = reset;
assign cond32_in =
  _guard4523 ? idx_between_11_19_reg_out :
  1'd0;
assign cond_wire37_in =
  _guard4526 ? cond37_out :
  _guard4527 ? idx_between_12_20_reg_out :
  1'd0;
assign cond50_write_en = _guard4528;
assign cond50_clk = clk;
assign cond50_reset = reset;
assign cond50_in =
  _guard4529 ? idx_between_8_16_reg_out :
  1'd0;
assign cond_wire60_in =
  _guard4530 ? idx_between_7_11_reg_out :
  _guard4533 ? cond60_out :
  1'd0;
assign cond_wire64_in =
  _guard4534 ? idx_between_8_12_reg_out :
  _guard4537 ? cond64_out :
  1'd0;
assign cond_wire81_in =
  _guard4540 ? cond81_out :
  _guard4541 ? idx_between_5_9_reg_out :
  1'd0;
assign cond_wire82_in =
  _guard4542 ? idx_between_5_13_reg_out :
  _guard4545 ? cond82_out :
  1'd0;
assign cond83_write_en = _guard4546;
assign cond83_clk = clk;
assign cond83_reset = reset;
assign cond83_in =
  _guard4547 ? idx_between_9_17_reg_out :
  1'd0;
assign cond_wire86_in =
  _guard4548 ? idx_between_6_14_reg_out :
  _guard4551 ? cond86_out :
  1'd0;
assign cond_wire87_in =
  _guard4552 ? idx_between_10_18_reg_out :
  _guard4555 ? cond87_out :
  1'd0;
assign cond91_write_en = _guard4556;
assign cond91_clk = clk;
assign cond91_reset = reset;
assign cond91_in =
  _guard4557 ? idx_between_11_19_reg_out :
  1'd0;
assign cond_wire105_in =
  _guard4560 ? cond105_out :
  _guard4561 ? idx_between_3_11_reg_out :
  1'd0;
assign cond116_write_en = _guard4562;
assign cond116_clk = clk;
assign cond116_reset = reset;
assign cond116_in =
  _guard4563 ? idx_between_10_18_reg_out :
  1'd0;
assign cond_wire117_in =
  _guard4564 ? idx_between_18_19_reg_out :
  _guard4567 ? cond117_out :
  1'd0;
assign cond_wire138_in =
  _guard4568 ? idx_between_4_12_reg_out :
  _guard4571 ? cond138_out :
  1'd0;
assign cond_wire140_in =
  _guard4572 ? idx_between_5_13_reg_out :
  _guard4575 ? cond140_out :
  1'd0;
assign cond_wire156_in =
  _guard4578 ? cond156_out :
  _guard4579 ? idx_between_9_17_reg_out :
  1'd0;
assign cond161_write_en = _guard4580;
assign cond161_clk = clk;
assign cond161_reset = reset;
assign cond161_in =
  _guard4581 ? idx_between_14_22_reg_out :
  1'd0;
assign cond174_write_en = _guard4582;
assign cond174_clk = clk;
assign cond174_reset = reset;
assign cond174_in =
  _guard4583 ? idx_between_10_18_reg_out :
  1'd0;
assign cond176_write_en = _guard4584;
assign cond176_clk = clk;
assign cond176_reset = reset;
assign cond176_in =
  _guard4585 ? idx_between_7_11_reg_out :
  1'd0;
assign cond_wire187_in =
  _guard4586 ? idx_between_21_22_reg_out :
  _guard4589 ? cond187_out :
  1'd0;
assign cond_wire190_in =
  _guard4592 ? cond190_out :
  _guard4593 ? idx_between_14_22_reg_out :
  1'd0;
assign cond194_write_en = _guard4594;
assign cond194_clk = clk;
assign cond194_reset = reset;
assign cond194_in =
  _guard4595 ? idx_between_15_23_reg_out :
  1'd0;
assign cond201_write_en = _guard4596;
assign cond201_clk = clk;
assign cond201_reset = reset;
assign cond201_in =
  _guard4597 ? idx_between_13_21_reg_out :
  1'd0;
assign cond205_write_en = _guard4598;
assign cond205_clk = clk;
assign cond205_reset = reset;
assign cond205_in =
  _guard4599 ? idx_between_7_11_reg_out :
  1'd0;
assign cond_wire207_in =
  _guard4600 ? idx_between_11_19_reg_out :
  _guard4603 ? cond207_out :
  1'd0;
assign cond_wire209_in =
  _guard4604 ? idx_between_8_12_reg_out :
  _guard4607 ? cond209_out :
  1'd0;
assign cond219_write_en = _guard4608;
assign cond219_clk = clk;
assign cond219_reset = reset;
assign cond219_in =
  _guard4609 ? idx_between_14_22_reg_out :
  1'd0;
assign cond221_write_en = _guard4610;
assign cond221_clk = clk;
assign cond221_reset = reset;
assign cond221_in =
  _guard4611 ? idx_between_11_15_reg_out :
  1'd0;
assign cond225_write_en = _guard4612;
assign cond225_clk = clk;
assign cond225_reset = reset;
assign cond225_in =
  _guard4613 ? idx_between_12_16_reg_out :
  1'd0;
assign cond256_write_en = _guard4614;
assign cond256_clk = clk;
assign cond256_reset = reset;
assign cond256_in =
  _guard4615 ? idx_between_16_24_reg_out :
  1'd0;
assign wrapper_early_reset_static_seq_done_in = _guard4618;
assign top_0_1_write_en = _guard4621;
assign top_0_1_clk = clk;
assign top_0_1_reset = reset;
assign top_0_1_in = t1_read_data;
assign left_0_2_write_en = _guard4627;
assign left_0_2_clk = clk;
assign left_0_2_reset = reset;
assign left_0_2_in = left_0_1_out;
assign pe_0_4_mul_ready =
  _guard4633 ? 1'd1 :
  _guard4636 ? 1'd0 :
  1'd0;
assign pe_0_4_clk = clk;
assign pe_0_4_top =
  _guard4649 ? top_0_4_out :
  32'd0;
assign pe_0_4_left =
  _guard4662 ? left_0_4_out :
  32'd0;
assign pe_0_4_reset = reset;
assign pe_0_4_go = _guard4675;
assign top_2_3_write_en = _guard4678;
assign top_2_3_clk = clk;
assign top_2_3_reset = reset;
assign top_2_3_in = top_1_3_out;
assign pe_2_6_mul_ready =
  _guard4684 ? 1'd1 :
  _guard4687 ? 1'd0 :
  1'd0;
assign pe_2_6_clk = clk;
assign pe_2_6_top =
  _guard4700 ? top_2_6_out :
  32'd0;
assign pe_2_6_left =
  _guard4713 ? left_2_6_out :
  32'd0;
assign pe_2_6_reset = reset;
assign pe_2_6_go = _guard4726;
assign left_3_0_write_en = _guard4729;
assign left_3_0_clk = clk;
assign left_3_0_reset = reset;
assign left_3_0_in = l3_read_data;
assign pe_4_2_mul_ready =
  _guard4735 ? 1'd1 :
  _guard4738 ? 1'd0 :
  1'd0;
assign pe_4_2_clk = clk;
assign pe_4_2_top =
  _guard4751 ? top_4_2_out :
  32'd0;
assign pe_4_2_left =
  _guard4764 ? left_4_2_out :
  32'd0;
assign pe_4_2_reset = reset;
assign pe_4_2_go = _guard4777;
assign top_5_1_write_en = _guard4780;
assign top_5_1_clk = clk;
assign top_5_1_reset = reset;
assign top_5_1_in = top_4_1_out;
assign left_5_4_write_en = _guard4786;
assign left_5_4_clk = clk;
assign left_5_4_reset = reset;
assign left_5_4_in = left_5_3_out;
assign pe_6_7_mul_ready =
  _guard4792 ? 1'd1 :
  _guard4795 ? 1'd0 :
  1'd0;
assign pe_6_7_clk = clk;
assign pe_6_7_top =
  _guard4808 ? top_6_7_out :
  32'd0;
assign pe_6_7_left =
  _guard4821 ? left_6_7_out :
  32'd0;
assign pe_6_7_reset = reset;
assign pe_6_7_go = _guard4834;
assign l7_add_left = 4'd1;
assign l7_add_right = l7_idx_out;
assign idx_between_18_26_reg_write_en = _guard4845;
assign idx_between_18_26_reg_clk = clk;
assign idx_between_18_26_reg_reset = reset;
assign idx_between_18_26_reg_in =
  _guard4846 ? idx_between_18_26_comb_out :
  _guard4849 ? 1'd0 :
  'x;
assign idx_between_3_7_comb_left = index_ge_3_out;
assign idx_between_3_7_comb_right = index_lt_7_out;
assign index_ge_4_left = idx_add_out;
assign index_ge_4_right = 5'd4;
assign idx_between_0_8_reg_write_en = _guard4858;
assign idx_between_0_8_reg_clk = clk;
assign idx_between_0_8_reg_reset = reset;
assign idx_between_0_8_reg_in =
  _guard4861 ? 1'd1 :
  _guard4862 ? index_lt_8_out :
  'x;
assign index_lt_8_left = idx_add_out;
assign index_lt_8_right = 5'd8;
assign index_lt_9_left = idx_add_out;
assign index_lt_9_right = 5'd9;
assign index_ge_1_left = idx_add_out;
assign index_ge_1_right = 5'd1;
assign idx_between_13_14_comb_left = index_ge_13_out;
assign idx_between_13_14_comb_right = index_lt_14_out;
assign idx_between_14_15_reg_write_en = _guard4875;
assign idx_between_14_15_reg_clk = clk;
assign idx_between_14_15_reg_reset = reset;
assign idx_between_14_15_reg_in =
  _guard4876 ? idx_between_14_15_comb_out :
  _guard4879 ? 1'd0 :
  'x;
assign idx_between_1_5_reg_write_en = _guard4884;
assign idx_between_1_5_reg_clk = clk;
assign idx_between_1_5_reg_reset = reset;
assign idx_between_1_5_reg_in =
  _guard4887 ? 1'd0 :
  _guard4888 ? idx_between_1_5_comb_out :
  'x;
assign idx_between_24_25_reg_write_en = _guard4893;
assign idx_between_24_25_reg_clk = clk;
assign idx_between_24_25_reg_reset = reset;
assign idx_between_24_25_reg_in =
  _guard4894 ? idx_between_24_25_comb_out :
  _guard4897 ? 1'd0 :
  'x;
assign idx_between_7_15_comb_left = index_ge_7_out;
assign idx_between_7_15_comb_right = index_lt_15_out;
assign idx_between_8_16_reg_write_en = _guard4904;
assign idx_between_8_16_reg_clk = clk;
assign idx_between_8_16_reg_reset = reset;
assign idx_between_8_16_reg_in =
  _guard4905 ? idx_between_8_16_comb_out :
  _guard4908 ? 1'd0 :
  'x;
assign index_lt_6_left = idx_add_out;
assign index_lt_6_right = 5'd6;
assign cond4_write_en = _guard4911;
assign cond4_clk = clk;
assign cond4_reset = reset;
assign cond4_in =
  _guard4912 ? idx_between_1_9_reg_out :
  1'd0;
assign cond5_write_en = _guard4913;
assign cond5_clk = clk;
assign cond5_reset = reset;
assign cond5_in =
  _guard4914 ? idx_between_2_6_reg_out :
  1'd0;
assign cond_wire6_in =
  _guard4917 ? cond6_out :
  _guard4918 ? idx_between_2_10_reg_out :
  1'd0;
assign cond20_write_en = _guard4919;
assign cond20_clk = clk;
assign cond20_reset = reset;
assign cond20_in =
  _guard4920 ? idx_between_5_9_reg_out :
  1'd0;
assign cond_wire36_in =
  _guard4921 ? idx_between_8_16_reg_out :
  _guard4924 ? cond36_out :
  1'd0;
assign cond46_write_en = _guard4925;
assign cond46_clk = clk;
assign cond46_reset = reset;
assign cond46_in =
  _guard4926 ? idx_between_7_15_reg_out :
  1'd0;
assign cond_wire62_in =
  _guard4927 ? idx_between_11_19_reg_out :
  _guard4930 ? cond62_out :
  1'd0;
assign cond63_write_en = _guard4931;
assign cond63_clk = clk;
assign cond63_reset = reset;
assign cond63_in =
  _guard4932 ? idx_between_19_20_reg_out :
  1'd0;
assign cond_wire66_in =
  _guard4935 ? cond66_out :
  _guard4936 ? idx_between_12_20_reg_out :
  1'd0;
assign cond_wire74_in =
  _guard4939 ? cond74_out :
  _guard4940 ? idx_between_3_11_reg_out :
  1'd0;
assign cond_wire75_in =
  _guard4941 ? idx_between_7_15_reg_out :
  _guard4944 ? cond75_out :
  1'd0;
assign cond78_write_en = _guard4945;
assign cond78_clk = clk;
assign cond78_reset = reset;
assign cond78_in =
  _guard4946 ? idx_between_4_12_reg_out :
  1'd0;
assign cond90_write_en = _guard4947;
assign cond90_clk = clk;
assign cond90_reset = reset;
assign cond90_in =
  _guard4948 ? idx_between_7_15_reg_out :
  1'd0;
assign cond_wire92_in =
  _guard4951 ? cond92_out :
  _guard4952 ? idx_between_19_20_reg_out :
  1'd0;
assign cond101_write_en = _guard4953;
assign cond101_clk = clk;
assign cond101_reset = reset;
assign cond101_in =
  _guard4954 ? idx_between_10_14_reg_out :
  1'd0;
assign cond106_write_en = _guard4955;
assign cond106_clk = clk;
assign cond106_reset = reset;
assign cond106_in =
  _guard4956 ? idx_between_4_8_reg_out :
  1'd0;
assign cond_wire108_in =
  _guard4957 ? idx_between_8_16_reg_out :
  _guard4960 ? cond108_out :
  1'd0;
assign cond112_write_en = _guard4961;
assign cond112_clk = clk;
assign cond112_reset = reset;
assign cond112_in =
  _guard4962 ? idx_between_9_17_reg_out :
  1'd0;
assign cond122_write_en = _guard4963;
assign cond122_clk = clk;
assign cond122_reset = reset;
assign cond122_in =
  _guard4964 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire122_in =
  _guard4965 ? idx_between_8_12_reg_out :
  _guard4968 ? cond122_out :
  1'd0;
assign cond_wire128_in =
  _guard4971 ? cond128_out :
  _guard4972 ? idx_between_13_21_reg_out :
  1'd0;
assign cond_wire139_in =
  _guard4975 ? cond139_out :
  _guard4976 ? idx_between_5_9_reg_out :
  1'd0;
assign cond143_write_en = _guard4977;
assign cond143_clk = clk;
assign cond143_reset = reset;
assign cond143_in =
  _guard4978 ? idx_between_6_10_reg_out :
  1'd0;
assign cond_wire143_in =
  _guard4979 ? idx_between_6_10_reg_out :
  _guard4982 ? cond143_out :
  1'd0;
assign cond148_write_en = _guard4983;
assign cond148_clk = clk;
assign cond148_reset = reset;
assign cond148_in =
  _guard4984 ? idx_between_7_15_reg_out :
  1'd0;
assign cond152_write_en = _guard4985;
assign cond152_clk = clk;
assign cond152_reset = reset;
assign cond152_in =
  _guard4986 ? idx_between_8_16_reg_out :
  1'd0;
assign cond_wire172_in =
  _guard4987 ? idx_between_6_10_reg_out :
  _guard4990 ? cond172_out :
  1'd0;
assign cond_wire178_in =
  _guard4991 ? idx_between_11_19_reg_out :
  _guard4994 ? cond178_out :
  1'd0;
assign cond_wire181_in =
  _guard4997 ? cond181_out :
  _guard4998 ? idx_between_8_16_reg_out :
  1'd0;
assign cond_wire189_in =
  _guard5001 ? cond189_out :
  _guard5002 ? idx_between_10_18_reg_out :
  1'd0;
assign cond192_write_en = _guard5003;
assign cond192_clk = clk;
assign cond192_reset = reset;
assign cond192_in =
  _guard5004 ? idx_between_11_15_reg_out :
  1'd0;
assign cond196_write_en = _guard5005;
assign cond196_clk = clk;
assign cond196_reset = reset;
assign cond196_in =
  _guard5006 ? idx_between_12_16_reg_out :
  1'd0;
assign cond203_write_en = _guard5007;
assign cond203_clk = clk;
assign cond203_reset = reset;
assign cond203_in =
  _guard5008 ? idx_between_25_26_reg_out :
  1'd0;
assign cond_wire203_in =
  _guard5009 ? idx_between_25_26_reg_out :
  _guard5012 ? cond203_out :
  1'd0;
assign cond208_write_en = _guard5013;
assign cond208_clk = clk;
assign cond208_reset = reset;
assign cond208_in =
  _guard5014 ? idx_between_19_20_reg_out :
  1'd0;
assign cond_wire210_in =
  _guard5015 ? idx_between_8_16_reg_out :
  _guard5018 ? cond210_out :
  1'd0;
assign cond_wire214_in =
  _guard5021 ? cond214_out :
  _guard5022 ? idx_between_9_17_reg_out :
  1'd0;
assign cond_wire233_in =
  _guard5025 ? cond233_out :
  _guard5026 ? idx_between_14_18_reg_out :
  1'd0;
assign cond235_write_en = _guard5027;
assign cond235_clk = clk;
assign cond235_reset = reset;
assign cond235_in =
  _guard5028 ? idx_between_18_26_reg_out :
  1'd0;
assign cond_wire248_in =
  _guard5031 ? cond248_out :
  _guard5032 ? idx_between_14_22_reg_out :
  1'd0;
assign cond250_write_en = _guard5033;
assign cond250_clk = clk;
assign cond250_reset = reset;
assign cond250_in =
  _guard5034 ? idx_between_11_15_reg_out :
  1'd0;
assign cond252_write_en = _guard5035;
assign cond252_clk = clk;
assign cond252_reset = reset;
assign cond252_in =
  _guard5036 ? idx_between_15_23_reg_out :
  1'd0;
assign cond_wire253_in =
  _guard5037 ? idx_between_23_24_reg_out :
  _guard5040 ? cond253_out :
  1'd0;
assign cond_wire256_in =
  _guard5043 ? cond256_out :
  _guard5044 ? idx_between_16_24_reg_out :
  1'd0;
assign cond_wire258_in =
  _guard5047 ? cond258_out :
  _guard5048 ? idx_between_13_17_reg_out :
  1'd0;
assign cond_wire268_in =
  _guard5049 ? idx_between_27_28_reg_out :
  _guard5052 ? cond268_out :
  1'd0;
assign adder0_left =
  _guard5053 ? fsm_out :
  1'd0;
assign adder0_right = _guard5054;
assign early_reset_static_seq_go_in = _guard5055;
assign top_0_2_write_en = _guard5058;
assign top_0_2_clk = clk;
assign top_0_2_reset = reset;
assign top_0_2_in = t2_read_data;
assign top_1_1_write_en = _guard5064;
assign top_1_1_clk = clk;
assign top_1_1_reset = reset;
assign top_1_1_in = top_0_1_out;
assign left_3_2_write_en = _guard5070;
assign left_3_2_clk = clk;
assign left_3_2_reset = reset;
assign left_3_2_in = left_3_1_out;
assign left_3_4_write_en = _guard5076;
assign left_3_4_clk = clk;
assign left_3_4_reset = reset;
assign left_3_4_in = left_3_3_out;
assign top_4_1_write_en = _guard5082;
assign top_4_1_clk = clk;
assign top_4_1_reset = reset;
assign top_4_1_in = top_3_1_out;
assign top_4_2_write_en = _guard5088;
assign top_4_2_clk = clk;
assign top_4_2_reset = reset;
assign top_4_2_in = top_3_2_out;
assign top_6_4_write_en = _guard5094;
assign top_6_4_clk = clk;
assign top_6_4_reset = reset;
assign top_6_4_in = top_5_4_out;
assign top_6_5_write_en = _guard5100;
assign top_6_5_clk = clk;
assign top_6_5_reset = reset;
assign top_6_5_in = top_5_5_out;
assign left_6_6_write_en = _guard5106;
assign left_6_6_clk = clk;
assign left_6_6_reset = reset;
assign left_6_6_in = left_6_5_out;
assign left_7_2_write_en = _guard5112;
assign left_7_2_clk = clk;
assign left_7_2_reset = reset;
assign left_7_2_in = left_7_1_out;
assign pe_7_5_mul_ready =
  _guard5118 ? 1'd1 :
  _guard5121 ? 1'd0 :
  1'd0;
assign pe_7_5_clk = clk;
assign pe_7_5_top =
  _guard5134 ? top_7_5_out :
  32'd0;
assign pe_7_5_left =
  _guard5147 ? left_7_5_out :
  32'd0;
assign pe_7_5_reset = reset;
assign pe_7_5_go = _guard5160;
assign pe_7_6_mul_ready =
  _guard5163 ? 1'd1 :
  _guard5166 ? 1'd0 :
  1'd0;
assign pe_7_6_clk = clk;
assign pe_7_6_top =
  _guard5179 ? top_7_6_out :
  32'd0;
assign pe_7_6_left =
  _guard5192 ? left_7_6_out :
  32'd0;
assign pe_7_6_reset = reset;
assign pe_7_6_go = _guard5205;
assign t0_add_left = 4'd1;
assign t0_add_right = t0_idx_out;
assign l0_add_left = 4'd1;
assign l0_add_right = l0_idx_out;
assign idx_between_5_13_comb_left = index_ge_5_out;
assign idx_between_5_13_comb_right = index_lt_13_out;
assign index_ge_9_left = idx_add_out;
assign index_ge_9_right = 5'd9;
assign idx_between_10_18_comb_left = index_ge_10_out;
assign idx_between_10_18_comb_right = index_lt_18_out;
assign idx_between_4_8_comb_left = index_ge_4_out;
assign idx_between_4_8_comb_right = index_lt_8_out;
assign index_ge_23_left = idx_add_out;
assign index_ge_23_right = 5'd23;
assign index_ge_11_left = idx_add_out;
assign index_ge_11_right = 5'd11;
assign index_lt_20_left = idx_add_out;
assign index_lt_20_right = 5'd20;
assign index_lt_21_left = idx_add_out;
assign index_lt_21_right = 5'd21;
assign idx_between_20_21_comb_left = index_ge_20_out;
assign idx_between_20_21_comb_right = index_lt_21_out;
assign idx_between_12_20_comb_left = index_ge_12_out;
assign idx_between_12_20_comb_right = index_lt_20_out;
assign idx_between_11_15_comb_left = index_ge_11_out;
assign idx_between_11_15_comb_right = index_lt_15_out;
assign idx_between_16_17_comb_left = index_ge_16_out;
assign idx_between_16_17_comb_right = index_lt_17_out;
assign cond_wire2_in =
  _guard5242 ? idx_between_5_13_reg_out :
  _guard5245 ? cond2_out :
  1'd0;
assign cond_wire9_in =
  _guard5248 ? cond9_out :
  _guard5249 ? idx_between_2_10_reg_out :
  1'd0;
assign cond10_write_en = _guard5250;
assign cond10_clk = clk;
assign cond10_reset = reset;
assign cond10_in =
  _guard5251 ? idx_between_3_7_reg_out :
  1'd0;
assign cond_wire11_in =
  _guard5254 ? cond11_out :
  _guard5255 ? idx_between_3_11_reg_out :
  1'd0;
assign cond21_write_en = _guard5256;
assign cond21_clk = clk;
assign cond21_reset = reset;
assign cond21_in =
  _guard5257 ? idx_between_5_13_reg_out :
  1'd0;
assign cond24_write_en = _guard5258;
assign cond24_clk = clk;
assign cond24_reset = reset;
assign cond24_in =
  _guard5259 ? idx_between_5_13_reg_out :
  1'd0;
assign cond31_write_en = _guard5260;
assign cond31_clk = clk;
assign cond31_reset = reset;
assign cond31_in =
  _guard5261 ? idx_between_7_15_reg_out :
  1'd0;
assign cond36_write_en = _guard5262;
assign cond36_clk = clk;
assign cond36_reset = reset;
assign cond36_in =
  _guard5263 ? idx_between_8_16_reg_out :
  1'd0;
assign cond_wire41_in =
  _guard5266 ? cond41_out :
  _guard5267 ? idx_between_2_10_reg_out :
  1'd0;
assign cond_wire45_in =
  _guard5270 ? cond45_out :
  _guard5271 ? idx_between_3_11_reg_out :
  1'd0;
assign cond51_write_en = _guard5272;
assign cond51_clk = clk;
assign cond51_reset = reset;
assign cond51_in =
  _guard5273 ? idx_between_16_17_reg_out :
  1'd0;
assign cond_wire57_in =
  _guard5274 ? idx_between_6_14_reg_out :
  _guard5277 ? cond57_out :
  1'd0;
assign cond_wire58_in =
  _guard5280 ? cond58_out :
  _guard5281 ? idx_between_10_18_reg_out :
  1'd0;
assign cond61_write_en = _guard5282;
assign cond61_clk = clk;
assign cond61_reset = reset;
assign cond61_in =
  _guard5283 ? idx_between_7_15_reg_out :
  1'd0;
assign cond80_write_en = _guard5284;
assign cond80_clk = clk;
assign cond80_reset = reset;
assign cond80_in =
  _guard5285 ? idx_between_16_17_reg_out :
  1'd0;
assign cond_wire80_in =
  _guard5286 ? idx_between_16_17_reg_out :
  _guard5289 ? cond80_out :
  1'd0;
assign cond86_write_en = _guard5290;
assign cond86_clk = clk;
assign cond86_reset = reset;
assign cond86_in =
  _guard5291 ? idx_between_6_14_reg_out :
  1'd0;
assign cond97_write_en = _guard5292;
assign cond97_clk = clk;
assign cond97_reset = reset;
assign cond97_in =
  _guard5293 ? idx_between_9_13_reg_out :
  1'd0;
assign cond_wire123_in =
  _guard5296 ? cond123_out :
  _guard5297 ? idx_between_8_16_reg_out :
  1'd0;
assign cond127_write_en = _guard5298;
assign cond127_clk = clk;
assign cond127_reset = reset;
assign cond127_in =
  _guard5299 ? idx_between_9_17_reg_out :
  1'd0;
assign cond129_write_en = _guard5300;
assign cond129_clk = clk;
assign cond129_reset = reset;
assign cond129_in =
  _guard5301 ? idx_between_21_22_reg_out :
  1'd0;
assign cond_wire129_in =
  _guard5302 ? idx_between_21_22_reg_out :
  _guard5305 ? cond129_out :
  1'd0;
assign cond_wire136_in =
  _guard5306 ? idx_between_15_23_reg_out :
  _guard5309 ? cond136_out :
  1'd0;
assign cond_wire145_in =
  _guard5310 ? idx_between_10_18_reg_out :
  _guard5313 ? cond145_out :
  1'd0;
assign cond170_write_en = _guard5314;
assign cond170_clk = clk;
assign cond170_reset = reset;
assign cond170_in =
  _guard5315 ? idx_between_24_25_reg_out :
  1'd0;
assign cond_wire184_in =
  _guard5318 ? cond184_out :
  _guard5319 ? idx_between_9_13_reg_out :
  1'd0;
assign cond_wire194_in =
  _guard5320 ? idx_between_15_23_reg_out :
  _guard5323 ? cond194_out :
  1'd0;
assign cond199_write_en = _guard5324;
assign cond199_clk = clk;
assign cond199_reset = reset;
assign cond199_in =
  _guard5325 ? idx_between_24_25_reg_out :
  1'd0;
assign cond_wire201_in =
  _guard5328 ? cond201_out :
  _guard5329 ? idx_between_13_21_reg_out :
  1'd0;
assign cond211_write_en = _guard5330;
assign cond211_clk = clk;
assign cond211_reset = reset;
assign cond211_in =
  _guard5331 ? idx_between_12_20_reg_out :
  1'd0;
assign cond_wire220_in =
  _guard5332 ? idx_between_22_23_reg_out :
  _guard5335 ? cond220_out :
  1'd0;
assign cond242_write_en = _guard5336;
assign cond242_clk = clk;
assign cond242_reset = reset;
assign cond242_in =
  _guard5337 ? idx_between_9_13_reg_out :
  1'd0;
assign cond_wire242_in =
  _guard5340 ? cond242_out :
  _guard5341 ? idx_between_9_13_reg_out :
  1'd0;
assign cond_wire246_in =
  _guard5342 ? idx_between_10_14_reg_out :
  _guard5345 ? cond246_out :
  1'd0;
assign cond249_write_en = _guard5346;
assign cond249_clk = clk;
assign cond249_reset = reset;
assign cond249_in =
  _guard5347 ? idx_between_22_23_reg_out :
  1'd0;
assign cond_wire249_in =
  _guard5348 ? idx_between_22_23_reg_out :
  _guard5351 ? cond249_out :
  1'd0;
assign cond_wire250_in =
  _guard5354 ? cond250_out :
  _guard5355 ? idx_between_11_15_reg_out :
  1'd0;
assign cond_wire251_in =
  _guard5356 ? idx_between_11_19_reg_out :
  _guard5359 ? cond251_out :
  1'd0;
assign cond268_write_en = _guard5360;
assign cond268_clk = clk;
assign cond268_reset = reset;
assign cond268_in =
  _guard5361 ? idx_between_27_28_reg_out :
  1'd0;
assign signal_reg_write_en = _guard5371;
assign signal_reg_clk = clk;
assign signal_reg_reset = reset;
assign signal_reg_in =
  _guard5377 ? 1'd1 :
  _guard5380 ? 1'd0 :
  1'd0;
assign top_0_4_write_en = _guard5383;
assign top_0_4_clk = clk;
assign top_0_4_reset = reset;
assign top_0_4_in = t4_read_data;
assign left_0_5_write_en = _guard5389;
assign left_0_5_clk = clk;
assign left_0_5_reset = reset;
assign left_0_5_in = left_0_4_out;
assign pe_2_0_mul_ready =
  _guard5395 ? 1'd1 :
  _guard5398 ? 1'd0 :
  1'd0;
assign pe_2_0_clk = clk;
assign pe_2_0_top =
  _guard5411 ? top_2_0_out :
  32'd0;
assign pe_2_0_left =
  _guard5424 ? left_2_0_out :
  32'd0;
assign pe_2_0_reset = reset;
assign pe_2_0_go = _guard5437;
assign left_2_1_write_en = _guard5440;
assign left_2_1_clk = clk;
assign left_2_1_reset = reset;
assign left_2_1_in = left_2_0_out;
assign top_2_2_write_en = _guard5446;
assign top_2_2_clk = clk;
assign top_2_2_reset = reset;
assign top_2_2_in = top_1_2_out;
assign left_2_5_write_en = _guard5452;
assign left_2_5_clk = clk;
assign left_2_5_reset = reset;
assign left_2_5_in = left_2_4_out;
assign left_3_6_write_en = _guard5458;
assign left_3_6_clk = clk;
assign left_3_6_reset = reset;
assign left_3_6_in = left_3_5_out;
assign pe_4_4_mul_ready =
  _guard5464 ? 1'd1 :
  _guard5467 ? 1'd0 :
  1'd0;
assign pe_4_4_clk = clk;
assign pe_4_4_top =
  _guard5480 ? top_4_4_out :
  32'd0;
assign pe_4_4_left =
  _guard5493 ? left_4_4_out :
  32'd0;
assign pe_4_4_reset = reset;
assign pe_4_4_go = _guard5506;
assign left_4_4_write_en = _guard5509;
assign left_4_4_clk = clk;
assign left_4_4_reset = reset;
assign left_4_4_in = left_4_3_out;
assign pe_4_7_mul_ready =
  _guard5515 ? 1'd1 :
  _guard5518 ? 1'd0 :
  1'd0;
assign pe_4_7_clk = clk;
assign pe_4_7_top =
  _guard5531 ? top_4_7_out :
  32'd0;
assign pe_4_7_left =
  _guard5544 ? left_4_7_out :
  32'd0;
assign pe_4_7_reset = reset;
assign pe_4_7_go = _guard5557;
assign left_5_5_write_en = _guard5560;
assign left_5_5_clk = clk;
assign left_5_5_reset = reset;
assign left_5_5_in = left_5_4_out;
assign left_7_0_write_en = _guard5566;
assign left_7_0_clk = clk;
assign left_7_0_reset = reset;
assign left_7_0_in = l7_read_data;
assign top_7_3_write_en = _guard5572;
assign top_7_3_clk = clk;
assign top_7_3_reset = reset;
assign top_7_3_in = top_6_3_out;
assign top_7_6_write_en = _guard5578;
assign top_7_6_clk = clk;
assign top_7_6_reset = reset;
assign top_7_6_in = top_6_6_out;
assign t1_add_left = 4'd1;
assign t1_add_right = t1_idx_out;
assign t3_idx_write_en = _guard5594;
assign t3_idx_clk = clk;
assign t3_idx_reset = reset;
assign t3_idx_in =
  _guard5597 ? t3_add_out :
  _guard5600 ? 4'd0 :
  'x;
assign l4_add_left = 4'd1;
assign l4_add_right = l4_idx_out;
assign idx_between_12_16_reg_write_en = _guard5611;
assign idx_between_12_16_reg_clk = clk;
assign idx_between_12_16_reg_reset = reset;
assign idx_between_12_16_reg_in =
  _guard5612 ? idx_between_12_16_comb_out :
  _guard5615 ? 1'd0 :
  'x;
assign index_lt_22_left = idx_add_out;
assign index_lt_22_right = 5'd22;
assign index_ge_22_left = idx_add_out;
assign index_ge_22_right = 5'd22;
assign idx_between_22_23_comb_left = index_ge_22_out;
assign idx_between_22_23_comb_right = index_lt_23_out;
assign index_ge_19_left = idx_add_out;
assign index_ge_19_right = 5'd19;
assign idx_between_19_27_comb_left = index_ge_19_out;
assign idx_between_19_27_comb_right = index_lt_27_out;
assign idx_between_13_17_reg_write_en = _guard5630;
assign idx_between_13_17_reg_clk = clk;
assign idx_between_13_17_reg_reset = reset;
assign idx_between_13_17_reg_in =
  _guard5631 ? idx_between_13_17_comb_out :
  _guard5634 ? 1'd0 :
  'x;
assign idx_between_18_19_comb_left = index_ge_18_out;
assign idx_between_18_19_comb_right = index_lt_19_out;
assign idx_between_2_10_reg_write_en = _guard5641;
assign idx_between_2_10_reg_clk = clk;
assign idx_between_2_10_reg_reset = reset;
assign idx_between_2_10_reg_in =
  _guard5642 ? idx_between_2_10_comb_out :
  _guard5645 ? 1'd0 :
  'x;
assign index_lt_10_left = idx_add_out;
assign index_lt_10_right = 5'd10;
assign index_ge_2_left = idx_add_out;
assign index_ge_2_right = 5'd2;
assign index_ge_16_left = idx_add_out;
assign index_ge_16_right = 5'd16;
assign cond_wire_in =
  _guard5654 ? cond_out :
  _guard5655 ? idx_between_0_8_reg_out :
  1'd0;
assign cond_wire15_in =
  _guard5658 ? cond15_out :
  _guard5659 ? idx_between_4_8_reg_out :
  1'd0;
assign cond16_write_en = _guard5660;
assign cond16_clk = clk;
assign cond16_reset = reset;
assign cond16_in =
  _guard5661 ? idx_between_4_12_reg_out :
  1'd0;
assign cond37_write_en = _guard5662;
assign cond37_clk = clk;
assign cond37_reset = reset;
assign cond37_in =
  _guard5663 ? idx_between_12_20_reg_out :
  1'd0;
assign cond_wire49_in =
  _guard5664 ? idx_between_4_12_reg_out :
  _guard5667 ? cond49_out :
  1'd0;
assign cond_wire55_in =
  _guard5668 ? idx_between_17_18_reg_out :
  _guard5671 ? cond55_out :
  1'd0;
assign cond_wire93_in =
  _guard5672 ? idx_between_8_12_reg_out :
  _guard5675 ? cond93_out :
  1'd0;
assign cond_wire95_in =
  _guard5678 ? cond95_out :
  _guard5679 ? idx_between_12_20_reg_out :
  1'd0;
assign cond_wire96_in =
  _guard5680 ? idx_between_20_21_reg_out :
  _guard5683 ? cond96_out :
  1'd0;
assign cond_wire99_in =
  _guard5684 ? idx_between_13_21_reg_out :
  _guard5687 ? cond99_out :
  1'd0;
assign cond110_write_en = _guard5688;
assign cond110_clk = clk;
assign cond110_reset = reset;
assign cond110_in =
  _guard5689 ? idx_between_5_9_reg_out :
  1'd0;
assign cond113_write_en = _guard5690;
assign cond113_clk = clk;
assign cond113_reset = reset;
assign cond113_in =
  _guard5691 ? idx_between_17_18_reg_out :
  1'd0;
assign cond_wire113_in =
  _guard5692 ? idx_between_17_18_reg_out :
  _guard5695 ? cond113_out :
  1'd0;
assign cond_wire114_in =
  _guard5696 ? idx_between_6_10_reg_out :
  _guard5699 ? cond114_out :
  1'd0;
assign cond125_write_en = _guard5700;
assign cond125_clk = clk;
assign cond125_reset = reset;
assign cond125_in =
  _guard5701 ? idx_between_20_21_reg_out :
  1'd0;
assign cond130_write_en = _guard5702;
assign cond130_clk = clk;
assign cond130_reset = reset;
assign cond130_in =
  _guard5703 ? idx_between_10_14_reg_out :
  1'd0;
assign cond_wire133_in =
  _guard5704 ? idx_between_22_23_reg_out :
  _guard5707 ? cond133_out :
  1'd0;
assign cond144_write_en = _guard5708;
assign cond144_clk = clk;
assign cond144_reset = reset;
assign cond144_in =
  _guard5709 ? idx_between_6_14_reg_out :
  1'd0;
assign cond_wire155_in =
  _guard5712 ? cond155_out :
  _guard5713 ? idx_between_9_13_reg_out :
  1'd0;
assign cond160_write_en = _guard5714;
assign cond160_clk = clk;
assign cond160_reset = reset;
assign cond160_in =
  _guard5715 ? idx_between_10_18_reg_out :
  1'd0;
assign cond163_write_en = _guard5716;
assign cond163_clk = clk;
assign cond163_reset = reset;
assign cond163_in =
  _guard5717 ? idx_between_11_15_reg_out :
  1'd0;
assign cond165_write_en = _guard5718;
assign cond165_clk = clk;
assign cond165_reset = reset;
assign cond165_in =
  _guard5719 ? idx_between_15_23_reg_out :
  1'd0;
assign cond168_write_en = _guard5720;
assign cond168_clk = clk;
assign cond168_reset = reset;
assign cond168_in =
  _guard5721 ? idx_between_12_20_reg_out :
  1'd0;
assign cond_wire173_in =
  _guard5722 ? idx_between_6_14_reg_out :
  _guard5725 ? cond173_out :
  1'd0;
assign cond_wire179_in =
  _guard5728 ? cond179_out :
  _guard5729 ? idx_between_19_20_reg_out :
  1'd0;
assign cond184_write_en = _guard5730;
assign cond184_clk = clk;
assign cond184_reset = reset;
assign cond184_in =
  _guard5731 ? idx_between_9_13_reg_out :
  1'd0;
assign cond185_write_en = _guard5732;
assign cond185_clk = clk;
assign cond185_reset = reset;
assign cond185_in =
  _guard5733 ? idx_between_9_17_reg_out :
  1'd0;
assign cond195_write_en = _guard5734;
assign cond195_clk = clk;
assign cond195_reset = reset;
assign cond195_in =
  _guard5735 ? idx_between_23_24_reg_out :
  1'd0;
assign cond197_write_en = _guard5736;
assign cond197_clk = clk;
assign cond197_reset = reset;
assign cond197_in =
  _guard5737 ? idx_between_12_20_reg_out :
  1'd0;
assign cond207_write_en = _guard5738;
assign cond207_clk = clk;
assign cond207_reset = reset;
assign cond207_in =
  _guard5739 ? idx_between_11_19_reg_out :
  1'd0;
assign cond_wire217_in =
  _guard5742 ? cond217_out :
  _guard5743 ? idx_between_10_14_reg_out :
  1'd0;
assign cond_wire219_in =
  _guard5746 ? cond219_out :
  _guard5747 ? idx_between_14_22_reg_out :
  1'd0;
assign cond_wire241_in =
  _guard5748 ? idx_between_20_21_reg_out :
  _guard5751 ? cond241_out :
  1'd0;
assign cond243_write_en = _guard5752;
assign cond243_clk = clk;
assign cond243_reset = reset;
assign cond243_in =
  _guard5753 ? idx_between_9_17_reg_out :
  1'd0;
assign cond_wire244_in =
  _guard5756 ? cond244_out :
  _guard5757 ? idx_between_13_21_reg_out :
  1'd0;
assign cond267_write_en = _guard5758;
assign cond267_clk = clk;
assign cond267_reset = reset;
assign cond267_in =
  _guard5759 ? idx_between_19_27_reg_out :
  1'd0;
assign pe_0_0_mul_ready =
  _guard5762 ? 1'd1 :
  _guard5765 ? 1'd0 :
  1'd0;
assign pe_0_0_clk = clk;
assign pe_0_0_top =
  _guard5778 ? top_0_0_out :
  32'd0;
assign pe_0_0_left =
  _guard5791 ? left_0_0_out :
  32'd0;
assign pe_0_0_reset = reset;
assign pe_0_0_go = _guard5804;
assign left_1_6_write_en = _guard5807;
assign left_1_6_clk = clk;
assign left_1_6_reset = reset;
assign left_1_6_in = left_1_5_out;
assign pe_3_3_mul_ready =
  _guard5813 ? 1'd1 :
  _guard5816 ? 1'd0 :
  1'd0;
assign pe_3_3_clk = clk;
assign pe_3_3_top =
  _guard5829 ? top_3_3_out :
  32'd0;
assign pe_3_3_left =
  _guard5842 ? left_3_3_out :
  32'd0;
assign pe_3_3_reset = reset;
assign pe_3_3_go = _guard5855;
assign top_3_3_write_en = _guard5858;
assign top_3_3_clk = clk;
assign top_3_3_reset = reset;
assign top_3_3_in = top_2_3_out;
assign top_4_3_write_en = _guard5864;
assign top_4_3_clk = clk;
assign top_4_3_reset = reset;
assign top_4_3_in = top_3_3_out;
assign top_4_6_write_en = _guard5870;
assign top_4_6_clk = clk;
assign top_4_6_reset = reset;
assign top_4_6_in = top_3_6_out;
assign pe_5_6_mul_ready =
  _guard5876 ? 1'd1 :
  _guard5879 ? 1'd0 :
  1'd0;
assign pe_5_6_clk = clk;
assign pe_5_6_top =
  _guard5892 ? top_5_6_out :
  32'd0;
assign pe_5_6_left =
  _guard5905 ? left_5_6_out :
  32'd0;
assign pe_5_6_reset = reset;
assign pe_5_6_go = _guard5918;
assign top_5_6_write_en = _guard5921;
assign top_5_6_clk = clk;
assign top_5_6_reset = reset;
assign top_5_6_in = top_4_6_out;
assign top_6_2_write_en = _guard5927;
assign top_6_2_clk = clk;
assign top_6_2_reset = reset;
assign top_6_2_in = top_5_2_out;
assign pe_7_1_mul_ready =
  _guard5933 ? 1'd1 :
  _guard5936 ? 1'd0 :
  1'd0;
assign pe_7_1_clk = clk;
assign pe_7_1_top =
  _guard5949 ? top_7_1_out :
  32'd0;
assign pe_7_1_left =
  _guard5962 ? left_7_1_out :
  32'd0;
assign pe_7_1_reset = reset;
assign pe_7_1_go = _guard5975;
assign t2_add_left = 4'd1;
assign t2_add_right = t2_idx_out;
assign t5_add_left = 4'd1;
assign t5_add_right = t5_idx_out;
assign index_lt_12_left = idx_add_out;
assign index_lt_12_right = 5'd12;
assign index_ge_5_left = idx_add_out;
assign index_ge_5_right = 5'd5;
assign index_ge_10_left = idx_add_out;
assign index_ge_10_right = 5'd10;
assign idx_between_27_28_comb_left = index_ge_27_out;
assign idx_between_27_28_comb_right = index_lt_28_out;
assign idx_between_7_11_comb_left = index_ge_7_out;
assign idx_between_7_11_comb_right = index_lt_11_out;
assign idx_between_17_25_reg_write_en = _guard6002;
assign idx_between_17_25_reg_clk = clk;
assign idx_between_17_25_reg_reset = reset;
assign idx_between_17_25_reg_in =
  _guard6003 ? idx_between_17_25_comb_out :
  _guard6006 ? 1'd0 :
  'x;
assign cond0_write_en = _guard6007;
assign cond0_clk = clk;
assign cond0_reset = reset;
assign cond0_in =
  _guard6008 ? idx_between_1_5_reg_out :
  1'd0;
assign cond_wire7_in =
  _guard6009 ? idx_between_6_14_reg_out :
  _guard6012 ? cond7_out :
  1'd0;
assign cond_wire10_in =
  _guard6013 ? idx_between_3_7_reg_out :
  _guard6016 ? cond10_out :
  1'd0;
assign cond_wire12_in =
  _guard6017 ? idx_between_7_15_reg_out :
  _guard6020 ? cond12_out :
  1'd0;
assign cond_wire17_in =
  _guard6023 ? cond17_out :
  _guard6024 ? idx_between_8_16_reg_out :
  1'd0;
assign cond_wire19_in =
  _guard6027 ? cond19_out :
  _guard6028 ? idx_between_4_12_reg_out :
  1'd0;
assign cond_wire23_in =
  _guard6029 ? idx_between_17_18_reg_out :
  _guard6032 ? cond23_out :
  1'd0;
assign cond_wire25_in =
  _guard6033 ? idx_between_6_10_reg_out :
  _guard6036 ? cond25_out :
  1'd0;
assign cond33_write_en = _guard6037;
assign cond33_clk = clk;
assign cond33_reset = reset;
assign cond33_in =
  _guard6038 ? idx_between_19_20_reg_out :
  1'd0;
assign cond_wire42_in =
  _guard6039 ? idx_between_6_14_reg_out :
  _guard6042 ? cond42_out :
  1'd0;
assign cond47_write_en = _guard6043;
assign cond47_clk = clk;
assign cond47_reset = reset;
assign cond47_in =
  _guard6044 ? idx_between_15_16_reg_out :
  1'd0;
assign cond48_write_en = _guard6045;
assign cond48_clk = clk;
assign cond48_reset = reset;
assign cond48_in =
  _guard6046 ? idx_between_4_8_reg_out :
  1'd0;
assign cond66_write_en = _guard6047;
assign cond66_clk = clk;
assign cond66_reset = reset;
assign cond66_in =
  _guard6048 ? idx_between_12_20_reg_out :
  1'd0;
assign cond_wire69_in =
  _guard6051 ? cond69_out :
  _guard6052 ? idx_between_9_17_reg_out :
  1'd0;
assign cond_wire71_in =
  _guard6055 ? cond71_out :
  _guard6056 ? idx_between_21_22_reg_out :
  1'd0;
assign cond82_write_en = _guard6057;
assign cond82_clk = clk;
assign cond82_reset = reset;
assign cond82_in =
  _guard6058 ? idx_between_5_13_reg_out :
  1'd0;
assign cond84_write_en = _guard6059;
assign cond84_clk = clk;
assign cond84_reset = reset;
assign cond84_in =
  _guard6060 ? idx_between_17_18_reg_out :
  1'd0;
assign cond_wire94_in =
  _guard6063 ? cond94_out :
  _guard6064 ? idx_between_8_16_reg_out :
  1'd0;
assign cond102_write_en = _guard6065;
assign cond102_clk = clk;
assign cond102_reset = reset;
assign cond102_in =
  _guard6066 ? idx_between_10_18_reg_out :
  1'd0;
assign cond_wire104_in =
  _guard6067 ? idx_between_22_23_reg_out :
  _guard6070 ? cond104_out :
  1'd0;
assign cond108_write_en = _guard6071;
assign cond108_clk = clk;
assign cond108_reset = reset;
assign cond108_in =
  _guard6072 ? idx_between_8_16_reg_out :
  1'd0;
assign cond_wire110_in =
  _guard6073 ? idx_between_5_9_reg_out :
  _guard6076 ? cond110_out :
  1'd0;
assign cond119_write_en = _guard6077;
assign cond119_clk = clk;
assign cond119_reset = reset;
assign cond119_in =
  _guard6078 ? idx_between_7_15_reg_out :
  1'd0;
assign cond120_write_en = _guard6079;
assign cond120_clk = clk;
assign cond120_reset = reset;
assign cond120_in =
  _guard6080 ? idx_between_11_19_reg_out :
  1'd0;
assign cond_wire130_in =
  _guard6083 ? cond130_out :
  _guard6084 ? idx_between_10_14_reg_out :
  1'd0;
assign cond_wire135_in =
  _guard6085 ? idx_between_11_19_reg_out :
  _guard6088 ? cond135_out :
  1'd0;
assign cond141_write_en = _guard6089;
assign cond141_clk = clk;
assign cond141_reset = reset;
assign cond141_in =
  _guard6090 ? idx_between_9_17_reg_out :
  1'd0;
assign cond_wire150_in =
  _guard6093 ? cond150_out :
  _guard6094 ? idx_between_19_20_reg_out :
  1'd0;
assign cond_wire152_in =
  _guard6095 ? idx_between_8_16_reg_out :
  _guard6098 ? cond152_out :
  1'd0;
assign cond_wire153_in =
  _guard6099 ? idx_between_12_20_reg_out :
  _guard6102 ? cond153_out :
  1'd0;
assign cond210_write_en = _guard6103;
assign cond210_clk = clk;
assign cond210_reset = reset;
assign cond210_in =
  _guard6104 ? idx_between_8_16_reg_out :
  1'd0;
assign cond218_write_en = _guard6105;
assign cond218_clk = clk;
assign cond218_reset = reset;
assign cond218_in =
  _guard6106 ? idx_between_10_18_reg_out :
  1'd0;
assign cond229_write_en = _guard6107;
assign cond229_clk = clk;
assign cond229_reset = reset;
assign cond229_in =
  _guard6108 ? idx_between_13_17_reg_out :
  1'd0;
assign cond_wire255_in =
  _guard6111 ? cond255_out :
  _guard6112 ? idx_between_12_20_reg_out :
  1'd0;
assign cond_wire266_in =
  _guard6113 ? idx_between_15_19_reg_out :
  _guard6116 ? cond266_out :
  1'd0;
assign early_reset_static_seq_done_in = ud_out;
assign top_0_3_write_en = _guard6119;
assign top_0_3_clk = clk;
assign top_0_3_reset = reset;
assign top_0_3_in = t3_read_data;
assign pe_0_6_mul_ready =
  _guard6125 ? 1'd1 :
  _guard6128 ? 1'd0 :
  1'd0;
assign pe_0_6_clk = clk;
assign pe_0_6_top =
  _guard6141 ? top_0_6_out :
  32'd0;
assign pe_0_6_left =
  _guard6154 ? left_0_6_out :
  32'd0;
assign pe_0_6_reset = reset;
assign pe_0_6_go = _guard6167;
assign top_1_7_write_en = _guard6170;
assign top_1_7_clk = clk;
assign top_1_7_reset = reset;
assign top_1_7_in = top_0_7_out;
assign top_2_1_write_en = _guard6176;
assign top_2_1_clk = clk;
assign top_2_1_reset = reset;
assign top_2_1_in = top_1_1_out;
assign left_3_3_write_en = _guard6182;
assign left_3_3_clk = clk;
assign left_3_3_reset = reset;
assign left_3_3_in = left_3_2_out;
assign top_3_7_write_en = _guard6188;
assign top_3_7_clk = clk;
assign top_3_7_reset = reset;
assign top_3_7_in = top_2_7_out;
assign left_4_1_write_en = _guard6194;
assign left_4_1_clk = clk;
assign left_4_1_reset = reset;
assign left_4_1_in = left_4_0_out;
assign pe_4_3_mul_ready =
  _guard6200 ? 1'd1 :
  _guard6203 ? 1'd0 :
  1'd0;
assign pe_4_3_clk = clk;
assign pe_4_3_top =
  _guard6216 ? top_4_3_out :
  32'd0;
assign pe_4_3_left =
  _guard6229 ? left_4_3_out :
  32'd0;
assign pe_4_3_reset = reset;
assign pe_4_3_go = _guard6242;
assign left_5_0_write_en = _guard6245;
assign left_5_0_clk = clk;
assign left_5_0_reset = reset;
assign left_5_0_in = l5_read_data;
assign pe_6_6_mul_ready =
  _guard6251 ? 1'd1 :
  _guard6254 ? 1'd0 :
  1'd0;
assign pe_6_6_clk = clk;
assign pe_6_6_top =
  _guard6267 ? top_6_6_out :
  32'd0;
assign pe_6_6_left =
  _guard6280 ? left_6_6_out :
  32'd0;
assign pe_6_6_reset = reset;
assign pe_6_6_go = _guard6293;
assign pe_7_2_mul_ready =
  _guard6296 ? 1'd1 :
  _guard6299 ? 1'd0 :
  1'd0;
assign pe_7_2_clk = clk;
assign pe_7_2_top =
  _guard6312 ? top_7_2_out :
  32'd0;
assign pe_7_2_left =
  _guard6325 ? left_7_2_out :
  32'd0;
assign pe_7_2_reset = reset;
assign pe_7_2_go = _guard6338;
assign pe_7_7_mul_ready =
  _guard6341 ? 1'd1 :
  _guard6344 ? 1'd0 :
  1'd0;
assign pe_7_7_clk = clk;
assign pe_7_7_top =
  _guard6357 ? top_7_7_out :
  32'd0;
assign pe_7_7_left =
  _guard6370 ? left_7_7_out :
  32'd0;
assign pe_7_7_reset = reset;
assign pe_7_7_go = _guard6383;
assign t2_idx_write_en = _guard6390;
assign t2_idx_clk = clk;
assign t2_idx_reset = reset;
assign t2_idx_in =
  _guard6393 ? 4'd0 :
  _guard6396 ? t2_add_out :
  'x;
assign l2_idx_write_en = _guard6403;
assign l2_idx_clk = clk;
assign l2_idx_reset = reset;
assign l2_idx_in =
  _guard6406 ? 4'd0 :
  _guard6409 ? l2_add_out :
  'x;
assign l6_idx_write_en = _guard6416;
assign l6_idx_clk = clk;
assign l6_idx_reset = reset;
assign l6_idx_in =
  _guard6419 ? 4'd0 :
  _guard6422 ? l6_add_out :
  'x;
assign index_lt_7_left = idx_add_out;
assign index_lt_7_right = 5'd7;
assign index_ge_26_left = idx_add_out;
assign index_ge_26_right = 5'd26;
assign idx_between_14_22_reg_write_en = _guard6431;
assign idx_between_14_22_reg_clk = clk;
assign idx_between_14_22_reg_reset = reset;
assign idx_between_14_22_reg_in =
  _guard6432 ? idx_between_14_22_comb_out :
  _guard6435 ? 1'd0 :
  'x;
assign idx_between_25_26_comb_left = index_ge_25_out;
assign idx_between_25_26_comb_right = index_lt_26_out;
assign index_ge_27_left = idx_add_out;
assign index_ge_27_right = 5'd27;
assign index_ge_6_left = idx_add_out;
assign index_ge_6_right = 5'd6;
assign idx_between_18_19_reg_write_en = _guard6446;
assign idx_between_18_19_reg_clk = clk;
assign idx_between_18_19_reg_reset = reset;
assign idx_between_18_19_reg_in =
  _guard6449 ? 1'd0 :
  _guard6450 ? idx_between_18_19_comb_out :
  'x;
assign idx_between_11_19_comb_left = index_ge_11_out;
assign idx_between_11_19_comb_right = index_lt_19_out;
assign idx_between_19_20_comb_left = index_ge_19_out;
assign idx_between_19_20_comb_right = index_lt_20_out;
assign idx_between_12_20_reg_write_en = _guard6459;
assign idx_between_12_20_reg_clk = clk;
assign idx_between_12_20_reg_reset = reset;
assign idx_between_12_20_reg_in =
  _guard6462 ? 1'd0 :
  _guard6463 ? idx_between_12_20_comb_out :
  'x;
assign idx_between_13_21_reg_write_en = _guard6468;
assign idx_between_13_21_reg_clk = clk;
assign idx_between_13_21_reg_reset = reset;
assign idx_between_13_21_reg_in =
  _guard6469 ? idx_between_13_21_comb_out :
  _guard6472 ? 1'd0 :
  'x;
assign cond1_write_en = _guard6473;
assign cond1_clk = clk;
assign cond1_reset = reset;
assign cond1_in =
  _guard6474 ? idx_between_1_9_reg_out :
  1'd0;
assign cond2_write_en = _guard6475;
assign cond2_clk = clk;
assign cond2_reset = reset;
assign cond2_in =
  _guard6476 ? idx_between_5_13_reg_out :
  1'd0;
assign cond_wire5_in =
  _guard6479 ? cond5_out :
  _guard6480 ? idx_between_2_6_reg_out :
  1'd0;
assign cond22_write_en = _guard6481;
assign cond22_clk = clk;
assign cond22_reset = reset;
assign cond22_in =
  _guard6482 ? idx_between_9_17_reg_out :
  1'd0;
assign cond26_write_en = _guard6483;
assign cond26_clk = clk;
assign cond26_reset = reset;
assign cond26_in =
  _guard6484 ? idx_between_6_14_reg_out :
  1'd0;
assign cond_wire34_in =
  _guard6485 ? idx_between_7_15_reg_out :
  _guard6488 ? cond34_out :
  1'd0;
assign cond39_write_en = _guard6489;
assign cond39_clk = clk;
assign cond39_reset = reset;
assign cond39_in =
  _guard6490 ? idx_between_1_9_reg_out :
  1'd0;
assign cond49_write_en = _guard6491;
assign cond49_clk = clk;
assign cond49_reset = reset;
assign cond49_in =
  _guard6492 ? idx_between_4_12_reg_out :
  1'd0;
assign cond_wire52_in =
  _guard6495 ? cond52_out :
  _guard6496 ? idx_between_5_9_reg_out :
  1'd0;
assign cond_wire68_in =
  _guard6499 ? cond68_out :
  _guard6500 ? idx_between_9_13_reg_out :
  1'd0;
assign cond_wire70_in =
  _guard6503 ? cond70_out :
  _guard6504 ? idx_between_13_21_reg_out :
  1'd0;
assign cond_wire83_in =
  _guard6507 ? cond83_out :
  _guard6508 ? idx_between_9_17_reg_out :
  1'd0;
assign cond87_write_en = _guard6509;
assign cond87_clk = clk;
assign cond87_reset = reset;
assign cond87_in =
  _guard6510 ? idx_between_10_18_reg_out :
  1'd0;
assign cond96_write_en = _guard6511;
assign cond96_clk = clk;
assign cond96_reset = reset;
assign cond96_in =
  _guard6512 ? idx_between_20_21_reg_out :
  1'd0;
assign cond_wire97_in =
  _guard6515 ? cond97_out :
  _guard6516 ? idx_between_9_13_reg_out :
  1'd0;
assign cond99_write_en = _guard6517;
assign cond99_clk = clk;
assign cond99_reset = reset;
assign cond99_in =
  _guard6518 ? idx_between_13_21_reg_out :
  1'd0;
assign cond104_write_en = _guard6519;
assign cond104_clk = clk;
assign cond104_reset = reset;
assign cond104_in =
  _guard6520 ? idx_between_22_23_reg_out :
  1'd0;
assign cond133_write_en = _guard6521;
assign cond133_clk = clk;
assign cond133_reset = reset;
assign cond133_in =
  _guard6522 ? idx_between_22_23_reg_out :
  1'd0;
assign cond138_write_en = _guard6523;
assign cond138_clk = clk;
assign cond138_reset = reset;
assign cond138_in =
  _guard6524 ? idx_between_4_12_reg_out :
  1'd0;
assign cond145_write_en = _guard6525;
assign cond145_clk = clk;
assign cond145_reset = reset;
assign cond145_in =
  _guard6526 ? idx_between_10_18_reg_out :
  1'd0;
assign cond147_write_en = _guard6527;
assign cond147_clk = clk;
assign cond147_reset = reset;
assign cond147_in =
  _guard6528 ? idx_between_7_11_reg_out :
  1'd0;
assign cond_wire147_in =
  _guard6529 ? idx_between_7_11_reg_out :
  _guard6532 ? cond147_out :
  1'd0;
assign cond154_write_en = _guard6533;
assign cond154_clk = clk;
assign cond154_reset = reset;
assign cond154_in =
  _guard6534 ? idx_between_20_21_reg_out :
  1'd0;
assign cond156_write_en = _guard6535;
assign cond156_clk = clk;
assign cond156_reset = reset;
assign cond156_in =
  _guard6536 ? idx_between_9_17_reg_out :
  1'd0;
assign cond_wire168_in =
  _guard6539 ? cond168_out :
  _guard6540 ? idx_between_12_20_reg_out :
  1'd0;
assign cond173_write_en = _guard6541;
assign cond173_clk = clk;
assign cond173_reset = reset;
assign cond173_in =
  _guard6542 ? idx_between_6_14_reg_out :
  1'd0;
assign cond175_write_en = _guard6543;
assign cond175_clk = clk;
assign cond175_reset = reset;
assign cond175_in =
  _guard6544 ? idx_between_18_19_reg_out :
  1'd0;
assign cond182_write_en = _guard6545;
assign cond182_clk = clk;
assign cond182_reset = reset;
assign cond182_in =
  _guard6546 ? idx_between_12_20_reg_out :
  1'd0;
assign cond_wire199_in =
  _guard6547 ? idx_between_24_25_reg_out :
  _guard6550 ? cond199_out :
  1'd0;
assign cond_wire206_in =
  _guard6553 ? cond206_out :
  _guard6554 ? idx_between_7_15_reg_out :
  1'd0;
assign cond212_write_en = _guard6555;
assign cond212_clk = clk;
assign cond212_reset = reset;
assign cond212_in =
  _guard6556 ? idx_between_20_21_reg_out :
  1'd0;
assign cond_wire212_in =
  _guard6557 ? idx_between_20_21_reg_out :
  _guard6560 ? cond212_out :
  1'd0;
assign cond224_write_en = _guard6561;
assign cond224_clk = clk;
assign cond224_reset = reset;
assign cond224_in =
  _guard6562 ? idx_between_23_24_reg_out :
  1'd0;
assign cond_wire229_in =
  _guard6563 ? idx_between_13_17_reg_out :
  _guard6566 ? cond229_out :
  1'd0;
assign cond_wire232_in =
  _guard6567 ? idx_between_25_26_reg_out :
  _guard6570 ? cond232_out :
  1'd0;
assign cond_wire247_in =
  _guard6573 ? cond247_out :
  _guard6574 ? idx_between_10_18_reg_out :
  1'd0;
assign cond259_write_en = _guard6575;
assign cond259_clk = clk;
assign cond259_reset = reset;
assign cond259_in =
  _guard6576 ? idx_between_13_21_reg_out :
  1'd0;
assign cond_wire259_in =
  _guard6577 ? idx_between_13_21_reg_out :
  _guard6580 ? cond259_out :
  1'd0;
assign cond260_write_en = _guard6581;
assign cond260_clk = clk;
assign cond260_reset = reset;
assign cond260_in =
  _guard6582 ? idx_between_17_25_reg_out :
  1'd0;
assign top_0_0_write_en = _guard6585;
assign top_0_0_clk = clk;
assign top_0_0_reset = reset;
assign top_0_0_in = t0_read_data;
assign top_0_5_write_en = _guard6591;
assign top_0_5_clk = clk;
assign top_0_5_reset = reset;
assign top_0_5_in = t5_read_data;
assign pe_1_1_mul_ready =
  _guard6597 ? 1'd1 :
  _guard6600 ? 1'd0 :
  1'd0;
assign pe_1_1_clk = clk;
assign pe_1_1_top =
  _guard6613 ? top_1_1_out :
  32'd0;
assign pe_1_1_left =
  _guard6626 ? left_1_1_out :
  32'd0;
assign pe_1_1_reset = reset;
assign pe_1_1_go = _guard6639;
assign top_2_7_write_en = _guard6642;
assign top_2_7_clk = clk;
assign top_2_7_reset = reset;
assign top_2_7_in = top_1_7_out;
assign left_5_2_write_en = _guard6648;
assign left_5_2_clk = clk;
assign left_5_2_reset = reset;
assign left_5_2_in = left_5_1_out;
assign top_5_7_write_en = _guard6654;
assign top_5_7_clk = clk;
assign top_5_7_reset = reset;
assign top_5_7_in = top_4_7_out;
assign left_5_7_write_en = _guard6660;
assign left_5_7_clk = clk;
assign left_5_7_reset = reset;
assign left_5_7_in = left_5_6_out;
assign left_6_0_write_en = _guard6666;
assign left_6_0_clk = clk;
assign left_6_0_reset = reset;
assign left_6_0_in = l6_read_data;
assign top_7_1_write_en = _guard6672;
assign top_7_1_clk = clk;
assign top_7_1_reset = reset;
assign top_7_1_in = top_6_1_out;
assign idx_between_8_12_comb_left = index_ge_8_out;
assign idx_between_8_12_comb_right = index_lt_12_out;
assign idx_between_9_17_reg_write_en = _guard6682;
assign idx_between_9_17_reg_clk = clk;
assign idx_between_9_17_reg_reset = reset;
assign idx_between_9_17_reg_in =
  _guard6683 ? idx_between_9_17_comb_out :
  _guard6686 ? 1'd0 :
  'x;
assign index_lt_18_left = idx_add_out;
assign index_lt_18_right = 5'd18;
assign index_lt_28_left = idx_add_out;
assign index_lt_28_right = 5'd28;
assign index_ge_13_left = idx_add_out;
assign index_ge_13_right = 5'd13;
assign idx_between_9_13_reg_write_en = _guard6697;
assign idx_between_9_13_reg_clk = clk;
assign idx_between_9_13_reg_reset = reset;
assign idx_between_9_13_reg_in =
  _guard6698 ? idx_between_9_13_comb_out :
  _guard6701 ? 1'd0 :
  'x;
assign idx_between_1_5_comb_left = index_ge_1_out;
assign idx_between_1_5_comb_right = index_lt_5_out;
assign idx_between_10_14_reg_write_en = _guard6708;
assign idx_between_10_14_reg_clk = clk;
assign idx_between_10_14_reg_reset = reset;
assign idx_between_10_14_reg_in =
  _guard6709 ? idx_between_10_14_comb_out :
  _guard6712 ? 1'd0 :
  'x;
assign idx_between_16_24_reg_write_en = _guard6717;
assign idx_between_16_24_reg_clk = clk;
assign idx_between_16_24_reg_reset = reset;
assign idx_between_16_24_reg_in =
  _guard6718 ? idx_between_16_24_comb_out :
  _guard6721 ? 1'd0 :
  'x;
assign idx_between_11_15_reg_write_en = _guard6726;
assign idx_between_11_15_reg_clk = clk;
assign idx_between_11_15_reg_reset = reset;
assign idx_between_11_15_reg_in =
  _guard6729 ? 1'd0 :
  _guard6730 ? idx_between_11_15_comb_out :
  'x;
assign cond_wire1_in =
  _guard6733 ? cond1_out :
  _guard6734 ? idx_between_1_9_reg_out :
  1'd0;
assign cond8_write_en = _guard6735;
assign cond8_clk = clk;
assign cond8_reset = reset;
assign cond8_in =
  _guard6736 ? idx_between_14_15_reg_out :
  1'd0;
assign cond12_write_en = _guard6737;
assign cond12_clk = clk;
assign cond12_reset = reset;
assign cond12_in =
  _guard6738 ? idx_between_7_15_reg_out :
  1'd0;
assign cond28_write_en = _guard6739;
assign cond28_clk = clk;
assign cond28_reset = reset;
assign cond28_in =
  _guard6740 ? idx_between_18_19_reg_out :
  1'd0;
assign cond_wire28_in =
  _guard6741 ? idx_between_18_19_reg_out :
  _guard6744 ? cond28_out :
  1'd0;
assign cond_wire53_in =
  _guard6747 ? cond53_out :
  _guard6748 ? idx_between_5_13_reg_out :
  1'd0;
assign cond55_write_en = _guard6749;
assign cond55_clk = clk;
assign cond55_reset = reset;
assign cond55_in =
  _guard6750 ? idx_between_17_18_reg_out :
  1'd0;
assign cond_wire65_in =
  _guard6753 ? cond65_out :
  _guard6754 ? idx_between_8_16_reg_out :
  1'd0;
assign cond79_write_en = _guard6755;
assign cond79_clk = clk;
assign cond79_reset = reset;
assign cond79_in =
  _guard6756 ? idx_between_8_16_reg_out :
  1'd0;
assign cond_wire84_in =
  _guard6757 ? idx_between_17_18_reg_out :
  _guard6760 ? cond84_out :
  1'd0;
assign cond_wire88_in =
  _guard6763 ? cond88_out :
  _guard6764 ? idx_between_18_19_reg_out :
  1'd0;
assign cond_wire91_in =
  _guard6765 ? idx_between_11_19_reg_out :
  _guard6768 ? cond91_out :
  1'd0;
assign cond_wire109_in =
  _guard6769 ? idx_between_16_17_reg_out :
  _guard6772 ? cond109_out :
  1'd0;
assign cond_wire115_in =
  _guard6775 ? cond115_out :
  _guard6776 ? idx_between_6_14_reg_out :
  1'd0;
assign cond117_write_en = _guard6777;
assign cond117_clk = clk;
assign cond117_reset = reset;
assign cond117_in =
  _guard6778 ? idx_between_18_19_reg_out :
  1'd0;
assign cond_wire119_in =
  _guard6779 ? idx_between_7_15_reg_out :
  _guard6782 ? cond119_out :
  1'd0;
assign cond126_write_en = _guard6783;
assign cond126_clk = clk;
assign cond126_reset = reset;
assign cond126_in =
  _guard6784 ? idx_between_9_13_reg_out :
  1'd0;
assign cond135_write_en = _guard6785;
assign cond135_clk = clk;
assign cond135_reset = reset;
assign cond135_in =
  _guard6786 ? idx_between_11_19_reg_out :
  1'd0;
assign cond_wire141_in =
  _guard6789 ? cond141_out :
  _guard6790 ? idx_between_9_17_reg_out :
  1'd0;
assign cond153_write_en = _guard6791;
assign cond153_clk = clk;
assign cond153_reset = reset;
assign cond153_in =
  _guard6792 ? idx_between_12_20_reg_out :
  1'd0;
assign cond_wire158_in =
  _guard6793 ? idx_between_21_22_reg_out :
  _guard6796 ? cond158_out :
  1'd0;
assign cond_wire159_in =
  _guard6799 ? cond159_out :
  _guard6800 ? idx_between_10_14_reg_out :
  1'd0;
assign cond_wire169_in =
  _guard6803 ? cond169_out :
  _guard6804 ? idx_between_16_24_reg_out :
  1'd0;
assign cond171_write_en = _guard6805;
assign cond171_clk = clk;
assign cond171_reset = reset;
assign cond171_in =
  _guard6806 ? idx_between_5_13_reg_out :
  1'd0;
assign cond186_write_en = _guard6807;
assign cond186_clk = clk;
assign cond186_reset = reset;
assign cond186_in =
  _guard6808 ? idx_between_13_21_reg_out :
  1'd0;
assign cond_wire186_in =
  _guard6809 ? idx_between_13_21_reg_out :
  _guard6812 ? cond186_out :
  1'd0;
assign cond_wire196_in =
  _guard6815 ? cond196_out :
  _guard6816 ? idx_between_12_16_reg_out :
  1'd0;
assign cond213_write_en = _guard6817;
assign cond213_clk = clk;
assign cond213_reset = reset;
assign cond213_in =
  _guard6818 ? idx_between_9_13_reg_out :
  1'd0;
assign cond234_write_en = _guard6819;
assign cond234_clk = clk;
assign cond234_reset = reset;
assign cond234_in =
  _guard6820 ? idx_between_14_22_reg_out :
  1'd0;
assign cond_wire235_in =
  _guard6821 ? idx_between_18_26_reg_out :
  _guard6824 ? cond235_out :
  1'd0;
assign cond246_write_en = _guard6825;
assign cond246_clk = clk;
assign cond246_reset = reset;
assign cond246_in =
  _guard6826 ? idx_between_10_14_reg_out :
  1'd0;
assign cond_wire257_in =
  _guard6829 ? cond257_out :
  _guard6830 ? idx_between_24_25_reg_out :
  1'd0;
assign cond261_write_en = _guard6831;
assign cond261_clk = clk;
assign cond261_reset = reset;
assign cond261_in =
  _guard6832 ? idx_between_25_26_reg_out :
  1'd0;
assign wrapper_early_reset_static_seq_go_in = go;
assign left_0_1_write_en = _guard6835;
assign left_0_1_clk = clk;
assign left_0_1_reset = reset;
assign left_0_1_in = left_0_0_out;
assign top_0_7_write_en = _guard6841;
assign top_0_7_clk = clk;
assign top_0_7_reset = reset;
assign top_0_7_in = t7_read_data;
assign left_1_7_write_en = _guard6847;
assign left_1_7_clk = clk;
assign left_1_7_reset = reset;
assign left_1_7_in = left_1_6_out;
assign pe_2_2_mul_ready =
  _guard6853 ? 1'd1 :
  _guard6856 ? 1'd0 :
  1'd0;
assign pe_2_2_clk = clk;
assign pe_2_2_top =
  _guard6869 ? top_2_2_out :
  32'd0;
assign pe_2_2_left =
  _guard6882 ? left_2_2_out :
  32'd0;
assign pe_2_2_reset = reset;
assign pe_2_2_go = _guard6895;
assign pe_4_1_mul_ready =
  _guard6898 ? 1'd1 :
  _guard6901 ? 1'd0 :
  1'd0;
assign pe_4_1_clk = clk;
assign pe_4_1_top =
  _guard6914 ? top_4_1_out :
  32'd0;
assign pe_4_1_left =
  _guard6927 ? left_4_1_out :
  32'd0;
assign pe_4_1_reset = reset;
assign pe_4_1_go = _guard6940;
assign left_4_3_write_en = _guard6943;
assign left_4_3_clk = clk;
assign left_4_3_reset = reset;
assign left_4_3_in = left_4_2_out;
assign left_6_3_write_en = _guard6949;
assign left_6_3_clk = clk;
assign left_6_3_reset = reset;
assign left_6_3_in = left_6_2_out;
assign l2_add_left = 4'd1;
assign l2_add_right = l2_idx_out;
assign l5_idx_write_en = _guard6965;
assign l5_idx_clk = clk;
assign l5_idx_reset = reset;
assign l5_idx_in =
  _guard6968 ? 4'd0 :
  _guard6971 ? l5_add_out :
  'x;
assign l6_add_left = 4'd1;
assign l6_add_right = l6_idx_out;
assign index_lt_26_left = idx_add_out;
assign index_lt_26_right = 5'd26;
assign index_lt_23_left = idx_add_out;
assign index_lt_23_right = 5'd23;
assign idx_between_1_9_reg_write_en = _guard6986;
assign idx_between_1_9_reg_clk = clk;
assign idx_between_1_9_reg_reset = reset;
assign idx_between_1_9_reg_in =
  _guard6987 ? idx_between_1_9_comb_out :
  _guard6990 ? 1'd0 :
  'x;
assign index_lt_14_left = idx_add_out;
assign index_lt_14_right = 5'd14;
assign idx_between_6_14_comb_left = index_ge_6_out;
assign idx_between_6_14_comb_right = index_lt_14_out;
assign index_lt_25_left = idx_add_out;
assign index_lt_25_right = 5'd25;
assign idx_between_3_11_reg_write_en = _guard7001;
assign idx_between_3_11_reg_clk = clk;
assign idx_between_3_11_reg_reset = reset;
assign idx_between_3_11_reg_in =
  _guard7002 ? idx_between_3_11_comb_out :
  _guard7005 ? 1'd0 :
  'x;
assign idx_between_2_6_reg_write_en = _guard7010;
assign idx_between_2_6_reg_clk = clk;
assign idx_between_2_6_reg_reset = reset;
assign idx_between_2_6_reg_in =
  _guard7013 ? 1'd0 :
  _guard7014 ? idx_between_2_6_comb_out :
  'x;
assign idx_between_2_6_comb_left = index_ge_2_out;
assign idx_between_2_6_comb_right = index_lt_6_out;
assign cond_wire14_in =
  _guard7019 ? cond14_out :
  _guard7020 ? idx_between_3_11_reg_out :
  1'd0;
assign cond_wire21_in =
  _guard7021 ? idx_between_5_13_reg_out :
  _guard7024 ? cond21_out :
  1'd0;
assign cond38_write_en = _guard7025;
assign cond38_clk = clk;
assign cond38_reset = reset;
assign cond38_in =
  _guard7026 ? idx_between_20_21_reg_out :
  1'd0;
assign cond42_write_en = _guard7027;
assign cond42_clk = clk;
assign cond42_reset = reset;
assign cond42_in =
  _guard7028 ? idx_between_6_14_reg_out :
  1'd0;
assign cond_wire51_in =
  _guard7029 ? idx_between_16_17_reg_out :
  _guard7032 ? cond51_out :
  1'd0;
assign cond59_write_en = _guard7033;
assign cond59_clk = clk;
assign cond59_reset = reset;
assign cond59_in =
  _guard7034 ? idx_between_18_19_reg_out :
  1'd0;
assign cond_wire78_in =
  _guard7035 ? idx_between_4_12_reg_out :
  _guard7038 ? cond78_out :
  1'd0;
assign cond_wire79_in =
  _guard7039 ? idx_between_8_16_reg_out :
  _guard7042 ? cond79_out :
  1'd0;
assign cond85_write_en = _guard7043;
assign cond85_clk = clk;
assign cond85_reset = reset;
assign cond85_in =
  _guard7044 ? idx_between_6_10_reg_out :
  1'd0;
assign cond_wire102_in =
  _guard7045 ? idx_between_10_18_reg_out :
  _guard7048 ? cond102_out :
  1'd0;
assign cond111_write_en = _guard7049;
assign cond111_clk = clk;
assign cond111_reset = reset;
assign cond111_in =
  _guard7050 ? idx_between_5_13_reg_out :
  1'd0;
assign cond_wire124_in =
  _guard7053 ? cond124_out :
  _guard7054 ? idx_between_12_20_reg_out :
  1'd0;
assign cond142_write_en = _guard7055;
assign cond142_clk = clk;
assign cond142_reset = reset;
assign cond142_in =
  _guard7056 ? idx_between_17_18_reg_out :
  1'd0;
assign cond157_write_en = _guard7057;
assign cond157_clk = clk;
assign cond157_reset = reset;
assign cond157_in =
  _guard7058 ? idx_between_13_21_reg_out :
  1'd0;
assign cond_wire166_in =
  _guard7059 ? idx_between_23_24_reg_out :
  _guard7062 ? cond166_out :
  1'd0;
assign cond_wire180_in =
  _guard7065 ? cond180_out :
  _guard7066 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire183_in =
  _guard7067 ? idx_between_20_21_reg_out :
  _guard7070 ? cond183_out :
  1'd0;
assign cond_wire188_in =
  _guard7073 ? cond188_out :
  _guard7074 ? idx_between_10_14_reg_out :
  1'd0;
assign cond200_write_en = _guard7075;
assign cond200_clk = clk;
assign cond200_reset = reset;
assign cond200_in =
  _guard7076 ? idx_between_13_17_reg_out :
  1'd0;
assign cond_wire202_in =
  _guard7079 ? cond202_out :
  _guard7080 ? idx_between_17_25_reg_out :
  1'd0;
assign cond_wire211_in =
  _guard7083 ? cond211_out :
  _guard7084 ? idx_between_12_20_reg_out :
  1'd0;
assign cond_wire215_in =
  _guard7087 ? cond215_out :
  _guard7088 ? idx_between_13_21_reg_out :
  1'd0;
assign cond_wire226_in =
  _guard7091 ? cond226_out :
  _guard7092 ? idx_between_12_20_reg_out :
  1'd0;
assign cond_wire227_in =
  _guard7095 ? cond227_out :
  _guard7096 ? idx_between_16_24_reg_out :
  1'd0;
assign cond253_write_en = _guard7097;
assign cond253_clk = clk;
assign cond253_reset = reset;
assign cond253_in =
  _guard7098 ? idx_between_23_24_reg_out :
  1'd0;
assign cond254_write_en = _guard7099;
assign cond254_clk = clk;
assign cond254_reset = reset;
assign cond254_in =
  _guard7100 ? idx_between_12_16_reg_out :
  1'd0;
assign cond_wire254_in =
  _guard7101 ? idx_between_12_16_reg_out :
  _guard7104 ? cond254_out :
  1'd0;
// COMPONENT END: main
endmodule

