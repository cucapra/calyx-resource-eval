
module std_fp_mult_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    input  logic             go,
    input  logic             clk,
    output logic [WIDTH-1:0] out,
    output logic             done
);
  logic [WIDTH-1:0]          rtmp;
  logic [WIDTH-1:0]          ltmp;
  logic [(WIDTH << 1) - 1:0] out_tmp;
  reg done_buf[1:0];
  always_ff @(posedge clk) begin
    if (go) begin
      rtmp <= right;
      ltmp <= left;
      out_tmp <= ltmp * rtmp;
      out <= out_tmp[(WIDTH << 1) - INT_WIDTH - 1 : WIDTH - INT_WIDTH];

      done <= done_buf[1];
      done_buf[0] <= 1'b1;
      done_buf[1] <= done_buf[0];
    end else begin
      rtmp <= 0;
      ltmp <= 0;
      out_tmp <= 0;
      out <= 0;

      done <= 0;
      done_buf[0] <= 0;
      done_buf[1] <= 0;
    end
  end
endmodule

module std_fp_add #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  assign out = left + right;
endmodule

module std_fp_sub #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module std_fp_gt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic             out
);
  assign out = left > right;
endmodule

module std_fp_add_dwidth #(
    parameter WIDTH1 = 32,
    parameter WIDTH2 = 32,
    parameter INT_WIDTH1 = 8,
    parameter FRACT_WIDTH1 = 24,
    parameter INT_WIDTH2 = 4,
    parameter FRACT_WIDTH2 = 28,
    parameter OUT_WIDTH = 36
) (
    input  logic [   WIDTH1-1:0] left,
    input  logic [   WIDTH2-1:0] right,
    output logic [OUT_WIDTH-1:0] out
);

  localparam BIG_INT = (INT_WIDTH1 >= INT_WIDTH2) ? INT_WIDTH1 : INT_WIDTH2;
  localparam BIG_FRACT = (FRACT_WIDTH1 >= FRACT_WIDTH2) ? FRACT_WIDTH1 : FRACT_WIDTH2;

  if (BIG_INT + BIG_FRACT != OUT_WIDTH)
    $error("std_fp_add_dwidth: Given output width not equal to computed output width");

  logic [INT_WIDTH1-1:0] left_int;
  logic [INT_WIDTH2-1:0] right_int;
  logic [FRACT_WIDTH1-1:0] left_fract;
  logic [FRACT_WIDTH2-1:0] right_fract;

  logic [BIG_INT-1:0] mod_right_int;
  logic [BIG_FRACT-1:0] mod_left_fract;

  logic [BIG_INT-1:0] whole_int;
  logic [BIG_FRACT-1:0] whole_fract;

  assign {left_int, left_fract} = left;
  assign {right_int, right_fract} = right;

  assign mod_left_fract = left_fract * (2 ** (FRACT_WIDTH2 - FRACT_WIDTH1));

  always_comb begin
    if ((mod_left_fract + right_fract) >= 2 ** FRACT_WIDTH2) begin
      whole_int = left_int + right_int + 1;
      whole_fract = mod_left_fract + right_fract - 2 ** FRACT_WIDTH2;
    end else begin
      whole_int = left_int + right_int;
      whole_fract = mod_left_fract + right_fract;
    end
  end

  assign out = {whole_int, whole_fract};
endmodule

/// ========================= Unsynthesizable primitives =====================

module std_fp_mult #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  logic [2*WIDTH-2:0] result;

  assign result = left * right;
  assign out = result[WIDTH+FRACT_WIDTH-1:FRACT_WIDTH];
endmodule

module std_fp_div #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  logic [2*WIDTH-2:0] result;

  assign result = left / right;
  assign out = result[WIDTH+FRACT_WIDTH-1:FRACT_WIDTH];
endmodule
module std_fp_smult_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  signed       [WIDTH-1:0] left,
    input  signed       [WIDTH-1:0] right,
    input  logic                    go,
    input  logic                    clk,
    output logic signed [WIDTH-1:0] out,
    output logic                    done
);
  logic signed [WIDTH-1:0] rtmp;
  logic signed [WIDTH-1:0] ltmp;
  logic signed [(WIDTH << 1) - 1:0] out_tmp;
  reg done_buf[1:0];
  always_ff @(posedge clk) begin
    if (go) begin
      ltmp <= left;
      rtmp <= right;
      // Sign extend by the first bit for the operands.
      out_tmp <= $signed(
                   { {WIDTH{ltmp[WIDTH-1]}}, ltmp} *
                   { {WIDTH{rtmp[WIDTH-1]}}, rtmp}
                 );
      out <= out_tmp[(WIDTH << 1) - INT_WIDTH - 1: WIDTH - INT_WIDTH];

      done <= done_buf[1];
      done_buf[0] <= 1'b1;
      done_buf[1] <= done_buf[0];
    end else begin
      rtmp <= 0;
      ltmp <= 0;
      out_tmp <= 0;
      out <= 0;

      done <= 0;
      done_buf[0] <= 0;
      done_buf[1] <= 0;
    end
  end
endmodule

module std_fp_sadd #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left + right);
endmodule

module std_fp_ssub #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);

  assign out = $signed(left - right);
endmodule

module std_fp_sadd_dwidth #(
    parameter WIDTH1 = 32,
    parameter WIDTH2 = 32,
    parameter INT_WIDTH1 = 8,
    parameter FRACT_WIDTH1 = 24,
    parameter INT_WIDTH2 = 4,
    parameter FRACT_WIDTH2 = 28,
    parameter OUT_WIDTH = 36
) (
    input  logic [   WIDTH1-1:0] left,
    input  logic [   WIDTH2-1:0] right,
    output logic [OUT_WIDTH-1:0] out
);

  logic signed [INT_WIDTH1-1:0] left_int;
  logic signed [INT_WIDTH2-1:0] right_int;
  logic [FRACT_WIDTH1-1:0] left_fract;
  logic [FRACT_WIDTH2-1:0] right_fract;

  localparam BIG_INT = (INT_WIDTH1 >= INT_WIDTH2) ? INT_WIDTH1 : INT_WIDTH2;
  localparam BIG_FRACT = (FRACT_WIDTH1 >= FRACT_WIDTH2) ? FRACT_WIDTH1 : FRACT_WIDTH2;

  logic [BIG_INT-1:0] mod_right_int;
  logic [BIG_FRACT-1:0] mod_left_fract;

  logic [BIG_INT-1:0] whole_int;
  logic [BIG_FRACT-1:0] whole_fract;

  assign {left_int, left_fract} = left;
  assign {right_int, right_fract} = right;

  assign mod_left_fract = left_fract * (2 ** (FRACT_WIDTH2 - FRACT_WIDTH1));

  always_comb begin
    if ((mod_left_fract + right_fract) >= 2 ** FRACT_WIDTH2) begin
      whole_int = $signed(left_int + right_int + 1);
      whole_fract = mod_left_fract + right_fract - 2 ** FRACT_WIDTH2;
    end else begin
      whole_int = $signed(left_int + right_int);
      whole_fract = mod_left_fract + right_fract;
    end
  end

  assign out = {whole_int, whole_fract};
endmodule

module std_fp_sgt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  logic signed [WIDTH-1:0] left,
    input  logic signed [WIDTH-1:0] right,
    output logic signed             out
);
  assign out = $signed(left > right);
endmodule

module std_fp_smult #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);

  logic [2*WIDTH-2:0] result;

  assign result = $signed(left * right);
  assign out = result[WIDTH+FRACT_WIDTH-1:FRACT_WIDTH];
endmodule

module std_fp_sdiv #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 8,
    parameter FRACT_WIDTH = 24
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);

  logic [2*WIDTH-2:0] result;

  assign result = $signed(left / right);
  assign out = result[WIDTH+FRACT_WIDTH-1:FRACT_WIDTH];
endmodule

/* verilator lint_off WIDTH */
module std_div_pipe #(
    parameter width = 32
) (
    input                    clk,
    input                    go,
    input        [width-1:0] left,
    input        [width-1:0] right,
    output logic [width-1:0] out_remainder,
    output logic [width-1:0] out_quotient,
    output logic             done
);

  logic [width-1:0] dividend;
  logic [(width-1)*2:0] divisor;
  logic [width-1:0] quotient;
  logic [width-1:0] quotient_msk;
  logic start, running, finished;

  assign start = go && !running;
  assign finished = !quotient_msk && running;

  always @(posedge clk) begin
    if (!go) begin
      running <= 0;
      done <= 0;
      out_remainder <= 0;
      out_quotient <= 0;
    end else if (start && left == 0) begin
      out_remainder <= 0;
      out_quotient <= 0;
      done <= 1;
    end

    if (start) begin
      running <= 1;
      dividend <= left;
      divisor <= right << width - 1;
      quotient <= 0;
      quotient_msk <= 1 << width - 1;
    end else if (finished) begin
      running <= 0;
      done <= 1;
      out_remainder <= dividend;
      out_quotient <= quotient;
    end else begin
      if (divisor <= dividend) begin
        dividend <= dividend - divisor;
        quotient <= quotient | quotient_msk;
      end
      divisor <= divisor >> 1;
      quotient_msk <= quotient_msk >> 1;
    end
  end

  `ifdef VERILATOR
    // Simulation self test against unsynthesizable implementation.
    always @(posedge clk) begin
      if (finished && dividend != $unsigned(left % right))
        $error(
          "\nstd_div_pipe (Remainder): Computed and golden outputs do not match!\n",
          "left: %0d", $unsigned(left),
          "  right: %0d\n", $unsigned(right),
          "expected: %0d", $unsigned(left % right),
          "  computed: %0d", $unsigned(dividend)
        );
      if (finished && quotient != $unsigned(left / right))
        $error(
          "\nstd_div_pipe (Quotient): Computed and golden outputs do not match!\n",
          "left: %0d", $unsigned(left),
          "  right: %0d\n", $unsigned(right),
          "expected: %0d", $unsigned(left / right),
          "  computed: %0d", $unsigned(quotient)
        );
    end
  `endif
endmodule

module std_mult_pipe #(
    parameter width = 32
) (
    input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    input  logic             go,
    input  logic             clk,
    output logic [width-1:0] out,
    output logic             done
);
  logic [width-1:0] rtmp;
  logic [width-1:0] ltmp;
  logic [width-1:0] out_tmp;
  reg done_buf[1:0];
  always_ff @(posedge clk) begin
    if (go) begin
      rtmp <= right;
      ltmp <= left;
      out_tmp <= rtmp * ltmp;
      out <= out_tmp;

      done <= done_buf[1];
      done_buf[0] <= 1'b1;
      done_buf[1] <= done_buf[0];
    end else begin
      rtmp <= 0;
      ltmp <= 0;
      out_tmp <= 0;
      out <= 0;

      done <= 0;
      done_buf[0] <= 0;
      done_buf[1] <= 0;
    end
  end
endmodule

// ===============Signed operations that wrap unsigned ones ===============

/* verilator lint_off WIDTH */
module std_sdiv_pipe #(
    parameter width = 32
) (
    input                     clk,
    input                     go,
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output logic  [width-1:0] out_quotient,
    output logic  [width-1:0] out_remainder,
    output logic              done
);

  logic signed [width-1:0] left_abs;
  logic signed [width-1:0] right_abs;
  logic signed [width-1:0] comp_out_q;
  logic signed [width-1:0] comp_out_r;

  assign right_abs = right[width-1] == 1 ? -right : right;
  assign left_abs = left[width-1] == 1 ? -left : left;
  assign out_quotient =
    (left[width-1] == 1) ^ (right[width-1] == 1) ? -comp_out_q : comp_out_q;
  assign out_remainder = left[width-1] == 1 ? $signed(right - comp_out_r) : comp_out_r;

  std_div_pipe #(
    .width(width)
  ) comp (
    .clk(clk),
    .done(done),
    .go(go),
    .left(left_abs),
    .right(right_abs),
    .out_quotient(comp_out_q),
    .out_remainder(comp_out_r)
  );

  `ifdef VERILATOR
    // Simulation self test against unsynthesizable implementation.
    always @(posedge clk) begin
      if (done && out_quotient != $signed(left / right))
        $error(
          "\nstd_sdiv_pipe (Quotient): Computed and golden outputs do not match!\n",
          "left: %0d", left,
          "  right: %0d\n", right,
          "expected: %0d", $signed(left / right),
          "  computed: %0d", $signed(out_quotient)
        );
      if (done && out_remainder != $signed(((left % right) + right) % right))
        $error(
          "\nstd_sdiv_pipe (Remainder): Computed and golden outputs do not match!\n",
          "left: %0d", left,
          "  right: %0d\n", right,
          "expected: %0d", $signed(((left % right) + right) % right),
          "  computed: %0d", $signed(out_remainder)
        );
    end
  `endif
endmodule


//==================== Unsynthesizable primitives =========================
module std_mult #(
    parameter width = 32
) (
    input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    output logic [width-1:0] out
);
  assign out = left * right;
endmodule

module std_div #(
    parameter width = 32
) (
    input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    output logic [width-1:0] out
);
  assign out = left / right;
endmodule

module std_mod #(
    parameter width = 32
) (
    input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    output logic [width-1:0] out
);
  assign out = left % right;
endmodule
/**
* Signed arthimetic primitives for FuTIL.
*/

module std_slsh #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed [width-1:0] out
);
  assign out = left <<< right;
endmodule

module std_srsh #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed [width-1:0] out
);
  assign out = left >>> right;
endmodule

module std_sadd #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed [width-1:0] out
);
  assign out = $signed(left + right);
endmodule

module std_ssub #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed [width-1:0] out
);
  assign out = $signed(left - right);
endmodule

module std_smult_pipe #(
    parameter width = 32
) (
    input  logic                    go,
    input  logic                    clk,
    input  signed       [width-1:0] left,
    input  signed       [width-1:0] right,
    output logic signed [width-1:0] out,
    output logic                    done
);
  logic signed [width-1:0] rtmp;
  logic signed [width-1:0] ltmp;
  logic signed [width-1:0] out_tmp;
  logic done_buf[1:0];

  always_ff @(posedge clk) begin
    if (go) begin
      rtmp <= right;
      ltmp <= left;
      out_tmp <= $signed(rtmp * ltmp);
      out <= out_tmp;

      done <= done_buf[1];
      done_buf[0] <= 1'b1;
      done_buf[1] <= done_buf[0];
    end else begin
      rtmp <= 0;
      ltmp <= 0;
      out_tmp <= 0;
      out <= 0;

      done <= 0;
      done_buf[0] <= 0;
      done_buf[1] <= 0;
    end
  end
endmodule

module std_sgt #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed             out
);
  assign out = $signed(left > right);
endmodule

module std_slt #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed             out
);
  assign out = $signed(left < right);
endmodule

module std_seq #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed             out
);
  assign out = $signed(left == right);
endmodule

module std_sneq #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed             out
);
  assign out = $signed(left != right);
endmodule

module std_sge #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed             out
);
  assign out = $signed(left >= right);
endmodule

module std_sle #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed             out
);
  assign out = $signed(left <= right);
endmodule

module std_sdiv #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed [width-1:0] out
);
  assign out = $signed(left / right);
endmodule

module std_smod #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed [width-1:0] out
);
  assign out = $signed(left % right);
endmodule


module std_smult #(
    parameter width = 32
) (
    input  signed [width-1:0] left,
    input  signed [width-1:0] right,
    output signed [width-1:0] out
);
  assign out = $signed(left * right);
endmodule

/**
 * Core primitives for FuTIL.
 * Implements core primitives used by the compiler.
 *
 * Conventions:
 * - All parameter names must be SNAKE_CASE and all caps.
 * - Port names must be snake_case, no caps.
 */
`default_nettype none

module std_mem_d1 #(
    parameter width = 32,
    parameter size = 16,
    parameter idx_size = 4
) (
   input wire                logic [idx_size-1:0] addr0,
   input wire                logic [ width-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   output logic [ width-1:0] read_data,
   output logic              done
);

  logic [width-1:0] mem[size-1:0];

  /* verilator lint_off WIDTH */
  assign read_data = mem[addr0];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0] <= write_data;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module std_mem_d2 #(
    parameter width = 32,
    parameter d0_size = 16,
    parameter d1_size = 16,
    parameter d0_idx_size = 4,
    parameter d1_idx_size = 4
) (
   input wire                logic [d0_idx_size-1:0] addr0,
   input wire                logic [d1_idx_size-1:0] addr1,
   input wire                logic [ width-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   output logic [ width-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [width-1:0] mem[d0_size-1:0][d1_size-1:0];

  assign read_data = mem[addr0][addr1];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0][addr1] <= write_data;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module std_mem_d3 #(
    parameter width = 32,
    parameter d0_size = 16,
    parameter d1_size = 16,
    parameter d2_size = 16,
    parameter d0_idx_size = 4,
    parameter d1_idx_size = 4,
    parameter d2_idx_size = 4
) (
   input wire                logic [d0_idx_size-1:0] addr0,
   input wire                logic [d1_idx_size-1:0] addr1,
   input wire                logic [d2_idx_size-1:0] addr2,
   input wire                logic [ width-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   output logic [ width-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [width-1:0] mem[d0_size-1:0][d1_size-1:0][d2_size-1:0];

  assign read_data = mem[addr0][addr1][addr2];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0][addr1][addr2] <= write_data;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module std_mem_d4 #(
    parameter width = 32,
    parameter d0_size = 16,
    parameter d1_size = 16,
    parameter d2_size = 16,
    parameter d3_size = 16,
    parameter d0_idx_size = 4,
    parameter d1_idx_size = 4,
    parameter d2_idx_size = 4,
    parameter d3_idx_size = 4
) (
   input wire                logic [d0_idx_size-1:0] addr0,
   input wire                logic [d1_idx_size-1:0] addr1,
   input wire                logic [d2_idx_size-1:0] addr2,
   input wire                logic [d3_idx_size-1:0] addr3,
   input wire                logic [ width-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   output logic [ width-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [width-1:0] mem[d0_size-1:0][d1_size-1:0][d2_size-1:0][d3_size-1:0];

  assign read_data = mem[addr0][addr1][addr2][addr3];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0][addr1][addr2][addr3] <= write_data;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module std_reg #(
    parameter width = 32
) (
   input wire [ width-1:0]    in,
   input wire                 write_en,
   input wire                 clk,
    // output
   output logic [width - 1:0] out,
   output logic               done
);

  always_ff @(posedge clk) begin
    if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module std_const #(
    parameter width = 32,
    parameter value = 0
) (
   output logic [width - 1:0] out
);
  assign out = value;
endmodule

module std_slice #(
    parameter in_width  = 32,
    parameter out_width = 32
) (
   input wire                   logic [ in_width-1:0] in,
   output logic [out_width-1:0] out
);
  assign out = in[out_width-1:0];

  `ifdef VERILATOR
    always_comb begin
      if (in_width < out_width)
        $error(
          "std_slice: Input width less than output width\n",
          "in_width: %0d", in_width,
          "out_width: %0d", out_width
        );
    end
  `endif
endmodule

module std_pad #(
    parameter in_width  = 32,
    parameter out_width = 32
) (
   input wire                   logic [ in_width-1:0] in,
   output logic [out_width-1:0] out
);
  localparam EXTEND = out_width - in_width;
  assign out = { {EXTEND {1'b0}}, in};

  `ifdef VERILATOR
    always_comb begin
      if (in_width > out_width)
        $error(
          "std_pad: Output width less than input width\n",
          "in_width: %0d", in_width,
          "out_width: %0d", out_width
        );
    end
  `endif
endmodule

module std_lsh #(
    parameter width = 32
) (
   input wire               logic [width-1:0] left,
   input wire               logic [width-1:0] right,
   output logic [width-1:0] out
);
  assign out = left << right;
endmodule

module std_rsh #(
    parameter width = 32
) (
   input wire               logic [width-1:0] left,
   input wire               logic [width-1:0] right,
   output logic [width-1:0] out
);
  assign out = left >> right;
endmodule

module std_add #(
    parameter width = 32
) (
   input wire               logic [width-1:0] left,
   input wire               logic [width-1:0] right,
   output logic [width-1:0] out
);
  assign out = left + right;
endmodule

module std_sub #(
    parameter width = 32
) (
   input wire               logic [width-1:0] left,
   input wire               logic [width-1:0] right,
   output logic [width-1:0] out
);
  assign out = left - right;
endmodule

module std_not #(
    parameter width = 32
) (
   input wire               logic [width-1:0] in,
   output logic [width-1:0] out
);
  assign out = ~in;
endmodule

module std_and #(
    parameter width = 32
) (
   input wire               logic [width-1:0] left,
   input wire               logic [width-1:0] right,
   output logic [width-1:0] out
);
  assign out = left & right;
endmodule

module std_or #(
    parameter width = 32
) (
   input wire               logic [width-1:0] left,
   input wire               logic [width-1:0] right,
   output logic [width-1:0] out
);
  assign out = left | right;
endmodule

module std_xor #(
    parameter width = 32
) (
   input wire               logic [width-1:0] left,
   input wire               logic [width-1:0] right,
   output logic [width-1:0] out
);
  assign out = left ^ right;
endmodule

module std_gt #(
    parameter width = 32
) (
   input wire   logic [width-1:0] left,
   input wire   logic [width-1:0] right,
   output logic out
);
  assign out = left > right;
endmodule

module std_lt #(
    parameter width = 32
) (
   input wire   logic [width-1:0] left,
   input wire   logic [width-1:0] right,
   output logic out
);
  assign out = left < right;
endmodule

module std_eq #(
    parameter width = 32
) (
   input wire   logic [width-1:0] left,
   input wire   logic [width-1:0] right,
   output logic out
);
  assign out = left == right;
endmodule

module std_neq #(
    parameter width = 32
) (
   input wire   logic [width-1:0] left,
   input wire   logic [width-1:0] right,
   output logic out
);
  assign out = left != right;
endmodule

module std_ge #(
    parameter width = 32
) (
    input wire   logic [width-1:0] left,
    input wire   logic [width-1:0] right,
    output logic out
);
  assign out = left >= right;
endmodule

module std_le #(
    parameter width = 32
) (
   input wire   logic [width-1:0] left,
   input wire   logic [width-1:0] right,
   output logic out
);
  assign out = left <= right;
endmodule

`default_nettype wire
module main (
    input logic go,
    input logic clk,
    output logic done,
    output logic [4:0] t0_addr0,
    output logic [31:0] t0_write_data,
    output logic t0_write_en,
    output logic t0_clk,
    input logic [31:0] t0_read_data,
    input logic t0_done,
    output logic [4:0] t1_addr0,
    output logic [31:0] t1_write_data,
    output logic t1_write_en,
    output logic t1_clk,
    input logic [31:0] t1_read_data,
    input logic t1_done,
    output logic [4:0] t2_addr0,
    output logic [31:0] t2_write_data,
    output logic t2_write_en,
    output logic t2_clk,
    input logic [31:0] t2_read_data,
    input logic t2_done,
    output logic [4:0] t3_addr0,
    output logic [31:0] t3_write_data,
    output logic t3_write_en,
    output logic t3_clk,
    input logic [31:0] t3_read_data,
    input logic t3_done,
    output logic [4:0] t4_addr0,
    output logic [31:0] t4_write_data,
    output logic t4_write_en,
    output logic t4_clk,
    input logic [31:0] t4_read_data,
    input logic t4_done,
    output logic [4:0] t5_addr0,
    output logic [31:0] t5_write_data,
    output logic t5_write_en,
    output logic t5_clk,
    input logic [31:0] t5_read_data,
    input logic t5_done,
    output logic [4:0] t6_addr0,
    output logic [31:0] t6_write_data,
    output logic t6_write_en,
    output logic t6_clk,
    input logic [31:0] t6_read_data,
    input logic t6_done,
    output logic [4:0] t7_addr0,
    output logic [31:0] t7_write_data,
    output logic t7_write_en,
    output logic t7_clk,
    input logic [31:0] t7_read_data,
    input logic t7_done,
    output logic [4:0] t8_addr0,
    output logic [31:0] t8_write_data,
    output logic t8_write_en,
    output logic t8_clk,
    input logic [31:0] t8_read_data,
    input logic t8_done,
    output logic [4:0] t9_addr0,
    output logic [31:0] t9_write_data,
    output logic t9_write_en,
    output logic t9_clk,
    input logic [31:0] t9_read_data,
    input logic t9_done,
    output logic [4:0] t10_addr0,
    output logic [31:0] t10_write_data,
    output logic t10_write_en,
    output logic t10_clk,
    input logic [31:0] t10_read_data,
    input logic t10_done,
    output logic [4:0] t11_addr0,
    output logic [31:0] t11_write_data,
    output logic t11_write_en,
    output logic t11_clk,
    input logic [31:0] t11_read_data,
    input logic t11_done,
    output logic [4:0] t12_addr0,
    output logic [31:0] t12_write_data,
    output logic t12_write_en,
    output logic t12_clk,
    input logic [31:0] t12_read_data,
    input logic t12_done,
    output logic [4:0] t13_addr0,
    output logic [31:0] t13_write_data,
    output logic t13_write_en,
    output logic t13_clk,
    input logic [31:0] t13_read_data,
    input logic t13_done,
    output logic [4:0] t14_addr0,
    output logic [31:0] t14_write_data,
    output logic t14_write_en,
    output logic t14_clk,
    input logic [31:0] t14_read_data,
    input logic t14_done,
    output logic [4:0] t15_addr0,
    output logic [31:0] t15_write_data,
    output logic t15_write_en,
    output logic t15_clk,
    input logic [31:0] t15_read_data,
    input logic t15_done,
    output logic [4:0] l0_addr0,
    output logic [31:0] l0_write_data,
    output logic l0_write_en,
    output logic l0_clk,
    input logic [31:0] l0_read_data,
    input logic l0_done,
    output logic [4:0] l1_addr0,
    output logic [31:0] l1_write_data,
    output logic l1_write_en,
    output logic l1_clk,
    input logic [31:0] l1_read_data,
    input logic l1_done,
    output logic [4:0] l2_addr0,
    output logic [31:0] l2_write_data,
    output logic l2_write_en,
    output logic l2_clk,
    input logic [31:0] l2_read_data,
    input logic l2_done,
    output logic [4:0] l3_addr0,
    output logic [31:0] l3_write_data,
    output logic l3_write_en,
    output logic l3_clk,
    input logic [31:0] l3_read_data,
    input logic l3_done,
    output logic [4:0] l4_addr0,
    output logic [31:0] l4_write_data,
    output logic l4_write_en,
    output logic l4_clk,
    input logic [31:0] l4_read_data,
    input logic l4_done,
    output logic [4:0] l5_addr0,
    output logic [31:0] l5_write_data,
    output logic l5_write_en,
    output logic l5_clk,
    input logic [31:0] l5_read_data,
    input logic l5_done,
    output logic [4:0] l6_addr0,
    output logic [31:0] l6_write_data,
    output logic l6_write_en,
    output logic l6_clk,
    input logic [31:0] l6_read_data,
    input logic l6_done,
    output logic [4:0] l7_addr0,
    output logic [31:0] l7_write_data,
    output logic l7_write_en,
    output logic l7_clk,
    input logic [31:0] l7_read_data,
    input logic l7_done,
    output logic [4:0] l8_addr0,
    output logic [31:0] l8_write_data,
    output logic l8_write_en,
    output logic l8_clk,
    input logic [31:0] l8_read_data,
    input logic l8_done,
    output logic [4:0] l9_addr0,
    output logic [31:0] l9_write_data,
    output logic l9_write_en,
    output logic l9_clk,
    input logic [31:0] l9_read_data,
    input logic l9_done,
    output logic [4:0] l10_addr0,
    output logic [31:0] l10_write_data,
    output logic l10_write_en,
    output logic l10_clk,
    input logic [31:0] l10_read_data,
    input logic l10_done,
    output logic [4:0] l11_addr0,
    output logic [31:0] l11_write_data,
    output logic l11_write_en,
    output logic l11_clk,
    input logic [31:0] l11_read_data,
    input logic l11_done,
    output logic [4:0] l12_addr0,
    output logic [31:0] l12_write_data,
    output logic l12_write_en,
    output logic l12_clk,
    input logic [31:0] l12_read_data,
    input logic l12_done,
    output logic [4:0] l13_addr0,
    output logic [31:0] l13_write_data,
    output logic l13_write_en,
    output logic l13_clk,
    input logic [31:0] l13_read_data,
    input logic l13_done,
    output logic [4:0] l14_addr0,
    output logic [31:0] l14_write_data,
    output logic l14_write_en,
    output logic l14_clk,
    input logic [31:0] l14_read_data,
    input logic l14_done,
    output logic [4:0] l15_addr0,
    output logic [31:0] l15_write_data,
    output logic l15_write_en,
    output logic l15_clk,
    input logic [31:0] l15_read_data,
    input logic l15_done,
    output logic [4:0] out_mem_addr0,
    output logic [4:0] out_mem_addr1,
    output logic [31:0] out_mem_write_data,
    output logic out_mem_write_en,
    output logic out_mem_clk,
    input logic [31:0] out_mem_read_data,
    input logic out_mem_done
);
    logic [4:0] t0_idx_in;
    logic t0_idx_write_en;
    logic t0_idx_clk;
    logic [4:0] t0_idx_out;
    logic t0_idx_done;
    logic [4:0] t0_add_left;
    logic [4:0] t0_add_right;
    logic [4:0] t0_add_out;
    logic [4:0] t1_idx_in;
    logic t1_idx_write_en;
    logic t1_idx_clk;
    logic [4:0] t1_idx_out;
    logic t1_idx_done;
    logic [4:0] t1_add_left;
    logic [4:0] t1_add_right;
    logic [4:0] t1_add_out;
    logic [4:0] t2_idx_in;
    logic t2_idx_write_en;
    logic t2_idx_clk;
    logic [4:0] t2_idx_out;
    logic t2_idx_done;
    logic [4:0] t2_add_left;
    logic [4:0] t2_add_right;
    logic [4:0] t2_add_out;
    logic [4:0] t3_idx_in;
    logic t3_idx_write_en;
    logic t3_idx_clk;
    logic [4:0] t3_idx_out;
    logic t3_idx_done;
    logic [4:0] t3_add_left;
    logic [4:0] t3_add_right;
    logic [4:0] t3_add_out;
    logic [4:0] t4_idx_in;
    logic t4_idx_write_en;
    logic t4_idx_clk;
    logic [4:0] t4_idx_out;
    logic t4_idx_done;
    logic [4:0] t4_add_left;
    logic [4:0] t4_add_right;
    logic [4:0] t4_add_out;
    logic [4:0] t5_idx_in;
    logic t5_idx_write_en;
    logic t5_idx_clk;
    logic [4:0] t5_idx_out;
    logic t5_idx_done;
    logic [4:0] t5_add_left;
    logic [4:0] t5_add_right;
    logic [4:0] t5_add_out;
    logic [4:0] t6_idx_in;
    logic t6_idx_write_en;
    logic t6_idx_clk;
    logic [4:0] t6_idx_out;
    logic t6_idx_done;
    logic [4:0] t6_add_left;
    logic [4:0] t6_add_right;
    logic [4:0] t6_add_out;
    logic [4:0] t7_idx_in;
    logic t7_idx_write_en;
    logic t7_idx_clk;
    logic [4:0] t7_idx_out;
    logic t7_idx_done;
    logic [4:0] t7_add_left;
    logic [4:0] t7_add_right;
    logic [4:0] t7_add_out;
    logic [4:0] t8_idx_in;
    logic t8_idx_write_en;
    logic t8_idx_clk;
    logic [4:0] t8_idx_out;
    logic t8_idx_done;
    logic [4:0] t8_add_left;
    logic [4:0] t8_add_right;
    logic [4:0] t8_add_out;
    logic [4:0] t9_idx_in;
    logic t9_idx_write_en;
    logic t9_idx_clk;
    logic [4:0] t9_idx_out;
    logic t9_idx_done;
    logic [4:0] t9_add_left;
    logic [4:0] t9_add_right;
    logic [4:0] t9_add_out;
    logic [4:0] t10_idx_in;
    logic t10_idx_write_en;
    logic t10_idx_clk;
    logic [4:0] t10_idx_out;
    logic t10_idx_done;
    logic [4:0] t10_add_left;
    logic [4:0] t10_add_right;
    logic [4:0] t10_add_out;
    logic [4:0] t11_idx_in;
    logic t11_idx_write_en;
    logic t11_idx_clk;
    logic [4:0] t11_idx_out;
    logic t11_idx_done;
    logic [4:0] t11_add_left;
    logic [4:0] t11_add_right;
    logic [4:0] t11_add_out;
    logic [4:0] t12_idx_in;
    logic t12_idx_write_en;
    logic t12_idx_clk;
    logic [4:0] t12_idx_out;
    logic t12_idx_done;
    logic [4:0] t12_add_left;
    logic [4:0] t12_add_right;
    logic [4:0] t12_add_out;
    logic [4:0] t13_idx_in;
    logic t13_idx_write_en;
    logic t13_idx_clk;
    logic [4:0] t13_idx_out;
    logic t13_idx_done;
    logic [4:0] t13_add_left;
    logic [4:0] t13_add_right;
    logic [4:0] t13_add_out;
    logic [4:0] t14_idx_in;
    logic t14_idx_write_en;
    logic t14_idx_clk;
    logic [4:0] t14_idx_out;
    logic t14_idx_done;
    logic [4:0] t14_add_left;
    logic [4:0] t14_add_right;
    logic [4:0] t14_add_out;
    logic [4:0] t15_idx_in;
    logic t15_idx_write_en;
    logic t15_idx_clk;
    logic [4:0] t15_idx_out;
    logic t15_idx_done;
    logic [4:0] t15_add_left;
    logic [4:0] t15_add_right;
    logic [4:0] t15_add_out;
    logic [4:0] l0_idx_in;
    logic l0_idx_write_en;
    logic l0_idx_clk;
    logic [4:0] l0_idx_out;
    logic l0_idx_done;
    logic [4:0] l0_add_left;
    logic [4:0] l0_add_right;
    logic [4:0] l0_add_out;
    logic [4:0] l1_idx_in;
    logic l1_idx_write_en;
    logic l1_idx_clk;
    logic [4:0] l1_idx_out;
    logic l1_idx_done;
    logic [4:0] l1_add_left;
    logic [4:0] l1_add_right;
    logic [4:0] l1_add_out;
    logic [4:0] l2_idx_in;
    logic l2_idx_write_en;
    logic l2_idx_clk;
    logic [4:0] l2_idx_out;
    logic l2_idx_done;
    logic [4:0] l2_add_left;
    logic [4:0] l2_add_right;
    logic [4:0] l2_add_out;
    logic [4:0] l3_idx_in;
    logic l3_idx_write_en;
    logic l3_idx_clk;
    logic [4:0] l3_idx_out;
    logic l3_idx_done;
    logic [4:0] l3_add_left;
    logic [4:0] l3_add_right;
    logic [4:0] l3_add_out;
    logic [4:0] l4_idx_in;
    logic l4_idx_write_en;
    logic l4_idx_clk;
    logic [4:0] l4_idx_out;
    logic l4_idx_done;
    logic [4:0] l4_add_left;
    logic [4:0] l4_add_right;
    logic [4:0] l4_add_out;
    logic [4:0] l5_idx_in;
    logic l5_idx_write_en;
    logic l5_idx_clk;
    logic [4:0] l5_idx_out;
    logic l5_idx_done;
    logic [4:0] l5_add_left;
    logic [4:0] l5_add_right;
    logic [4:0] l5_add_out;
    logic [4:0] l6_idx_in;
    logic l6_idx_write_en;
    logic l6_idx_clk;
    logic [4:0] l6_idx_out;
    logic l6_idx_done;
    logic [4:0] l6_add_left;
    logic [4:0] l6_add_right;
    logic [4:0] l6_add_out;
    logic [4:0] l7_idx_in;
    logic l7_idx_write_en;
    logic l7_idx_clk;
    logic [4:0] l7_idx_out;
    logic l7_idx_done;
    logic [4:0] l7_add_left;
    logic [4:0] l7_add_right;
    logic [4:0] l7_add_out;
    logic [4:0] l8_idx_in;
    logic l8_idx_write_en;
    logic l8_idx_clk;
    logic [4:0] l8_idx_out;
    logic l8_idx_done;
    logic [4:0] l8_add_left;
    logic [4:0] l8_add_right;
    logic [4:0] l8_add_out;
    logic [4:0] l9_idx_in;
    logic l9_idx_write_en;
    logic l9_idx_clk;
    logic [4:0] l9_idx_out;
    logic l9_idx_done;
    logic [4:0] l9_add_left;
    logic [4:0] l9_add_right;
    logic [4:0] l9_add_out;
    logic [4:0] l10_idx_in;
    logic l10_idx_write_en;
    logic l10_idx_clk;
    logic [4:0] l10_idx_out;
    logic l10_idx_done;
    logic [4:0] l10_add_left;
    logic [4:0] l10_add_right;
    logic [4:0] l10_add_out;
    logic [4:0] l11_idx_in;
    logic l11_idx_write_en;
    logic l11_idx_clk;
    logic [4:0] l11_idx_out;
    logic l11_idx_done;
    logic [4:0] l11_add_left;
    logic [4:0] l11_add_right;
    logic [4:0] l11_add_out;
    logic [4:0] l12_idx_in;
    logic l12_idx_write_en;
    logic l12_idx_clk;
    logic [4:0] l12_idx_out;
    logic l12_idx_done;
    logic [4:0] l12_add_left;
    logic [4:0] l12_add_right;
    logic [4:0] l12_add_out;
    logic [4:0] l13_idx_in;
    logic l13_idx_write_en;
    logic l13_idx_clk;
    logic [4:0] l13_idx_out;
    logic l13_idx_done;
    logic [4:0] l13_add_left;
    logic [4:0] l13_add_right;
    logic [4:0] l13_add_out;
    logic [4:0] l14_idx_in;
    logic l14_idx_write_en;
    logic l14_idx_clk;
    logic [4:0] l14_idx_out;
    logic l14_idx_done;
    logic [4:0] l14_add_left;
    logic [4:0] l14_add_right;
    logic [4:0] l14_add_out;
    logic [4:0] l15_idx_in;
    logic l15_idx_write_en;
    logic l15_idx_clk;
    logic [4:0] l15_idx_out;
    logic l15_idx_done;
    logic [4:0] l15_add_left;
    logic [4:0] l15_add_right;
    logic [4:0] l15_add_out;
    logic [31:0] pe_0_0_top;
    logic [31:0] pe_0_0_left;
    logic [31:0] pe_0_0_out;
    logic pe_0_0_go;
    logic pe_0_0_clk;
    logic pe_0_0_done;
    logic [31:0] top_0_0_in;
    logic top_0_0_write_en;
    logic top_0_0_clk;
    logic [31:0] top_0_0_out;
    logic top_0_0_done;
    logic [31:0] left_0_0_in;
    logic left_0_0_write_en;
    logic left_0_0_clk;
    logic [31:0] left_0_0_out;
    logic left_0_0_done;
    logic [31:0] pe_0_1_top;
    logic [31:0] pe_0_1_left;
    logic [31:0] pe_0_1_out;
    logic pe_0_1_go;
    logic pe_0_1_clk;
    logic pe_0_1_done;
    logic [31:0] top_0_1_in;
    logic top_0_1_write_en;
    logic top_0_1_clk;
    logic [31:0] top_0_1_out;
    logic top_0_1_done;
    logic [31:0] left_0_1_in;
    logic left_0_1_write_en;
    logic left_0_1_clk;
    logic [31:0] left_0_1_out;
    logic left_0_1_done;
    logic [31:0] pe_0_2_top;
    logic [31:0] pe_0_2_left;
    logic [31:0] pe_0_2_out;
    logic pe_0_2_go;
    logic pe_0_2_clk;
    logic pe_0_2_done;
    logic [31:0] top_0_2_in;
    logic top_0_2_write_en;
    logic top_0_2_clk;
    logic [31:0] top_0_2_out;
    logic top_0_2_done;
    logic [31:0] left_0_2_in;
    logic left_0_2_write_en;
    logic left_0_2_clk;
    logic [31:0] left_0_2_out;
    logic left_0_2_done;
    logic [31:0] pe_0_3_top;
    logic [31:0] pe_0_3_left;
    logic [31:0] pe_0_3_out;
    logic pe_0_3_go;
    logic pe_0_3_clk;
    logic pe_0_3_done;
    logic [31:0] top_0_3_in;
    logic top_0_3_write_en;
    logic top_0_3_clk;
    logic [31:0] top_0_3_out;
    logic top_0_3_done;
    logic [31:0] left_0_3_in;
    logic left_0_3_write_en;
    logic left_0_3_clk;
    logic [31:0] left_0_3_out;
    logic left_0_3_done;
    logic [31:0] pe_0_4_top;
    logic [31:0] pe_0_4_left;
    logic [31:0] pe_0_4_out;
    logic pe_0_4_go;
    logic pe_0_4_clk;
    logic pe_0_4_done;
    logic [31:0] top_0_4_in;
    logic top_0_4_write_en;
    logic top_0_4_clk;
    logic [31:0] top_0_4_out;
    logic top_0_4_done;
    logic [31:0] left_0_4_in;
    logic left_0_4_write_en;
    logic left_0_4_clk;
    logic [31:0] left_0_4_out;
    logic left_0_4_done;
    logic [31:0] pe_0_5_top;
    logic [31:0] pe_0_5_left;
    logic [31:0] pe_0_5_out;
    logic pe_0_5_go;
    logic pe_0_5_clk;
    logic pe_0_5_done;
    logic [31:0] top_0_5_in;
    logic top_0_5_write_en;
    logic top_0_5_clk;
    logic [31:0] top_0_5_out;
    logic top_0_5_done;
    logic [31:0] left_0_5_in;
    logic left_0_5_write_en;
    logic left_0_5_clk;
    logic [31:0] left_0_5_out;
    logic left_0_5_done;
    logic [31:0] pe_0_6_top;
    logic [31:0] pe_0_6_left;
    logic [31:0] pe_0_6_out;
    logic pe_0_6_go;
    logic pe_0_6_clk;
    logic pe_0_6_done;
    logic [31:0] top_0_6_in;
    logic top_0_6_write_en;
    logic top_0_6_clk;
    logic [31:0] top_0_6_out;
    logic top_0_6_done;
    logic [31:0] left_0_6_in;
    logic left_0_6_write_en;
    logic left_0_6_clk;
    logic [31:0] left_0_6_out;
    logic left_0_6_done;
    logic [31:0] pe_0_7_top;
    logic [31:0] pe_0_7_left;
    logic [31:0] pe_0_7_out;
    logic pe_0_7_go;
    logic pe_0_7_clk;
    logic pe_0_7_done;
    logic [31:0] top_0_7_in;
    logic top_0_7_write_en;
    logic top_0_7_clk;
    logic [31:0] top_0_7_out;
    logic top_0_7_done;
    logic [31:0] left_0_7_in;
    logic left_0_7_write_en;
    logic left_0_7_clk;
    logic [31:0] left_0_7_out;
    logic left_0_7_done;
    logic [31:0] pe_0_8_top;
    logic [31:0] pe_0_8_left;
    logic [31:0] pe_0_8_out;
    logic pe_0_8_go;
    logic pe_0_8_clk;
    logic pe_0_8_done;
    logic [31:0] top_0_8_in;
    logic top_0_8_write_en;
    logic top_0_8_clk;
    logic [31:0] top_0_8_out;
    logic top_0_8_done;
    logic [31:0] left_0_8_in;
    logic left_0_8_write_en;
    logic left_0_8_clk;
    logic [31:0] left_0_8_out;
    logic left_0_8_done;
    logic [31:0] pe_0_9_top;
    logic [31:0] pe_0_9_left;
    logic [31:0] pe_0_9_out;
    logic pe_0_9_go;
    logic pe_0_9_clk;
    logic pe_0_9_done;
    logic [31:0] top_0_9_in;
    logic top_0_9_write_en;
    logic top_0_9_clk;
    logic [31:0] top_0_9_out;
    logic top_0_9_done;
    logic [31:0] left_0_9_in;
    logic left_0_9_write_en;
    logic left_0_9_clk;
    logic [31:0] left_0_9_out;
    logic left_0_9_done;
    logic [31:0] pe_0_10_top;
    logic [31:0] pe_0_10_left;
    logic [31:0] pe_0_10_out;
    logic pe_0_10_go;
    logic pe_0_10_clk;
    logic pe_0_10_done;
    logic [31:0] top_0_10_in;
    logic top_0_10_write_en;
    logic top_0_10_clk;
    logic [31:0] top_0_10_out;
    logic top_0_10_done;
    logic [31:0] left_0_10_in;
    logic left_0_10_write_en;
    logic left_0_10_clk;
    logic [31:0] left_0_10_out;
    logic left_0_10_done;
    logic [31:0] pe_0_11_top;
    logic [31:0] pe_0_11_left;
    logic [31:0] pe_0_11_out;
    logic pe_0_11_go;
    logic pe_0_11_clk;
    logic pe_0_11_done;
    logic [31:0] top_0_11_in;
    logic top_0_11_write_en;
    logic top_0_11_clk;
    logic [31:0] top_0_11_out;
    logic top_0_11_done;
    logic [31:0] left_0_11_in;
    logic left_0_11_write_en;
    logic left_0_11_clk;
    logic [31:0] left_0_11_out;
    logic left_0_11_done;
    logic [31:0] pe_0_12_top;
    logic [31:0] pe_0_12_left;
    logic [31:0] pe_0_12_out;
    logic pe_0_12_go;
    logic pe_0_12_clk;
    logic pe_0_12_done;
    logic [31:0] top_0_12_in;
    logic top_0_12_write_en;
    logic top_0_12_clk;
    logic [31:0] top_0_12_out;
    logic top_0_12_done;
    logic [31:0] left_0_12_in;
    logic left_0_12_write_en;
    logic left_0_12_clk;
    logic [31:0] left_0_12_out;
    logic left_0_12_done;
    logic [31:0] pe_0_13_top;
    logic [31:0] pe_0_13_left;
    logic [31:0] pe_0_13_out;
    logic pe_0_13_go;
    logic pe_0_13_clk;
    logic pe_0_13_done;
    logic [31:0] top_0_13_in;
    logic top_0_13_write_en;
    logic top_0_13_clk;
    logic [31:0] top_0_13_out;
    logic top_0_13_done;
    logic [31:0] left_0_13_in;
    logic left_0_13_write_en;
    logic left_0_13_clk;
    logic [31:0] left_0_13_out;
    logic left_0_13_done;
    logic [31:0] pe_0_14_top;
    logic [31:0] pe_0_14_left;
    logic [31:0] pe_0_14_out;
    logic pe_0_14_go;
    logic pe_0_14_clk;
    logic pe_0_14_done;
    logic [31:0] top_0_14_in;
    logic top_0_14_write_en;
    logic top_0_14_clk;
    logic [31:0] top_0_14_out;
    logic top_0_14_done;
    logic [31:0] left_0_14_in;
    logic left_0_14_write_en;
    logic left_0_14_clk;
    logic [31:0] left_0_14_out;
    logic left_0_14_done;
    logic [31:0] pe_0_15_top;
    logic [31:0] pe_0_15_left;
    logic [31:0] pe_0_15_out;
    logic pe_0_15_go;
    logic pe_0_15_clk;
    logic pe_0_15_done;
    logic [31:0] top_0_15_in;
    logic top_0_15_write_en;
    logic top_0_15_clk;
    logic [31:0] top_0_15_out;
    logic top_0_15_done;
    logic [31:0] left_0_15_in;
    logic left_0_15_write_en;
    logic left_0_15_clk;
    logic [31:0] left_0_15_out;
    logic left_0_15_done;
    logic [31:0] pe_1_0_top;
    logic [31:0] pe_1_0_left;
    logic [31:0] pe_1_0_out;
    logic pe_1_0_go;
    logic pe_1_0_clk;
    logic pe_1_0_done;
    logic [31:0] top_1_0_in;
    logic top_1_0_write_en;
    logic top_1_0_clk;
    logic [31:0] top_1_0_out;
    logic top_1_0_done;
    logic [31:0] left_1_0_in;
    logic left_1_0_write_en;
    logic left_1_0_clk;
    logic [31:0] left_1_0_out;
    logic left_1_0_done;
    logic [31:0] pe_1_1_top;
    logic [31:0] pe_1_1_left;
    logic [31:0] pe_1_1_out;
    logic pe_1_1_go;
    logic pe_1_1_clk;
    logic pe_1_1_done;
    logic [31:0] top_1_1_in;
    logic top_1_1_write_en;
    logic top_1_1_clk;
    logic [31:0] top_1_1_out;
    logic top_1_1_done;
    logic [31:0] left_1_1_in;
    logic left_1_1_write_en;
    logic left_1_1_clk;
    logic [31:0] left_1_1_out;
    logic left_1_1_done;
    logic [31:0] pe_1_2_top;
    logic [31:0] pe_1_2_left;
    logic [31:0] pe_1_2_out;
    logic pe_1_2_go;
    logic pe_1_2_clk;
    logic pe_1_2_done;
    logic [31:0] top_1_2_in;
    logic top_1_2_write_en;
    logic top_1_2_clk;
    logic [31:0] top_1_2_out;
    logic top_1_2_done;
    logic [31:0] left_1_2_in;
    logic left_1_2_write_en;
    logic left_1_2_clk;
    logic [31:0] left_1_2_out;
    logic left_1_2_done;
    logic [31:0] pe_1_3_top;
    logic [31:0] pe_1_3_left;
    logic [31:0] pe_1_3_out;
    logic pe_1_3_go;
    logic pe_1_3_clk;
    logic pe_1_3_done;
    logic [31:0] top_1_3_in;
    logic top_1_3_write_en;
    logic top_1_3_clk;
    logic [31:0] top_1_3_out;
    logic top_1_3_done;
    logic [31:0] left_1_3_in;
    logic left_1_3_write_en;
    logic left_1_3_clk;
    logic [31:0] left_1_3_out;
    logic left_1_3_done;
    logic [31:0] pe_1_4_top;
    logic [31:0] pe_1_4_left;
    logic [31:0] pe_1_4_out;
    logic pe_1_4_go;
    logic pe_1_4_clk;
    logic pe_1_4_done;
    logic [31:0] top_1_4_in;
    logic top_1_4_write_en;
    logic top_1_4_clk;
    logic [31:0] top_1_4_out;
    logic top_1_4_done;
    logic [31:0] left_1_4_in;
    logic left_1_4_write_en;
    logic left_1_4_clk;
    logic [31:0] left_1_4_out;
    logic left_1_4_done;
    logic [31:0] pe_1_5_top;
    logic [31:0] pe_1_5_left;
    logic [31:0] pe_1_5_out;
    logic pe_1_5_go;
    logic pe_1_5_clk;
    logic pe_1_5_done;
    logic [31:0] top_1_5_in;
    logic top_1_5_write_en;
    logic top_1_5_clk;
    logic [31:0] top_1_5_out;
    logic top_1_5_done;
    logic [31:0] left_1_5_in;
    logic left_1_5_write_en;
    logic left_1_5_clk;
    logic [31:0] left_1_5_out;
    logic left_1_5_done;
    logic [31:0] pe_1_6_top;
    logic [31:0] pe_1_6_left;
    logic [31:0] pe_1_6_out;
    logic pe_1_6_go;
    logic pe_1_6_clk;
    logic pe_1_6_done;
    logic [31:0] top_1_6_in;
    logic top_1_6_write_en;
    logic top_1_6_clk;
    logic [31:0] top_1_6_out;
    logic top_1_6_done;
    logic [31:0] left_1_6_in;
    logic left_1_6_write_en;
    logic left_1_6_clk;
    logic [31:0] left_1_6_out;
    logic left_1_6_done;
    logic [31:0] pe_1_7_top;
    logic [31:0] pe_1_7_left;
    logic [31:0] pe_1_7_out;
    logic pe_1_7_go;
    logic pe_1_7_clk;
    logic pe_1_7_done;
    logic [31:0] top_1_7_in;
    logic top_1_7_write_en;
    logic top_1_7_clk;
    logic [31:0] top_1_7_out;
    logic top_1_7_done;
    logic [31:0] left_1_7_in;
    logic left_1_7_write_en;
    logic left_1_7_clk;
    logic [31:0] left_1_7_out;
    logic left_1_7_done;
    logic [31:0] pe_1_8_top;
    logic [31:0] pe_1_8_left;
    logic [31:0] pe_1_8_out;
    logic pe_1_8_go;
    logic pe_1_8_clk;
    logic pe_1_8_done;
    logic [31:0] top_1_8_in;
    logic top_1_8_write_en;
    logic top_1_8_clk;
    logic [31:0] top_1_8_out;
    logic top_1_8_done;
    logic [31:0] left_1_8_in;
    logic left_1_8_write_en;
    logic left_1_8_clk;
    logic [31:0] left_1_8_out;
    logic left_1_8_done;
    logic [31:0] pe_1_9_top;
    logic [31:0] pe_1_9_left;
    logic [31:0] pe_1_9_out;
    logic pe_1_9_go;
    logic pe_1_9_clk;
    logic pe_1_9_done;
    logic [31:0] top_1_9_in;
    logic top_1_9_write_en;
    logic top_1_9_clk;
    logic [31:0] top_1_9_out;
    logic top_1_9_done;
    logic [31:0] left_1_9_in;
    logic left_1_9_write_en;
    logic left_1_9_clk;
    logic [31:0] left_1_9_out;
    logic left_1_9_done;
    logic [31:0] pe_1_10_top;
    logic [31:0] pe_1_10_left;
    logic [31:0] pe_1_10_out;
    logic pe_1_10_go;
    logic pe_1_10_clk;
    logic pe_1_10_done;
    logic [31:0] top_1_10_in;
    logic top_1_10_write_en;
    logic top_1_10_clk;
    logic [31:0] top_1_10_out;
    logic top_1_10_done;
    logic [31:0] left_1_10_in;
    logic left_1_10_write_en;
    logic left_1_10_clk;
    logic [31:0] left_1_10_out;
    logic left_1_10_done;
    logic [31:0] pe_1_11_top;
    logic [31:0] pe_1_11_left;
    logic [31:0] pe_1_11_out;
    logic pe_1_11_go;
    logic pe_1_11_clk;
    logic pe_1_11_done;
    logic [31:0] top_1_11_in;
    logic top_1_11_write_en;
    logic top_1_11_clk;
    logic [31:0] top_1_11_out;
    logic top_1_11_done;
    logic [31:0] left_1_11_in;
    logic left_1_11_write_en;
    logic left_1_11_clk;
    logic [31:0] left_1_11_out;
    logic left_1_11_done;
    logic [31:0] pe_1_12_top;
    logic [31:0] pe_1_12_left;
    logic [31:0] pe_1_12_out;
    logic pe_1_12_go;
    logic pe_1_12_clk;
    logic pe_1_12_done;
    logic [31:0] top_1_12_in;
    logic top_1_12_write_en;
    logic top_1_12_clk;
    logic [31:0] top_1_12_out;
    logic top_1_12_done;
    logic [31:0] left_1_12_in;
    logic left_1_12_write_en;
    logic left_1_12_clk;
    logic [31:0] left_1_12_out;
    logic left_1_12_done;
    logic [31:0] pe_1_13_top;
    logic [31:0] pe_1_13_left;
    logic [31:0] pe_1_13_out;
    logic pe_1_13_go;
    logic pe_1_13_clk;
    logic pe_1_13_done;
    logic [31:0] top_1_13_in;
    logic top_1_13_write_en;
    logic top_1_13_clk;
    logic [31:0] top_1_13_out;
    logic top_1_13_done;
    logic [31:0] left_1_13_in;
    logic left_1_13_write_en;
    logic left_1_13_clk;
    logic [31:0] left_1_13_out;
    logic left_1_13_done;
    logic [31:0] pe_1_14_top;
    logic [31:0] pe_1_14_left;
    logic [31:0] pe_1_14_out;
    logic pe_1_14_go;
    logic pe_1_14_clk;
    logic pe_1_14_done;
    logic [31:0] top_1_14_in;
    logic top_1_14_write_en;
    logic top_1_14_clk;
    logic [31:0] top_1_14_out;
    logic top_1_14_done;
    logic [31:0] left_1_14_in;
    logic left_1_14_write_en;
    logic left_1_14_clk;
    logic [31:0] left_1_14_out;
    logic left_1_14_done;
    logic [31:0] pe_1_15_top;
    logic [31:0] pe_1_15_left;
    logic [31:0] pe_1_15_out;
    logic pe_1_15_go;
    logic pe_1_15_clk;
    logic pe_1_15_done;
    logic [31:0] top_1_15_in;
    logic top_1_15_write_en;
    logic top_1_15_clk;
    logic [31:0] top_1_15_out;
    logic top_1_15_done;
    logic [31:0] left_1_15_in;
    logic left_1_15_write_en;
    logic left_1_15_clk;
    logic [31:0] left_1_15_out;
    logic left_1_15_done;
    logic [31:0] pe_2_0_top;
    logic [31:0] pe_2_0_left;
    logic [31:0] pe_2_0_out;
    logic pe_2_0_go;
    logic pe_2_0_clk;
    logic pe_2_0_done;
    logic [31:0] top_2_0_in;
    logic top_2_0_write_en;
    logic top_2_0_clk;
    logic [31:0] top_2_0_out;
    logic top_2_0_done;
    logic [31:0] left_2_0_in;
    logic left_2_0_write_en;
    logic left_2_0_clk;
    logic [31:0] left_2_0_out;
    logic left_2_0_done;
    logic [31:0] pe_2_1_top;
    logic [31:0] pe_2_1_left;
    logic [31:0] pe_2_1_out;
    logic pe_2_1_go;
    logic pe_2_1_clk;
    logic pe_2_1_done;
    logic [31:0] top_2_1_in;
    logic top_2_1_write_en;
    logic top_2_1_clk;
    logic [31:0] top_2_1_out;
    logic top_2_1_done;
    logic [31:0] left_2_1_in;
    logic left_2_1_write_en;
    logic left_2_1_clk;
    logic [31:0] left_2_1_out;
    logic left_2_1_done;
    logic [31:0] pe_2_2_top;
    logic [31:0] pe_2_2_left;
    logic [31:0] pe_2_2_out;
    logic pe_2_2_go;
    logic pe_2_2_clk;
    logic pe_2_2_done;
    logic [31:0] top_2_2_in;
    logic top_2_2_write_en;
    logic top_2_2_clk;
    logic [31:0] top_2_2_out;
    logic top_2_2_done;
    logic [31:0] left_2_2_in;
    logic left_2_2_write_en;
    logic left_2_2_clk;
    logic [31:0] left_2_2_out;
    logic left_2_2_done;
    logic [31:0] pe_2_3_top;
    logic [31:0] pe_2_3_left;
    logic [31:0] pe_2_3_out;
    logic pe_2_3_go;
    logic pe_2_3_clk;
    logic pe_2_3_done;
    logic [31:0] top_2_3_in;
    logic top_2_3_write_en;
    logic top_2_3_clk;
    logic [31:0] top_2_3_out;
    logic top_2_3_done;
    logic [31:0] left_2_3_in;
    logic left_2_3_write_en;
    logic left_2_3_clk;
    logic [31:0] left_2_3_out;
    logic left_2_3_done;
    logic [31:0] pe_2_4_top;
    logic [31:0] pe_2_4_left;
    logic [31:0] pe_2_4_out;
    logic pe_2_4_go;
    logic pe_2_4_clk;
    logic pe_2_4_done;
    logic [31:0] top_2_4_in;
    logic top_2_4_write_en;
    logic top_2_4_clk;
    logic [31:0] top_2_4_out;
    logic top_2_4_done;
    logic [31:0] left_2_4_in;
    logic left_2_4_write_en;
    logic left_2_4_clk;
    logic [31:0] left_2_4_out;
    logic left_2_4_done;
    logic [31:0] pe_2_5_top;
    logic [31:0] pe_2_5_left;
    logic [31:0] pe_2_5_out;
    logic pe_2_5_go;
    logic pe_2_5_clk;
    logic pe_2_5_done;
    logic [31:0] top_2_5_in;
    logic top_2_5_write_en;
    logic top_2_5_clk;
    logic [31:0] top_2_5_out;
    logic top_2_5_done;
    logic [31:0] left_2_5_in;
    logic left_2_5_write_en;
    logic left_2_5_clk;
    logic [31:0] left_2_5_out;
    logic left_2_5_done;
    logic [31:0] pe_2_6_top;
    logic [31:0] pe_2_6_left;
    logic [31:0] pe_2_6_out;
    logic pe_2_6_go;
    logic pe_2_6_clk;
    logic pe_2_6_done;
    logic [31:0] top_2_6_in;
    logic top_2_6_write_en;
    logic top_2_6_clk;
    logic [31:0] top_2_6_out;
    logic top_2_6_done;
    logic [31:0] left_2_6_in;
    logic left_2_6_write_en;
    logic left_2_6_clk;
    logic [31:0] left_2_6_out;
    logic left_2_6_done;
    logic [31:0] pe_2_7_top;
    logic [31:0] pe_2_7_left;
    logic [31:0] pe_2_7_out;
    logic pe_2_7_go;
    logic pe_2_7_clk;
    logic pe_2_7_done;
    logic [31:0] top_2_7_in;
    logic top_2_7_write_en;
    logic top_2_7_clk;
    logic [31:0] top_2_7_out;
    logic top_2_7_done;
    logic [31:0] left_2_7_in;
    logic left_2_7_write_en;
    logic left_2_7_clk;
    logic [31:0] left_2_7_out;
    logic left_2_7_done;
    logic [31:0] pe_2_8_top;
    logic [31:0] pe_2_8_left;
    logic [31:0] pe_2_8_out;
    logic pe_2_8_go;
    logic pe_2_8_clk;
    logic pe_2_8_done;
    logic [31:0] top_2_8_in;
    logic top_2_8_write_en;
    logic top_2_8_clk;
    logic [31:0] top_2_8_out;
    logic top_2_8_done;
    logic [31:0] left_2_8_in;
    logic left_2_8_write_en;
    logic left_2_8_clk;
    logic [31:0] left_2_8_out;
    logic left_2_8_done;
    logic [31:0] pe_2_9_top;
    logic [31:0] pe_2_9_left;
    logic [31:0] pe_2_9_out;
    logic pe_2_9_go;
    logic pe_2_9_clk;
    logic pe_2_9_done;
    logic [31:0] top_2_9_in;
    logic top_2_9_write_en;
    logic top_2_9_clk;
    logic [31:0] top_2_9_out;
    logic top_2_9_done;
    logic [31:0] left_2_9_in;
    logic left_2_9_write_en;
    logic left_2_9_clk;
    logic [31:0] left_2_9_out;
    logic left_2_9_done;
    logic [31:0] pe_2_10_top;
    logic [31:0] pe_2_10_left;
    logic [31:0] pe_2_10_out;
    logic pe_2_10_go;
    logic pe_2_10_clk;
    logic pe_2_10_done;
    logic [31:0] top_2_10_in;
    logic top_2_10_write_en;
    logic top_2_10_clk;
    logic [31:0] top_2_10_out;
    logic top_2_10_done;
    logic [31:0] left_2_10_in;
    logic left_2_10_write_en;
    logic left_2_10_clk;
    logic [31:0] left_2_10_out;
    logic left_2_10_done;
    logic [31:0] pe_2_11_top;
    logic [31:0] pe_2_11_left;
    logic [31:0] pe_2_11_out;
    logic pe_2_11_go;
    logic pe_2_11_clk;
    logic pe_2_11_done;
    logic [31:0] top_2_11_in;
    logic top_2_11_write_en;
    logic top_2_11_clk;
    logic [31:0] top_2_11_out;
    logic top_2_11_done;
    logic [31:0] left_2_11_in;
    logic left_2_11_write_en;
    logic left_2_11_clk;
    logic [31:0] left_2_11_out;
    logic left_2_11_done;
    logic [31:0] pe_2_12_top;
    logic [31:0] pe_2_12_left;
    logic [31:0] pe_2_12_out;
    logic pe_2_12_go;
    logic pe_2_12_clk;
    logic pe_2_12_done;
    logic [31:0] top_2_12_in;
    logic top_2_12_write_en;
    logic top_2_12_clk;
    logic [31:0] top_2_12_out;
    logic top_2_12_done;
    logic [31:0] left_2_12_in;
    logic left_2_12_write_en;
    logic left_2_12_clk;
    logic [31:0] left_2_12_out;
    logic left_2_12_done;
    logic [31:0] pe_2_13_top;
    logic [31:0] pe_2_13_left;
    logic [31:0] pe_2_13_out;
    logic pe_2_13_go;
    logic pe_2_13_clk;
    logic pe_2_13_done;
    logic [31:0] top_2_13_in;
    logic top_2_13_write_en;
    logic top_2_13_clk;
    logic [31:0] top_2_13_out;
    logic top_2_13_done;
    logic [31:0] left_2_13_in;
    logic left_2_13_write_en;
    logic left_2_13_clk;
    logic [31:0] left_2_13_out;
    logic left_2_13_done;
    logic [31:0] pe_2_14_top;
    logic [31:0] pe_2_14_left;
    logic [31:0] pe_2_14_out;
    logic pe_2_14_go;
    logic pe_2_14_clk;
    logic pe_2_14_done;
    logic [31:0] top_2_14_in;
    logic top_2_14_write_en;
    logic top_2_14_clk;
    logic [31:0] top_2_14_out;
    logic top_2_14_done;
    logic [31:0] left_2_14_in;
    logic left_2_14_write_en;
    logic left_2_14_clk;
    logic [31:0] left_2_14_out;
    logic left_2_14_done;
    logic [31:0] pe_2_15_top;
    logic [31:0] pe_2_15_left;
    logic [31:0] pe_2_15_out;
    logic pe_2_15_go;
    logic pe_2_15_clk;
    logic pe_2_15_done;
    logic [31:0] top_2_15_in;
    logic top_2_15_write_en;
    logic top_2_15_clk;
    logic [31:0] top_2_15_out;
    logic top_2_15_done;
    logic [31:0] left_2_15_in;
    logic left_2_15_write_en;
    logic left_2_15_clk;
    logic [31:0] left_2_15_out;
    logic left_2_15_done;
    logic [31:0] pe_3_0_top;
    logic [31:0] pe_3_0_left;
    logic [31:0] pe_3_0_out;
    logic pe_3_0_go;
    logic pe_3_0_clk;
    logic pe_3_0_done;
    logic [31:0] top_3_0_in;
    logic top_3_0_write_en;
    logic top_3_0_clk;
    logic [31:0] top_3_0_out;
    logic top_3_0_done;
    logic [31:0] left_3_0_in;
    logic left_3_0_write_en;
    logic left_3_0_clk;
    logic [31:0] left_3_0_out;
    logic left_3_0_done;
    logic [31:0] pe_3_1_top;
    logic [31:0] pe_3_1_left;
    logic [31:0] pe_3_1_out;
    logic pe_3_1_go;
    logic pe_3_1_clk;
    logic pe_3_1_done;
    logic [31:0] top_3_1_in;
    logic top_3_1_write_en;
    logic top_3_1_clk;
    logic [31:0] top_3_1_out;
    logic top_3_1_done;
    logic [31:0] left_3_1_in;
    logic left_3_1_write_en;
    logic left_3_1_clk;
    logic [31:0] left_3_1_out;
    logic left_3_1_done;
    logic [31:0] pe_3_2_top;
    logic [31:0] pe_3_2_left;
    logic [31:0] pe_3_2_out;
    logic pe_3_2_go;
    logic pe_3_2_clk;
    logic pe_3_2_done;
    logic [31:0] top_3_2_in;
    logic top_3_2_write_en;
    logic top_3_2_clk;
    logic [31:0] top_3_2_out;
    logic top_3_2_done;
    logic [31:0] left_3_2_in;
    logic left_3_2_write_en;
    logic left_3_2_clk;
    logic [31:0] left_3_2_out;
    logic left_3_2_done;
    logic [31:0] pe_3_3_top;
    logic [31:0] pe_3_3_left;
    logic [31:0] pe_3_3_out;
    logic pe_3_3_go;
    logic pe_3_3_clk;
    logic pe_3_3_done;
    logic [31:0] top_3_3_in;
    logic top_3_3_write_en;
    logic top_3_3_clk;
    logic [31:0] top_3_3_out;
    logic top_3_3_done;
    logic [31:0] left_3_3_in;
    logic left_3_3_write_en;
    logic left_3_3_clk;
    logic [31:0] left_3_3_out;
    logic left_3_3_done;
    logic [31:0] pe_3_4_top;
    logic [31:0] pe_3_4_left;
    logic [31:0] pe_3_4_out;
    logic pe_3_4_go;
    logic pe_3_4_clk;
    logic pe_3_4_done;
    logic [31:0] top_3_4_in;
    logic top_3_4_write_en;
    logic top_3_4_clk;
    logic [31:0] top_3_4_out;
    logic top_3_4_done;
    logic [31:0] left_3_4_in;
    logic left_3_4_write_en;
    logic left_3_4_clk;
    logic [31:0] left_3_4_out;
    logic left_3_4_done;
    logic [31:0] pe_3_5_top;
    logic [31:0] pe_3_5_left;
    logic [31:0] pe_3_5_out;
    logic pe_3_5_go;
    logic pe_3_5_clk;
    logic pe_3_5_done;
    logic [31:0] top_3_5_in;
    logic top_3_5_write_en;
    logic top_3_5_clk;
    logic [31:0] top_3_5_out;
    logic top_3_5_done;
    logic [31:0] left_3_5_in;
    logic left_3_5_write_en;
    logic left_3_5_clk;
    logic [31:0] left_3_5_out;
    logic left_3_5_done;
    logic [31:0] pe_3_6_top;
    logic [31:0] pe_3_6_left;
    logic [31:0] pe_3_6_out;
    logic pe_3_6_go;
    logic pe_3_6_clk;
    logic pe_3_6_done;
    logic [31:0] top_3_6_in;
    logic top_3_6_write_en;
    logic top_3_6_clk;
    logic [31:0] top_3_6_out;
    logic top_3_6_done;
    logic [31:0] left_3_6_in;
    logic left_3_6_write_en;
    logic left_3_6_clk;
    logic [31:0] left_3_6_out;
    logic left_3_6_done;
    logic [31:0] pe_3_7_top;
    logic [31:0] pe_3_7_left;
    logic [31:0] pe_3_7_out;
    logic pe_3_7_go;
    logic pe_3_7_clk;
    logic pe_3_7_done;
    logic [31:0] top_3_7_in;
    logic top_3_7_write_en;
    logic top_3_7_clk;
    logic [31:0] top_3_7_out;
    logic top_3_7_done;
    logic [31:0] left_3_7_in;
    logic left_3_7_write_en;
    logic left_3_7_clk;
    logic [31:0] left_3_7_out;
    logic left_3_7_done;
    logic [31:0] pe_3_8_top;
    logic [31:0] pe_3_8_left;
    logic [31:0] pe_3_8_out;
    logic pe_3_8_go;
    logic pe_3_8_clk;
    logic pe_3_8_done;
    logic [31:0] top_3_8_in;
    logic top_3_8_write_en;
    logic top_3_8_clk;
    logic [31:0] top_3_8_out;
    logic top_3_8_done;
    logic [31:0] left_3_8_in;
    logic left_3_8_write_en;
    logic left_3_8_clk;
    logic [31:0] left_3_8_out;
    logic left_3_8_done;
    logic [31:0] pe_3_9_top;
    logic [31:0] pe_3_9_left;
    logic [31:0] pe_3_9_out;
    logic pe_3_9_go;
    logic pe_3_9_clk;
    logic pe_3_9_done;
    logic [31:0] top_3_9_in;
    logic top_3_9_write_en;
    logic top_3_9_clk;
    logic [31:0] top_3_9_out;
    logic top_3_9_done;
    logic [31:0] left_3_9_in;
    logic left_3_9_write_en;
    logic left_3_9_clk;
    logic [31:0] left_3_9_out;
    logic left_3_9_done;
    logic [31:0] pe_3_10_top;
    logic [31:0] pe_3_10_left;
    logic [31:0] pe_3_10_out;
    logic pe_3_10_go;
    logic pe_3_10_clk;
    logic pe_3_10_done;
    logic [31:0] top_3_10_in;
    logic top_3_10_write_en;
    logic top_3_10_clk;
    logic [31:0] top_3_10_out;
    logic top_3_10_done;
    logic [31:0] left_3_10_in;
    logic left_3_10_write_en;
    logic left_3_10_clk;
    logic [31:0] left_3_10_out;
    logic left_3_10_done;
    logic [31:0] pe_3_11_top;
    logic [31:0] pe_3_11_left;
    logic [31:0] pe_3_11_out;
    logic pe_3_11_go;
    logic pe_3_11_clk;
    logic pe_3_11_done;
    logic [31:0] top_3_11_in;
    logic top_3_11_write_en;
    logic top_3_11_clk;
    logic [31:0] top_3_11_out;
    logic top_3_11_done;
    logic [31:0] left_3_11_in;
    logic left_3_11_write_en;
    logic left_3_11_clk;
    logic [31:0] left_3_11_out;
    logic left_3_11_done;
    logic [31:0] pe_3_12_top;
    logic [31:0] pe_3_12_left;
    logic [31:0] pe_3_12_out;
    logic pe_3_12_go;
    logic pe_3_12_clk;
    logic pe_3_12_done;
    logic [31:0] top_3_12_in;
    logic top_3_12_write_en;
    logic top_3_12_clk;
    logic [31:0] top_3_12_out;
    logic top_3_12_done;
    logic [31:0] left_3_12_in;
    logic left_3_12_write_en;
    logic left_3_12_clk;
    logic [31:0] left_3_12_out;
    logic left_3_12_done;
    logic [31:0] pe_3_13_top;
    logic [31:0] pe_3_13_left;
    logic [31:0] pe_3_13_out;
    logic pe_3_13_go;
    logic pe_3_13_clk;
    logic pe_3_13_done;
    logic [31:0] top_3_13_in;
    logic top_3_13_write_en;
    logic top_3_13_clk;
    logic [31:0] top_3_13_out;
    logic top_3_13_done;
    logic [31:0] left_3_13_in;
    logic left_3_13_write_en;
    logic left_3_13_clk;
    logic [31:0] left_3_13_out;
    logic left_3_13_done;
    logic [31:0] pe_3_14_top;
    logic [31:0] pe_3_14_left;
    logic [31:0] pe_3_14_out;
    logic pe_3_14_go;
    logic pe_3_14_clk;
    logic pe_3_14_done;
    logic [31:0] top_3_14_in;
    logic top_3_14_write_en;
    logic top_3_14_clk;
    logic [31:0] top_3_14_out;
    logic top_3_14_done;
    logic [31:0] left_3_14_in;
    logic left_3_14_write_en;
    logic left_3_14_clk;
    logic [31:0] left_3_14_out;
    logic left_3_14_done;
    logic [31:0] pe_3_15_top;
    logic [31:0] pe_3_15_left;
    logic [31:0] pe_3_15_out;
    logic pe_3_15_go;
    logic pe_3_15_clk;
    logic pe_3_15_done;
    logic [31:0] top_3_15_in;
    logic top_3_15_write_en;
    logic top_3_15_clk;
    logic [31:0] top_3_15_out;
    logic top_3_15_done;
    logic [31:0] left_3_15_in;
    logic left_3_15_write_en;
    logic left_3_15_clk;
    logic [31:0] left_3_15_out;
    logic left_3_15_done;
    logic [31:0] pe_4_0_top;
    logic [31:0] pe_4_0_left;
    logic [31:0] pe_4_0_out;
    logic pe_4_0_go;
    logic pe_4_0_clk;
    logic pe_4_0_done;
    logic [31:0] top_4_0_in;
    logic top_4_0_write_en;
    logic top_4_0_clk;
    logic [31:0] top_4_0_out;
    logic top_4_0_done;
    logic [31:0] left_4_0_in;
    logic left_4_0_write_en;
    logic left_4_0_clk;
    logic [31:0] left_4_0_out;
    logic left_4_0_done;
    logic [31:0] pe_4_1_top;
    logic [31:0] pe_4_1_left;
    logic [31:0] pe_4_1_out;
    logic pe_4_1_go;
    logic pe_4_1_clk;
    logic pe_4_1_done;
    logic [31:0] top_4_1_in;
    logic top_4_1_write_en;
    logic top_4_1_clk;
    logic [31:0] top_4_1_out;
    logic top_4_1_done;
    logic [31:0] left_4_1_in;
    logic left_4_1_write_en;
    logic left_4_1_clk;
    logic [31:0] left_4_1_out;
    logic left_4_1_done;
    logic [31:0] pe_4_2_top;
    logic [31:0] pe_4_2_left;
    logic [31:0] pe_4_2_out;
    logic pe_4_2_go;
    logic pe_4_2_clk;
    logic pe_4_2_done;
    logic [31:0] top_4_2_in;
    logic top_4_2_write_en;
    logic top_4_2_clk;
    logic [31:0] top_4_2_out;
    logic top_4_2_done;
    logic [31:0] left_4_2_in;
    logic left_4_2_write_en;
    logic left_4_2_clk;
    logic [31:0] left_4_2_out;
    logic left_4_2_done;
    logic [31:0] pe_4_3_top;
    logic [31:0] pe_4_3_left;
    logic [31:0] pe_4_3_out;
    logic pe_4_3_go;
    logic pe_4_3_clk;
    logic pe_4_3_done;
    logic [31:0] top_4_3_in;
    logic top_4_3_write_en;
    logic top_4_3_clk;
    logic [31:0] top_4_3_out;
    logic top_4_3_done;
    logic [31:0] left_4_3_in;
    logic left_4_3_write_en;
    logic left_4_3_clk;
    logic [31:0] left_4_3_out;
    logic left_4_3_done;
    logic [31:0] pe_4_4_top;
    logic [31:0] pe_4_4_left;
    logic [31:0] pe_4_4_out;
    logic pe_4_4_go;
    logic pe_4_4_clk;
    logic pe_4_4_done;
    logic [31:0] top_4_4_in;
    logic top_4_4_write_en;
    logic top_4_4_clk;
    logic [31:0] top_4_4_out;
    logic top_4_4_done;
    logic [31:0] left_4_4_in;
    logic left_4_4_write_en;
    logic left_4_4_clk;
    logic [31:0] left_4_4_out;
    logic left_4_4_done;
    logic [31:0] pe_4_5_top;
    logic [31:0] pe_4_5_left;
    logic [31:0] pe_4_5_out;
    logic pe_4_5_go;
    logic pe_4_5_clk;
    logic pe_4_5_done;
    logic [31:0] top_4_5_in;
    logic top_4_5_write_en;
    logic top_4_5_clk;
    logic [31:0] top_4_5_out;
    logic top_4_5_done;
    logic [31:0] left_4_5_in;
    logic left_4_5_write_en;
    logic left_4_5_clk;
    logic [31:0] left_4_5_out;
    logic left_4_5_done;
    logic [31:0] pe_4_6_top;
    logic [31:0] pe_4_6_left;
    logic [31:0] pe_4_6_out;
    logic pe_4_6_go;
    logic pe_4_6_clk;
    logic pe_4_6_done;
    logic [31:0] top_4_6_in;
    logic top_4_6_write_en;
    logic top_4_6_clk;
    logic [31:0] top_4_6_out;
    logic top_4_6_done;
    logic [31:0] left_4_6_in;
    logic left_4_6_write_en;
    logic left_4_6_clk;
    logic [31:0] left_4_6_out;
    logic left_4_6_done;
    logic [31:0] pe_4_7_top;
    logic [31:0] pe_4_7_left;
    logic [31:0] pe_4_7_out;
    logic pe_4_7_go;
    logic pe_4_7_clk;
    logic pe_4_7_done;
    logic [31:0] top_4_7_in;
    logic top_4_7_write_en;
    logic top_4_7_clk;
    logic [31:0] top_4_7_out;
    logic top_4_7_done;
    logic [31:0] left_4_7_in;
    logic left_4_7_write_en;
    logic left_4_7_clk;
    logic [31:0] left_4_7_out;
    logic left_4_7_done;
    logic [31:0] pe_4_8_top;
    logic [31:0] pe_4_8_left;
    logic [31:0] pe_4_8_out;
    logic pe_4_8_go;
    logic pe_4_8_clk;
    logic pe_4_8_done;
    logic [31:0] top_4_8_in;
    logic top_4_8_write_en;
    logic top_4_8_clk;
    logic [31:0] top_4_8_out;
    logic top_4_8_done;
    logic [31:0] left_4_8_in;
    logic left_4_8_write_en;
    logic left_4_8_clk;
    logic [31:0] left_4_8_out;
    logic left_4_8_done;
    logic [31:0] pe_4_9_top;
    logic [31:0] pe_4_9_left;
    logic [31:0] pe_4_9_out;
    logic pe_4_9_go;
    logic pe_4_9_clk;
    logic pe_4_9_done;
    logic [31:0] top_4_9_in;
    logic top_4_9_write_en;
    logic top_4_9_clk;
    logic [31:0] top_4_9_out;
    logic top_4_9_done;
    logic [31:0] left_4_9_in;
    logic left_4_9_write_en;
    logic left_4_9_clk;
    logic [31:0] left_4_9_out;
    logic left_4_9_done;
    logic [31:0] pe_4_10_top;
    logic [31:0] pe_4_10_left;
    logic [31:0] pe_4_10_out;
    logic pe_4_10_go;
    logic pe_4_10_clk;
    logic pe_4_10_done;
    logic [31:0] top_4_10_in;
    logic top_4_10_write_en;
    logic top_4_10_clk;
    logic [31:0] top_4_10_out;
    logic top_4_10_done;
    logic [31:0] left_4_10_in;
    logic left_4_10_write_en;
    logic left_4_10_clk;
    logic [31:0] left_4_10_out;
    logic left_4_10_done;
    logic [31:0] pe_4_11_top;
    logic [31:0] pe_4_11_left;
    logic [31:0] pe_4_11_out;
    logic pe_4_11_go;
    logic pe_4_11_clk;
    logic pe_4_11_done;
    logic [31:0] top_4_11_in;
    logic top_4_11_write_en;
    logic top_4_11_clk;
    logic [31:0] top_4_11_out;
    logic top_4_11_done;
    logic [31:0] left_4_11_in;
    logic left_4_11_write_en;
    logic left_4_11_clk;
    logic [31:0] left_4_11_out;
    logic left_4_11_done;
    logic [31:0] pe_4_12_top;
    logic [31:0] pe_4_12_left;
    logic [31:0] pe_4_12_out;
    logic pe_4_12_go;
    logic pe_4_12_clk;
    logic pe_4_12_done;
    logic [31:0] top_4_12_in;
    logic top_4_12_write_en;
    logic top_4_12_clk;
    logic [31:0] top_4_12_out;
    logic top_4_12_done;
    logic [31:0] left_4_12_in;
    logic left_4_12_write_en;
    logic left_4_12_clk;
    logic [31:0] left_4_12_out;
    logic left_4_12_done;
    logic [31:0] pe_4_13_top;
    logic [31:0] pe_4_13_left;
    logic [31:0] pe_4_13_out;
    logic pe_4_13_go;
    logic pe_4_13_clk;
    logic pe_4_13_done;
    logic [31:0] top_4_13_in;
    logic top_4_13_write_en;
    logic top_4_13_clk;
    logic [31:0] top_4_13_out;
    logic top_4_13_done;
    logic [31:0] left_4_13_in;
    logic left_4_13_write_en;
    logic left_4_13_clk;
    logic [31:0] left_4_13_out;
    logic left_4_13_done;
    logic [31:0] pe_4_14_top;
    logic [31:0] pe_4_14_left;
    logic [31:0] pe_4_14_out;
    logic pe_4_14_go;
    logic pe_4_14_clk;
    logic pe_4_14_done;
    logic [31:0] top_4_14_in;
    logic top_4_14_write_en;
    logic top_4_14_clk;
    logic [31:0] top_4_14_out;
    logic top_4_14_done;
    logic [31:0] left_4_14_in;
    logic left_4_14_write_en;
    logic left_4_14_clk;
    logic [31:0] left_4_14_out;
    logic left_4_14_done;
    logic [31:0] pe_4_15_top;
    logic [31:0] pe_4_15_left;
    logic [31:0] pe_4_15_out;
    logic pe_4_15_go;
    logic pe_4_15_clk;
    logic pe_4_15_done;
    logic [31:0] top_4_15_in;
    logic top_4_15_write_en;
    logic top_4_15_clk;
    logic [31:0] top_4_15_out;
    logic top_4_15_done;
    logic [31:0] left_4_15_in;
    logic left_4_15_write_en;
    logic left_4_15_clk;
    logic [31:0] left_4_15_out;
    logic left_4_15_done;
    logic [31:0] pe_5_0_top;
    logic [31:0] pe_5_0_left;
    logic [31:0] pe_5_0_out;
    logic pe_5_0_go;
    logic pe_5_0_clk;
    logic pe_5_0_done;
    logic [31:0] top_5_0_in;
    logic top_5_0_write_en;
    logic top_5_0_clk;
    logic [31:0] top_5_0_out;
    logic top_5_0_done;
    logic [31:0] left_5_0_in;
    logic left_5_0_write_en;
    logic left_5_0_clk;
    logic [31:0] left_5_0_out;
    logic left_5_0_done;
    logic [31:0] pe_5_1_top;
    logic [31:0] pe_5_1_left;
    logic [31:0] pe_5_1_out;
    logic pe_5_1_go;
    logic pe_5_1_clk;
    logic pe_5_1_done;
    logic [31:0] top_5_1_in;
    logic top_5_1_write_en;
    logic top_5_1_clk;
    logic [31:0] top_5_1_out;
    logic top_5_1_done;
    logic [31:0] left_5_1_in;
    logic left_5_1_write_en;
    logic left_5_1_clk;
    logic [31:0] left_5_1_out;
    logic left_5_1_done;
    logic [31:0] pe_5_2_top;
    logic [31:0] pe_5_2_left;
    logic [31:0] pe_5_2_out;
    logic pe_5_2_go;
    logic pe_5_2_clk;
    logic pe_5_2_done;
    logic [31:0] top_5_2_in;
    logic top_5_2_write_en;
    logic top_5_2_clk;
    logic [31:0] top_5_2_out;
    logic top_5_2_done;
    logic [31:0] left_5_2_in;
    logic left_5_2_write_en;
    logic left_5_2_clk;
    logic [31:0] left_5_2_out;
    logic left_5_2_done;
    logic [31:0] pe_5_3_top;
    logic [31:0] pe_5_3_left;
    logic [31:0] pe_5_3_out;
    logic pe_5_3_go;
    logic pe_5_3_clk;
    logic pe_5_3_done;
    logic [31:0] top_5_3_in;
    logic top_5_3_write_en;
    logic top_5_3_clk;
    logic [31:0] top_5_3_out;
    logic top_5_3_done;
    logic [31:0] left_5_3_in;
    logic left_5_3_write_en;
    logic left_5_3_clk;
    logic [31:0] left_5_3_out;
    logic left_5_3_done;
    logic [31:0] pe_5_4_top;
    logic [31:0] pe_5_4_left;
    logic [31:0] pe_5_4_out;
    logic pe_5_4_go;
    logic pe_5_4_clk;
    logic pe_5_4_done;
    logic [31:0] top_5_4_in;
    logic top_5_4_write_en;
    logic top_5_4_clk;
    logic [31:0] top_5_4_out;
    logic top_5_4_done;
    logic [31:0] left_5_4_in;
    logic left_5_4_write_en;
    logic left_5_4_clk;
    logic [31:0] left_5_4_out;
    logic left_5_4_done;
    logic [31:0] pe_5_5_top;
    logic [31:0] pe_5_5_left;
    logic [31:0] pe_5_5_out;
    logic pe_5_5_go;
    logic pe_5_5_clk;
    logic pe_5_5_done;
    logic [31:0] top_5_5_in;
    logic top_5_5_write_en;
    logic top_5_5_clk;
    logic [31:0] top_5_5_out;
    logic top_5_5_done;
    logic [31:0] left_5_5_in;
    logic left_5_5_write_en;
    logic left_5_5_clk;
    logic [31:0] left_5_5_out;
    logic left_5_5_done;
    logic [31:0] pe_5_6_top;
    logic [31:0] pe_5_6_left;
    logic [31:0] pe_5_6_out;
    logic pe_5_6_go;
    logic pe_5_6_clk;
    logic pe_5_6_done;
    logic [31:0] top_5_6_in;
    logic top_5_6_write_en;
    logic top_5_6_clk;
    logic [31:0] top_5_6_out;
    logic top_5_6_done;
    logic [31:0] left_5_6_in;
    logic left_5_6_write_en;
    logic left_5_6_clk;
    logic [31:0] left_5_6_out;
    logic left_5_6_done;
    logic [31:0] pe_5_7_top;
    logic [31:0] pe_5_7_left;
    logic [31:0] pe_5_7_out;
    logic pe_5_7_go;
    logic pe_5_7_clk;
    logic pe_5_7_done;
    logic [31:0] top_5_7_in;
    logic top_5_7_write_en;
    logic top_5_7_clk;
    logic [31:0] top_5_7_out;
    logic top_5_7_done;
    logic [31:0] left_5_7_in;
    logic left_5_7_write_en;
    logic left_5_7_clk;
    logic [31:0] left_5_7_out;
    logic left_5_7_done;
    logic [31:0] pe_5_8_top;
    logic [31:0] pe_5_8_left;
    logic [31:0] pe_5_8_out;
    logic pe_5_8_go;
    logic pe_5_8_clk;
    logic pe_5_8_done;
    logic [31:0] top_5_8_in;
    logic top_5_8_write_en;
    logic top_5_8_clk;
    logic [31:0] top_5_8_out;
    logic top_5_8_done;
    logic [31:0] left_5_8_in;
    logic left_5_8_write_en;
    logic left_5_8_clk;
    logic [31:0] left_5_8_out;
    logic left_5_8_done;
    logic [31:0] pe_5_9_top;
    logic [31:0] pe_5_9_left;
    logic [31:0] pe_5_9_out;
    logic pe_5_9_go;
    logic pe_5_9_clk;
    logic pe_5_9_done;
    logic [31:0] top_5_9_in;
    logic top_5_9_write_en;
    logic top_5_9_clk;
    logic [31:0] top_5_9_out;
    logic top_5_9_done;
    logic [31:0] left_5_9_in;
    logic left_5_9_write_en;
    logic left_5_9_clk;
    logic [31:0] left_5_9_out;
    logic left_5_9_done;
    logic [31:0] pe_5_10_top;
    logic [31:0] pe_5_10_left;
    logic [31:0] pe_5_10_out;
    logic pe_5_10_go;
    logic pe_5_10_clk;
    logic pe_5_10_done;
    logic [31:0] top_5_10_in;
    logic top_5_10_write_en;
    logic top_5_10_clk;
    logic [31:0] top_5_10_out;
    logic top_5_10_done;
    logic [31:0] left_5_10_in;
    logic left_5_10_write_en;
    logic left_5_10_clk;
    logic [31:0] left_5_10_out;
    logic left_5_10_done;
    logic [31:0] pe_5_11_top;
    logic [31:0] pe_5_11_left;
    logic [31:0] pe_5_11_out;
    logic pe_5_11_go;
    logic pe_5_11_clk;
    logic pe_5_11_done;
    logic [31:0] top_5_11_in;
    logic top_5_11_write_en;
    logic top_5_11_clk;
    logic [31:0] top_5_11_out;
    logic top_5_11_done;
    logic [31:0] left_5_11_in;
    logic left_5_11_write_en;
    logic left_5_11_clk;
    logic [31:0] left_5_11_out;
    logic left_5_11_done;
    logic [31:0] pe_5_12_top;
    logic [31:0] pe_5_12_left;
    logic [31:0] pe_5_12_out;
    logic pe_5_12_go;
    logic pe_5_12_clk;
    logic pe_5_12_done;
    logic [31:0] top_5_12_in;
    logic top_5_12_write_en;
    logic top_5_12_clk;
    logic [31:0] top_5_12_out;
    logic top_5_12_done;
    logic [31:0] left_5_12_in;
    logic left_5_12_write_en;
    logic left_5_12_clk;
    logic [31:0] left_5_12_out;
    logic left_5_12_done;
    logic [31:0] pe_5_13_top;
    logic [31:0] pe_5_13_left;
    logic [31:0] pe_5_13_out;
    logic pe_5_13_go;
    logic pe_5_13_clk;
    logic pe_5_13_done;
    logic [31:0] top_5_13_in;
    logic top_5_13_write_en;
    logic top_5_13_clk;
    logic [31:0] top_5_13_out;
    logic top_5_13_done;
    logic [31:0] left_5_13_in;
    logic left_5_13_write_en;
    logic left_5_13_clk;
    logic [31:0] left_5_13_out;
    logic left_5_13_done;
    logic [31:0] pe_5_14_top;
    logic [31:0] pe_5_14_left;
    logic [31:0] pe_5_14_out;
    logic pe_5_14_go;
    logic pe_5_14_clk;
    logic pe_5_14_done;
    logic [31:0] top_5_14_in;
    logic top_5_14_write_en;
    logic top_5_14_clk;
    logic [31:0] top_5_14_out;
    logic top_5_14_done;
    logic [31:0] left_5_14_in;
    logic left_5_14_write_en;
    logic left_5_14_clk;
    logic [31:0] left_5_14_out;
    logic left_5_14_done;
    logic [31:0] pe_5_15_top;
    logic [31:0] pe_5_15_left;
    logic [31:0] pe_5_15_out;
    logic pe_5_15_go;
    logic pe_5_15_clk;
    logic pe_5_15_done;
    logic [31:0] top_5_15_in;
    logic top_5_15_write_en;
    logic top_5_15_clk;
    logic [31:0] top_5_15_out;
    logic top_5_15_done;
    logic [31:0] left_5_15_in;
    logic left_5_15_write_en;
    logic left_5_15_clk;
    logic [31:0] left_5_15_out;
    logic left_5_15_done;
    logic [31:0] pe_6_0_top;
    logic [31:0] pe_6_0_left;
    logic [31:0] pe_6_0_out;
    logic pe_6_0_go;
    logic pe_6_0_clk;
    logic pe_6_0_done;
    logic [31:0] top_6_0_in;
    logic top_6_0_write_en;
    logic top_6_0_clk;
    logic [31:0] top_6_0_out;
    logic top_6_0_done;
    logic [31:0] left_6_0_in;
    logic left_6_0_write_en;
    logic left_6_0_clk;
    logic [31:0] left_6_0_out;
    logic left_6_0_done;
    logic [31:0] pe_6_1_top;
    logic [31:0] pe_6_1_left;
    logic [31:0] pe_6_1_out;
    logic pe_6_1_go;
    logic pe_6_1_clk;
    logic pe_6_1_done;
    logic [31:0] top_6_1_in;
    logic top_6_1_write_en;
    logic top_6_1_clk;
    logic [31:0] top_6_1_out;
    logic top_6_1_done;
    logic [31:0] left_6_1_in;
    logic left_6_1_write_en;
    logic left_6_1_clk;
    logic [31:0] left_6_1_out;
    logic left_6_1_done;
    logic [31:0] pe_6_2_top;
    logic [31:0] pe_6_2_left;
    logic [31:0] pe_6_2_out;
    logic pe_6_2_go;
    logic pe_6_2_clk;
    logic pe_6_2_done;
    logic [31:0] top_6_2_in;
    logic top_6_2_write_en;
    logic top_6_2_clk;
    logic [31:0] top_6_2_out;
    logic top_6_2_done;
    logic [31:0] left_6_2_in;
    logic left_6_2_write_en;
    logic left_6_2_clk;
    logic [31:0] left_6_2_out;
    logic left_6_2_done;
    logic [31:0] pe_6_3_top;
    logic [31:0] pe_6_3_left;
    logic [31:0] pe_6_3_out;
    logic pe_6_3_go;
    logic pe_6_3_clk;
    logic pe_6_3_done;
    logic [31:0] top_6_3_in;
    logic top_6_3_write_en;
    logic top_6_3_clk;
    logic [31:0] top_6_3_out;
    logic top_6_3_done;
    logic [31:0] left_6_3_in;
    logic left_6_3_write_en;
    logic left_6_3_clk;
    logic [31:0] left_6_3_out;
    logic left_6_3_done;
    logic [31:0] pe_6_4_top;
    logic [31:0] pe_6_4_left;
    logic [31:0] pe_6_4_out;
    logic pe_6_4_go;
    logic pe_6_4_clk;
    logic pe_6_4_done;
    logic [31:0] top_6_4_in;
    logic top_6_4_write_en;
    logic top_6_4_clk;
    logic [31:0] top_6_4_out;
    logic top_6_4_done;
    logic [31:0] left_6_4_in;
    logic left_6_4_write_en;
    logic left_6_4_clk;
    logic [31:0] left_6_4_out;
    logic left_6_4_done;
    logic [31:0] pe_6_5_top;
    logic [31:0] pe_6_5_left;
    logic [31:0] pe_6_5_out;
    logic pe_6_5_go;
    logic pe_6_5_clk;
    logic pe_6_5_done;
    logic [31:0] top_6_5_in;
    logic top_6_5_write_en;
    logic top_6_5_clk;
    logic [31:0] top_6_5_out;
    logic top_6_5_done;
    logic [31:0] left_6_5_in;
    logic left_6_5_write_en;
    logic left_6_5_clk;
    logic [31:0] left_6_5_out;
    logic left_6_5_done;
    logic [31:0] pe_6_6_top;
    logic [31:0] pe_6_6_left;
    logic [31:0] pe_6_6_out;
    logic pe_6_6_go;
    logic pe_6_6_clk;
    logic pe_6_6_done;
    logic [31:0] top_6_6_in;
    logic top_6_6_write_en;
    logic top_6_6_clk;
    logic [31:0] top_6_6_out;
    logic top_6_6_done;
    logic [31:0] left_6_6_in;
    logic left_6_6_write_en;
    logic left_6_6_clk;
    logic [31:0] left_6_6_out;
    logic left_6_6_done;
    logic [31:0] pe_6_7_top;
    logic [31:0] pe_6_7_left;
    logic [31:0] pe_6_7_out;
    logic pe_6_7_go;
    logic pe_6_7_clk;
    logic pe_6_7_done;
    logic [31:0] top_6_7_in;
    logic top_6_7_write_en;
    logic top_6_7_clk;
    logic [31:0] top_6_7_out;
    logic top_6_7_done;
    logic [31:0] left_6_7_in;
    logic left_6_7_write_en;
    logic left_6_7_clk;
    logic [31:0] left_6_7_out;
    logic left_6_7_done;
    logic [31:0] pe_6_8_top;
    logic [31:0] pe_6_8_left;
    logic [31:0] pe_6_8_out;
    logic pe_6_8_go;
    logic pe_6_8_clk;
    logic pe_6_8_done;
    logic [31:0] top_6_8_in;
    logic top_6_8_write_en;
    logic top_6_8_clk;
    logic [31:0] top_6_8_out;
    logic top_6_8_done;
    logic [31:0] left_6_8_in;
    logic left_6_8_write_en;
    logic left_6_8_clk;
    logic [31:0] left_6_8_out;
    logic left_6_8_done;
    logic [31:0] pe_6_9_top;
    logic [31:0] pe_6_9_left;
    logic [31:0] pe_6_9_out;
    logic pe_6_9_go;
    logic pe_6_9_clk;
    logic pe_6_9_done;
    logic [31:0] top_6_9_in;
    logic top_6_9_write_en;
    logic top_6_9_clk;
    logic [31:0] top_6_9_out;
    logic top_6_9_done;
    logic [31:0] left_6_9_in;
    logic left_6_9_write_en;
    logic left_6_9_clk;
    logic [31:0] left_6_9_out;
    logic left_6_9_done;
    logic [31:0] pe_6_10_top;
    logic [31:0] pe_6_10_left;
    logic [31:0] pe_6_10_out;
    logic pe_6_10_go;
    logic pe_6_10_clk;
    logic pe_6_10_done;
    logic [31:0] top_6_10_in;
    logic top_6_10_write_en;
    logic top_6_10_clk;
    logic [31:0] top_6_10_out;
    logic top_6_10_done;
    logic [31:0] left_6_10_in;
    logic left_6_10_write_en;
    logic left_6_10_clk;
    logic [31:0] left_6_10_out;
    logic left_6_10_done;
    logic [31:0] pe_6_11_top;
    logic [31:0] pe_6_11_left;
    logic [31:0] pe_6_11_out;
    logic pe_6_11_go;
    logic pe_6_11_clk;
    logic pe_6_11_done;
    logic [31:0] top_6_11_in;
    logic top_6_11_write_en;
    logic top_6_11_clk;
    logic [31:0] top_6_11_out;
    logic top_6_11_done;
    logic [31:0] left_6_11_in;
    logic left_6_11_write_en;
    logic left_6_11_clk;
    logic [31:0] left_6_11_out;
    logic left_6_11_done;
    logic [31:0] pe_6_12_top;
    logic [31:0] pe_6_12_left;
    logic [31:0] pe_6_12_out;
    logic pe_6_12_go;
    logic pe_6_12_clk;
    logic pe_6_12_done;
    logic [31:0] top_6_12_in;
    logic top_6_12_write_en;
    logic top_6_12_clk;
    logic [31:0] top_6_12_out;
    logic top_6_12_done;
    logic [31:0] left_6_12_in;
    logic left_6_12_write_en;
    logic left_6_12_clk;
    logic [31:0] left_6_12_out;
    logic left_6_12_done;
    logic [31:0] pe_6_13_top;
    logic [31:0] pe_6_13_left;
    logic [31:0] pe_6_13_out;
    logic pe_6_13_go;
    logic pe_6_13_clk;
    logic pe_6_13_done;
    logic [31:0] top_6_13_in;
    logic top_6_13_write_en;
    logic top_6_13_clk;
    logic [31:0] top_6_13_out;
    logic top_6_13_done;
    logic [31:0] left_6_13_in;
    logic left_6_13_write_en;
    logic left_6_13_clk;
    logic [31:0] left_6_13_out;
    logic left_6_13_done;
    logic [31:0] pe_6_14_top;
    logic [31:0] pe_6_14_left;
    logic [31:0] pe_6_14_out;
    logic pe_6_14_go;
    logic pe_6_14_clk;
    logic pe_6_14_done;
    logic [31:0] top_6_14_in;
    logic top_6_14_write_en;
    logic top_6_14_clk;
    logic [31:0] top_6_14_out;
    logic top_6_14_done;
    logic [31:0] left_6_14_in;
    logic left_6_14_write_en;
    logic left_6_14_clk;
    logic [31:0] left_6_14_out;
    logic left_6_14_done;
    logic [31:0] pe_6_15_top;
    logic [31:0] pe_6_15_left;
    logic [31:0] pe_6_15_out;
    logic pe_6_15_go;
    logic pe_6_15_clk;
    logic pe_6_15_done;
    logic [31:0] top_6_15_in;
    logic top_6_15_write_en;
    logic top_6_15_clk;
    logic [31:0] top_6_15_out;
    logic top_6_15_done;
    logic [31:0] left_6_15_in;
    logic left_6_15_write_en;
    logic left_6_15_clk;
    logic [31:0] left_6_15_out;
    logic left_6_15_done;
    logic [31:0] pe_7_0_top;
    logic [31:0] pe_7_0_left;
    logic [31:0] pe_7_0_out;
    logic pe_7_0_go;
    logic pe_7_0_clk;
    logic pe_7_0_done;
    logic [31:0] top_7_0_in;
    logic top_7_0_write_en;
    logic top_7_0_clk;
    logic [31:0] top_7_0_out;
    logic top_7_0_done;
    logic [31:0] left_7_0_in;
    logic left_7_0_write_en;
    logic left_7_0_clk;
    logic [31:0] left_7_0_out;
    logic left_7_0_done;
    logic [31:0] pe_7_1_top;
    logic [31:0] pe_7_1_left;
    logic [31:0] pe_7_1_out;
    logic pe_7_1_go;
    logic pe_7_1_clk;
    logic pe_7_1_done;
    logic [31:0] top_7_1_in;
    logic top_7_1_write_en;
    logic top_7_1_clk;
    logic [31:0] top_7_1_out;
    logic top_7_1_done;
    logic [31:0] left_7_1_in;
    logic left_7_1_write_en;
    logic left_7_1_clk;
    logic [31:0] left_7_1_out;
    logic left_7_1_done;
    logic [31:0] pe_7_2_top;
    logic [31:0] pe_7_2_left;
    logic [31:0] pe_7_2_out;
    logic pe_7_2_go;
    logic pe_7_2_clk;
    logic pe_7_2_done;
    logic [31:0] top_7_2_in;
    logic top_7_2_write_en;
    logic top_7_2_clk;
    logic [31:0] top_7_2_out;
    logic top_7_2_done;
    logic [31:0] left_7_2_in;
    logic left_7_2_write_en;
    logic left_7_2_clk;
    logic [31:0] left_7_2_out;
    logic left_7_2_done;
    logic [31:0] pe_7_3_top;
    logic [31:0] pe_7_3_left;
    logic [31:0] pe_7_3_out;
    logic pe_7_3_go;
    logic pe_7_3_clk;
    logic pe_7_3_done;
    logic [31:0] top_7_3_in;
    logic top_7_3_write_en;
    logic top_7_3_clk;
    logic [31:0] top_7_3_out;
    logic top_7_3_done;
    logic [31:0] left_7_3_in;
    logic left_7_3_write_en;
    logic left_7_3_clk;
    logic [31:0] left_7_3_out;
    logic left_7_3_done;
    logic [31:0] pe_7_4_top;
    logic [31:0] pe_7_4_left;
    logic [31:0] pe_7_4_out;
    logic pe_7_4_go;
    logic pe_7_4_clk;
    logic pe_7_4_done;
    logic [31:0] top_7_4_in;
    logic top_7_4_write_en;
    logic top_7_4_clk;
    logic [31:0] top_7_4_out;
    logic top_7_4_done;
    logic [31:0] left_7_4_in;
    logic left_7_4_write_en;
    logic left_7_4_clk;
    logic [31:0] left_7_4_out;
    logic left_7_4_done;
    logic [31:0] pe_7_5_top;
    logic [31:0] pe_7_5_left;
    logic [31:0] pe_7_5_out;
    logic pe_7_5_go;
    logic pe_7_5_clk;
    logic pe_7_5_done;
    logic [31:0] top_7_5_in;
    logic top_7_5_write_en;
    logic top_7_5_clk;
    logic [31:0] top_7_5_out;
    logic top_7_5_done;
    logic [31:0] left_7_5_in;
    logic left_7_5_write_en;
    logic left_7_5_clk;
    logic [31:0] left_7_5_out;
    logic left_7_5_done;
    logic [31:0] pe_7_6_top;
    logic [31:0] pe_7_6_left;
    logic [31:0] pe_7_6_out;
    logic pe_7_6_go;
    logic pe_7_6_clk;
    logic pe_7_6_done;
    logic [31:0] top_7_6_in;
    logic top_7_6_write_en;
    logic top_7_6_clk;
    logic [31:0] top_7_6_out;
    logic top_7_6_done;
    logic [31:0] left_7_6_in;
    logic left_7_6_write_en;
    logic left_7_6_clk;
    logic [31:0] left_7_6_out;
    logic left_7_6_done;
    logic [31:0] pe_7_7_top;
    logic [31:0] pe_7_7_left;
    logic [31:0] pe_7_7_out;
    logic pe_7_7_go;
    logic pe_7_7_clk;
    logic pe_7_7_done;
    logic [31:0] top_7_7_in;
    logic top_7_7_write_en;
    logic top_7_7_clk;
    logic [31:0] top_7_7_out;
    logic top_7_7_done;
    logic [31:0] left_7_7_in;
    logic left_7_7_write_en;
    logic left_7_7_clk;
    logic [31:0] left_7_7_out;
    logic left_7_7_done;
    logic [31:0] pe_7_8_top;
    logic [31:0] pe_7_8_left;
    logic [31:0] pe_7_8_out;
    logic pe_7_8_go;
    logic pe_7_8_clk;
    logic pe_7_8_done;
    logic [31:0] top_7_8_in;
    logic top_7_8_write_en;
    logic top_7_8_clk;
    logic [31:0] top_7_8_out;
    logic top_7_8_done;
    logic [31:0] left_7_8_in;
    logic left_7_8_write_en;
    logic left_7_8_clk;
    logic [31:0] left_7_8_out;
    logic left_7_8_done;
    logic [31:0] pe_7_9_top;
    logic [31:0] pe_7_9_left;
    logic [31:0] pe_7_9_out;
    logic pe_7_9_go;
    logic pe_7_9_clk;
    logic pe_7_9_done;
    logic [31:0] top_7_9_in;
    logic top_7_9_write_en;
    logic top_7_9_clk;
    logic [31:0] top_7_9_out;
    logic top_7_9_done;
    logic [31:0] left_7_9_in;
    logic left_7_9_write_en;
    logic left_7_9_clk;
    logic [31:0] left_7_9_out;
    logic left_7_9_done;
    logic [31:0] pe_7_10_top;
    logic [31:0] pe_7_10_left;
    logic [31:0] pe_7_10_out;
    logic pe_7_10_go;
    logic pe_7_10_clk;
    logic pe_7_10_done;
    logic [31:0] top_7_10_in;
    logic top_7_10_write_en;
    logic top_7_10_clk;
    logic [31:0] top_7_10_out;
    logic top_7_10_done;
    logic [31:0] left_7_10_in;
    logic left_7_10_write_en;
    logic left_7_10_clk;
    logic [31:0] left_7_10_out;
    logic left_7_10_done;
    logic [31:0] pe_7_11_top;
    logic [31:0] pe_7_11_left;
    logic [31:0] pe_7_11_out;
    logic pe_7_11_go;
    logic pe_7_11_clk;
    logic pe_7_11_done;
    logic [31:0] top_7_11_in;
    logic top_7_11_write_en;
    logic top_7_11_clk;
    logic [31:0] top_7_11_out;
    logic top_7_11_done;
    logic [31:0] left_7_11_in;
    logic left_7_11_write_en;
    logic left_7_11_clk;
    logic [31:0] left_7_11_out;
    logic left_7_11_done;
    logic [31:0] pe_7_12_top;
    logic [31:0] pe_7_12_left;
    logic [31:0] pe_7_12_out;
    logic pe_7_12_go;
    logic pe_7_12_clk;
    logic pe_7_12_done;
    logic [31:0] top_7_12_in;
    logic top_7_12_write_en;
    logic top_7_12_clk;
    logic [31:0] top_7_12_out;
    logic top_7_12_done;
    logic [31:0] left_7_12_in;
    logic left_7_12_write_en;
    logic left_7_12_clk;
    logic [31:0] left_7_12_out;
    logic left_7_12_done;
    logic [31:0] pe_7_13_top;
    logic [31:0] pe_7_13_left;
    logic [31:0] pe_7_13_out;
    logic pe_7_13_go;
    logic pe_7_13_clk;
    logic pe_7_13_done;
    logic [31:0] top_7_13_in;
    logic top_7_13_write_en;
    logic top_7_13_clk;
    logic [31:0] top_7_13_out;
    logic top_7_13_done;
    logic [31:0] left_7_13_in;
    logic left_7_13_write_en;
    logic left_7_13_clk;
    logic [31:0] left_7_13_out;
    logic left_7_13_done;
    logic [31:0] pe_7_14_top;
    logic [31:0] pe_7_14_left;
    logic [31:0] pe_7_14_out;
    logic pe_7_14_go;
    logic pe_7_14_clk;
    logic pe_7_14_done;
    logic [31:0] top_7_14_in;
    logic top_7_14_write_en;
    logic top_7_14_clk;
    logic [31:0] top_7_14_out;
    logic top_7_14_done;
    logic [31:0] left_7_14_in;
    logic left_7_14_write_en;
    logic left_7_14_clk;
    logic [31:0] left_7_14_out;
    logic left_7_14_done;
    logic [31:0] pe_7_15_top;
    logic [31:0] pe_7_15_left;
    logic [31:0] pe_7_15_out;
    logic pe_7_15_go;
    logic pe_7_15_clk;
    logic pe_7_15_done;
    logic [31:0] top_7_15_in;
    logic top_7_15_write_en;
    logic top_7_15_clk;
    logic [31:0] top_7_15_out;
    logic top_7_15_done;
    logic [31:0] left_7_15_in;
    logic left_7_15_write_en;
    logic left_7_15_clk;
    logic [31:0] left_7_15_out;
    logic left_7_15_done;
    logic [31:0] pe_8_0_top;
    logic [31:0] pe_8_0_left;
    logic [31:0] pe_8_0_out;
    logic pe_8_0_go;
    logic pe_8_0_clk;
    logic pe_8_0_done;
    logic [31:0] top_8_0_in;
    logic top_8_0_write_en;
    logic top_8_0_clk;
    logic [31:0] top_8_0_out;
    logic top_8_0_done;
    logic [31:0] left_8_0_in;
    logic left_8_0_write_en;
    logic left_8_0_clk;
    logic [31:0] left_8_0_out;
    logic left_8_0_done;
    logic [31:0] pe_8_1_top;
    logic [31:0] pe_8_1_left;
    logic [31:0] pe_8_1_out;
    logic pe_8_1_go;
    logic pe_8_1_clk;
    logic pe_8_1_done;
    logic [31:0] top_8_1_in;
    logic top_8_1_write_en;
    logic top_8_1_clk;
    logic [31:0] top_8_1_out;
    logic top_8_1_done;
    logic [31:0] left_8_1_in;
    logic left_8_1_write_en;
    logic left_8_1_clk;
    logic [31:0] left_8_1_out;
    logic left_8_1_done;
    logic [31:0] pe_8_2_top;
    logic [31:0] pe_8_2_left;
    logic [31:0] pe_8_2_out;
    logic pe_8_2_go;
    logic pe_8_2_clk;
    logic pe_8_2_done;
    logic [31:0] top_8_2_in;
    logic top_8_2_write_en;
    logic top_8_2_clk;
    logic [31:0] top_8_2_out;
    logic top_8_2_done;
    logic [31:0] left_8_2_in;
    logic left_8_2_write_en;
    logic left_8_2_clk;
    logic [31:0] left_8_2_out;
    logic left_8_2_done;
    logic [31:0] pe_8_3_top;
    logic [31:0] pe_8_3_left;
    logic [31:0] pe_8_3_out;
    logic pe_8_3_go;
    logic pe_8_3_clk;
    logic pe_8_3_done;
    logic [31:0] top_8_3_in;
    logic top_8_3_write_en;
    logic top_8_3_clk;
    logic [31:0] top_8_3_out;
    logic top_8_3_done;
    logic [31:0] left_8_3_in;
    logic left_8_3_write_en;
    logic left_8_3_clk;
    logic [31:0] left_8_3_out;
    logic left_8_3_done;
    logic [31:0] pe_8_4_top;
    logic [31:0] pe_8_4_left;
    logic [31:0] pe_8_4_out;
    logic pe_8_4_go;
    logic pe_8_4_clk;
    logic pe_8_4_done;
    logic [31:0] top_8_4_in;
    logic top_8_4_write_en;
    logic top_8_4_clk;
    logic [31:0] top_8_4_out;
    logic top_8_4_done;
    logic [31:0] left_8_4_in;
    logic left_8_4_write_en;
    logic left_8_4_clk;
    logic [31:0] left_8_4_out;
    logic left_8_4_done;
    logic [31:0] pe_8_5_top;
    logic [31:0] pe_8_5_left;
    logic [31:0] pe_8_5_out;
    logic pe_8_5_go;
    logic pe_8_5_clk;
    logic pe_8_5_done;
    logic [31:0] top_8_5_in;
    logic top_8_5_write_en;
    logic top_8_5_clk;
    logic [31:0] top_8_5_out;
    logic top_8_5_done;
    logic [31:0] left_8_5_in;
    logic left_8_5_write_en;
    logic left_8_5_clk;
    logic [31:0] left_8_5_out;
    logic left_8_5_done;
    logic [31:0] pe_8_6_top;
    logic [31:0] pe_8_6_left;
    logic [31:0] pe_8_6_out;
    logic pe_8_6_go;
    logic pe_8_6_clk;
    logic pe_8_6_done;
    logic [31:0] top_8_6_in;
    logic top_8_6_write_en;
    logic top_8_6_clk;
    logic [31:0] top_8_6_out;
    logic top_8_6_done;
    logic [31:0] left_8_6_in;
    logic left_8_6_write_en;
    logic left_8_6_clk;
    logic [31:0] left_8_6_out;
    logic left_8_6_done;
    logic [31:0] pe_8_7_top;
    logic [31:0] pe_8_7_left;
    logic [31:0] pe_8_7_out;
    logic pe_8_7_go;
    logic pe_8_7_clk;
    logic pe_8_7_done;
    logic [31:0] top_8_7_in;
    logic top_8_7_write_en;
    logic top_8_7_clk;
    logic [31:0] top_8_7_out;
    logic top_8_7_done;
    logic [31:0] left_8_7_in;
    logic left_8_7_write_en;
    logic left_8_7_clk;
    logic [31:0] left_8_7_out;
    logic left_8_7_done;
    logic [31:0] pe_8_8_top;
    logic [31:0] pe_8_8_left;
    logic [31:0] pe_8_8_out;
    logic pe_8_8_go;
    logic pe_8_8_clk;
    logic pe_8_8_done;
    logic [31:0] top_8_8_in;
    logic top_8_8_write_en;
    logic top_8_8_clk;
    logic [31:0] top_8_8_out;
    logic top_8_8_done;
    logic [31:0] left_8_8_in;
    logic left_8_8_write_en;
    logic left_8_8_clk;
    logic [31:0] left_8_8_out;
    logic left_8_8_done;
    logic [31:0] pe_8_9_top;
    logic [31:0] pe_8_9_left;
    logic [31:0] pe_8_9_out;
    logic pe_8_9_go;
    logic pe_8_9_clk;
    logic pe_8_9_done;
    logic [31:0] top_8_9_in;
    logic top_8_9_write_en;
    logic top_8_9_clk;
    logic [31:0] top_8_9_out;
    logic top_8_9_done;
    logic [31:0] left_8_9_in;
    logic left_8_9_write_en;
    logic left_8_9_clk;
    logic [31:0] left_8_9_out;
    logic left_8_9_done;
    logic [31:0] pe_8_10_top;
    logic [31:0] pe_8_10_left;
    logic [31:0] pe_8_10_out;
    logic pe_8_10_go;
    logic pe_8_10_clk;
    logic pe_8_10_done;
    logic [31:0] top_8_10_in;
    logic top_8_10_write_en;
    logic top_8_10_clk;
    logic [31:0] top_8_10_out;
    logic top_8_10_done;
    logic [31:0] left_8_10_in;
    logic left_8_10_write_en;
    logic left_8_10_clk;
    logic [31:0] left_8_10_out;
    logic left_8_10_done;
    logic [31:0] pe_8_11_top;
    logic [31:0] pe_8_11_left;
    logic [31:0] pe_8_11_out;
    logic pe_8_11_go;
    logic pe_8_11_clk;
    logic pe_8_11_done;
    logic [31:0] top_8_11_in;
    logic top_8_11_write_en;
    logic top_8_11_clk;
    logic [31:0] top_8_11_out;
    logic top_8_11_done;
    logic [31:0] left_8_11_in;
    logic left_8_11_write_en;
    logic left_8_11_clk;
    logic [31:0] left_8_11_out;
    logic left_8_11_done;
    logic [31:0] pe_8_12_top;
    logic [31:0] pe_8_12_left;
    logic [31:0] pe_8_12_out;
    logic pe_8_12_go;
    logic pe_8_12_clk;
    logic pe_8_12_done;
    logic [31:0] top_8_12_in;
    logic top_8_12_write_en;
    logic top_8_12_clk;
    logic [31:0] top_8_12_out;
    logic top_8_12_done;
    logic [31:0] left_8_12_in;
    logic left_8_12_write_en;
    logic left_8_12_clk;
    logic [31:0] left_8_12_out;
    logic left_8_12_done;
    logic [31:0] pe_8_13_top;
    logic [31:0] pe_8_13_left;
    logic [31:0] pe_8_13_out;
    logic pe_8_13_go;
    logic pe_8_13_clk;
    logic pe_8_13_done;
    logic [31:0] top_8_13_in;
    logic top_8_13_write_en;
    logic top_8_13_clk;
    logic [31:0] top_8_13_out;
    logic top_8_13_done;
    logic [31:0] left_8_13_in;
    logic left_8_13_write_en;
    logic left_8_13_clk;
    logic [31:0] left_8_13_out;
    logic left_8_13_done;
    logic [31:0] pe_8_14_top;
    logic [31:0] pe_8_14_left;
    logic [31:0] pe_8_14_out;
    logic pe_8_14_go;
    logic pe_8_14_clk;
    logic pe_8_14_done;
    logic [31:0] top_8_14_in;
    logic top_8_14_write_en;
    logic top_8_14_clk;
    logic [31:0] top_8_14_out;
    logic top_8_14_done;
    logic [31:0] left_8_14_in;
    logic left_8_14_write_en;
    logic left_8_14_clk;
    logic [31:0] left_8_14_out;
    logic left_8_14_done;
    logic [31:0] pe_8_15_top;
    logic [31:0] pe_8_15_left;
    logic [31:0] pe_8_15_out;
    logic pe_8_15_go;
    logic pe_8_15_clk;
    logic pe_8_15_done;
    logic [31:0] top_8_15_in;
    logic top_8_15_write_en;
    logic top_8_15_clk;
    logic [31:0] top_8_15_out;
    logic top_8_15_done;
    logic [31:0] left_8_15_in;
    logic left_8_15_write_en;
    logic left_8_15_clk;
    logic [31:0] left_8_15_out;
    logic left_8_15_done;
    logic [31:0] pe_9_0_top;
    logic [31:0] pe_9_0_left;
    logic [31:0] pe_9_0_out;
    logic pe_9_0_go;
    logic pe_9_0_clk;
    logic pe_9_0_done;
    logic [31:0] top_9_0_in;
    logic top_9_0_write_en;
    logic top_9_0_clk;
    logic [31:0] top_9_0_out;
    logic top_9_0_done;
    logic [31:0] left_9_0_in;
    logic left_9_0_write_en;
    logic left_9_0_clk;
    logic [31:0] left_9_0_out;
    logic left_9_0_done;
    logic [31:0] pe_9_1_top;
    logic [31:0] pe_9_1_left;
    logic [31:0] pe_9_1_out;
    logic pe_9_1_go;
    logic pe_9_1_clk;
    logic pe_9_1_done;
    logic [31:0] top_9_1_in;
    logic top_9_1_write_en;
    logic top_9_1_clk;
    logic [31:0] top_9_1_out;
    logic top_9_1_done;
    logic [31:0] left_9_1_in;
    logic left_9_1_write_en;
    logic left_9_1_clk;
    logic [31:0] left_9_1_out;
    logic left_9_1_done;
    logic [31:0] pe_9_2_top;
    logic [31:0] pe_9_2_left;
    logic [31:0] pe_9_2_out;
    logic pe_9_2_go;
    logic pe_9_2_clk;
    logic pe_9_2_done;
    logic [31:0] top_9_2_in;
    logic top_9_2_write_en;
    logic top_9_2_clk;
    logic [31:0] top_9_2_out;
    logic top_9_2_done;
    logic [31:0] left_9_2_in;
    logic left_9_2_write_en;
    logic left_9_2_clk;
    logic [31:0] left_9_2_out;
    logic left_9_2_done;
    logic [31:0] pe_9_3_top;
    logic [31:0] pe_9_3_left;
    logic [31:0] pe_9_3_out;
    logic pe_9_3_go;
    logic pe_9_3_clk;
    logic pe_9_3_done;
    logic [31:0] top_9_3_in;
    logic top_9_3_write_en;
    logic top_9_3_clk;
    logic [31:0] top_9_3_out;
    logic top_9_3_done;
    logic [31:0] left_9_3_in;
    logic left_9_3_write_en;
    logic left_9_3_clk;
    logic [31:0] left_9_3_out;
    logic left_9_3_done;
    logic [31:0] pe_9_4_top;
    logic [31:0] pe_9_4_left;
    logic [31:0] pe_9_4_out;
    logic pe_9_4_go;
    logic pe_9_4_clk;
    logic pe_9_4_done;
    logic [31:0] top_9_4_in;
    logic top_9_4_write_en;
    logic top_9_4_clk;
    logic [31:0] top_9_4_out;
    logic top_9_4_done;
    logic [31:0] left_9_4_in;
    logic left_9_4_write_en;
    logic left_9_4_clk;
    logic [31:0] left_9_4_out;
    logic left_9_4_done;
    logic [31:0] pe_9_5_top;
    logic [31:0] pe_9_5_left;
    logic [31:0] pe_9_5_out;
    logic pe_9_5_go;
    logic pe_9_5_clk;
    logic pe_9_5_done;
    logic [31:0] top_9_5_in;
    logic top_9_5_write_en;
    logic top_9_5_clk;
    logic [31:0] top_9_5_out;
    logic top_9_5_done;
    logic [31:0] left_9_5_in;
    logic left_9_5_write_en;
    logic left_9_5_clk;
    logic [31:0] left_9_5_out;
    logic left_9_5_done;
    logic [31:0] pe_9_6_top;
    logic [31:0] pe_9_6_left;
    logic [31:0] pe_9_6_out;
    logic pe_9_6_go;
    logic pe_9_6_clk;
    logic pe_9_6_done;
    logic [31:0] top_9_6_in;
    logic top_9_6_write_en;
    logic top_9_6_clk;
    logic [31:0] top_9_6_out;
    logic top_9_6_done;
    logic [31:0] left_9_6_in;
    logic left_9_6_write_en;
    logic left_9_6_clk;
    logic [31:0] left_9_6_out;
    logic left_9_6_done;
    logic [31:0] pe_9_7_top;
    logic [31:0] pe_9_7_left;
    logic [31:0] pe_9_7_out;
    logic pe_9_7_go;
    logic pe_9_7_clk;
    logic pe_9_7_done;
    logic [31:0] top_9_7_in;
    logic top_9_7_write_en;
    logic top_9_7_clk;
    logic [31:0] top_9_7_out;
    logic top_9_7_done;
    logic [31:0] left_9_7_in;
    logic left_9_7_write_en;
    logic left_9_7_clk;
    logic [31:0] left_9_7_out;
    logic left_9_7_done;
    logic [31:0] pe_9_8_top;
    logic [31:0] pe_9_8_left;
    logic [31:0] pe_9_8_out;
    logic pe_9_8_go;
    logic pe_9_8_clk;
    logic pe_9_8_done;
    logic [31:0] top_9_8_in;
    logic top_9_8_write_en;
    logic top_9_8_clk;
    logic [31:0] top_9_8_out;
    logic top_9_8_done;
    logic [31:0] left_9_8_in;
    logic left_9_8_write_en;
    logic left_9_8_clk;
    logic [31:0] left_9_8_out;
    logic left_9_8_done;
    logic [31:0] pe_9_9_top;
    logic [31:0] pe_9_9_left;
    logic [31:0] pe_9_9_out;
    logic pe_9_9_go;
    logic pe_9_9_clk;
    logic pe_9_9_done;
    logic [31:0] top_9_9_in;
    logic top_9_9_write_en;
    logic top_9_9_clk;
    logic [31:0] top_9_9_out;
    logic top_9_9_done;
    logic [31:0] left_9_9_in;
    logic left_9_9_write_en;
    logic left_9_9_clk;
    logic [31:0] left_9_9_out;
    logic left_9_9_done;
    logic [31:0] pe_9_10_top;
    logic [31:0] pe_9_10_left;
    logic [31:0] pe_9_10_out;
    logic pe_9_10_go;
    logic pe_9_10_clk;
    logic pe_9_10_done;
    logic [31:0] top_9_10_in;
    logic top_9_10_write_en;
    logic top_9_10_clk;
    logic [31:0] top_9_10_out;
    logic top_9_10_done;
    logic [31:0] left_9_10_in;
    logic left_9_10_write_en;
    logic left_9_10_clk;
    logic [31:0] left_9_10_out;
    logic left_9_10_done;
    logic [31:0] pe_9_11_top;
    logic [31:0] pe_9_11_left;
    logic [31:0] pe_9_11_out;
    logic pe_9_11_go;
    logic pe_9_11_clk;
    logic pe_9_11_done;
    logic [31:0] top_9_11_in;
    logic top_9_11_write_en;
    logic top_9_11_clk;
    logic [31:0] top_9_11_out;
    logic top_9_11_done;
    logic [31:0] left_9_11_in;
    logic left_9_11_write_en;
    logic left_9_11_clk;
    logic [31:0] left_9_11_out;
    logic left_9_11_done;
    logic [31:0] pe_9_12_top;
    logic [31:0] pe_9_12_left;
    logic [31:0] pe_9_12_out;
    logic pe_9_12_go;
    logic pe_9_12_clk;
    logic pe_9_12_done;
    logic [31:0] top_9_12_in;
    logic top_9_12_write_en;
    logic top_9_12_clk;
    logic [31:0] top_9_12_out;
    logic top_9_12_done;
    logic [31:0] left_9_12_in;
    logic left_9_12_write_en;
    logic left_9_12_clk;
    logic [31:0] left_9_12_out;
    logic left_9_12_done;
    logic [31:0] pe_9_13_top;
    logic [31:0] pe_9_13_left;
    logic [31:0] pe_9_13_out;
    logic pe_9_13_go;
    logic pe_9_13_clk;
    logic pe_9_13_done;
    logic [31:0] top_9_13_in;
    logic top_9_13_write_en;
    logic top_9_13_clk;
    logic [31:0] top_9_13_out;
    logic top_9_13_done;
    logic [31:0] left_9_13_in;
    logic left_9_13_write_en;
    logic left_9_13_clk;
    logic [31:0] left_9_13_out;
    logic left_9_13_done;
    logic [31:0] pe_9_14_top;
    logic [31:0] pe_9_14_left;
    logic [31:0] pe_9_14_out;
    logic pe_9_14_go;
    logic pe_9_14_clk;
    logic pe_9_14_done;
    logic [31:0] top_9_14_in;
    logic top_9_14_write_en;
    logic top_9_14_clk;
    logic [31:0] top_9_14_out;
    logic top_9_14_done;
    logic [31:0] left_9_14_in;
    logic left_9_14_write_en;
    logic left_9_14_clk;
    logic [31:0] left_9_14_out;
    logic left_9_14_done;
    logic [31:0] pe_9_15_top;
    logic [31:0] pe_9_15_left;
    logic [31:0] pe_9_15_out;
    logic pe_9_15_go;
    logic pe_9_15_clk;
    logic pe_9_15_done;
    logic [31:0] top_9_15_in;
    logic top_9_15_write_en;
    logic top_9_15_clk;
    logic [31:0] top_9_15_out;
    logic top_9_15_done;
    logic [31:0] left_9_15_in;
    logic left_9_15_write_en;
    logic left_9_15_clk;
    logic [31:0] left_9_15_out;
    logic left_9_15_done;
    logic [31:0] pe_10_0_top;
    logic [31:0] pe_10_0_left;
    logic [31:0] pe_10_0_out;
    logic pe_10_0_go;
    logic pe_10_0_clk;
    logic pe_10_0_done;
    logic [31:0] top_10_0_in;
    logic top_10_0_write_en;
    logic top_10_0_clk;
    logic [31:0] top_10_0_out;
    logic top_10_0_done;
    logic [31:0] left_10_0_in;
    logic left_10_0_write_en;
    logic left_10_0_clk;
    logic [31:0] left_10_0_out;
    logic left_10_0_done;
    logic [31:0] pe_10_1_top;
    logic [31:0] pe_10_1_left;
    logic [31:0] pe_10_1_out;
    logic pe_10_1_go;
    logic pe_10_1_clk;
    logic pe_10_1_done;
    logic [31:0] top_10_1_in;
    logic top_10_1_write_en;
    logic top_10_1_clk;
    logic [31:0] top_10_1_out;
    logic top_10_1_done;
    logic [31:0] left_10_1_in;
    logic left_10_1_write_en;
    logic left_10_1_clk;
    logic [31:0] left_10_1_out;
    logic left_10_1_done;
    logic [31:0] pe_10_2_top;
    logic [31:0] pe_10_2_left;
    logic [31:0] pe_10_2_out;
    logic pe_10_2_go;
    logic pe_10_2_clk;
    logic pe_10_2_done;
    logic [31:0] top_10_2_in;
    logic top_10_2_write_en;
    logic top_10_2_clk;
    logic [31:0] top_10_2_out;
    logic top_10_2_done;
    logic [31:0] left_10_2_in;
    logic left_10_2_write_en;
    logic left_10_2_clk;
    logic [31:0] left_10_2_out;
    logic left_10_2_done;
    logic [31:0] pe_10_3_top;
    logic [31:0] pe_10_3_left;
    logic [31:0] pe_10_3_out;
    logic pe_10_3_go;
    logic pe_10_3_clk;
    logic pe_10_3_done;
    logic [31:0] top_10_3_in;
    logic top_10_3_write_en;
    logic top_10_3_clk;
    logic [31:0] top_10_3_out;
    logic top_10_3_done;
    logic [31:0] left_10_3_in;
    logic left_10_3_write_en;
    logic left_10_3_clk;
    logic [31:0] left_10_3_out;
    logic left_10_3_done;
    logic [31:0] pe_10_4_top;
    logic [31:0] pe_10_4_left;
    logic [31:0] pe_10_4_out;
    logic pe_10_4_go;
    logic pe_10_4_clk;
    logic pe_10_4_done;
    logic [31:0] top_10_4_in;
    logic top_10_4_write_en;
    logic top_10_4_clk;
    logic [31:0] top_10_4_out;
    logic top_10_4_done;
    logic [31:0] left_10_4_in;
    logic left_10_4_write_en;
    logic left_10_4_clk;
    logic [31:0] left_10_4_out;
    logic left_10_4_done;
    logic [31:0] pe_10_5_top;
    logic [31:0] pe_10_5_left;
    logic [31:0] pe_10_5_out;
    logic pe_10_5_go;
    logic pe_10_5_clk;
    logic pe_10_5_done;
    logic [31:0] top_10_5_in;
    logic top_10_5_write_en;
    logic top_10_5_clk;
    logic [31:0] top_10_5_out;
    logic top_10_5_done;
    logic [31:0] left_10_5_in;
    logic left_10_5_write_en;
    logic left_10_5_clk;
    logic [31:0] left_10_5_out;
    logic left_10_5_done;
    logic [31:0] pe_10_6_top;
    logic [31:0] pe_10_6_left;
    logic [31:0] pe_10_6_out;
    logic pe_10_6_go;
    logic pe_10_6_clk;
    logic pe_10_6_done;
    logic [31:0] top_10_6_in;
    logic top_10_6_write_en;
    logic top_10_6_clk;
    logic [31:0] top_10_6_out;
    logic top_10_6_done;
    logic [31:0] left_10_6_in;
    logic left_10_6_write_en;
    logic left_10_6_clk;
    logic [31:0] left_10_6_out;
    logic left_10_6_done;
    logic [31:0] pe_10_7_top;
    logic [31:0] pe_10_7_left;
    logic [31:0] pe_10_7_out;
    logic pe_10_7_go;
    logic pe_10_7_clk;
    logic pe_10_7_done;
    logic [31:0] top_10_7_in;
    logic top_10_7_write_en;
    logic top_10_7_clk;
    logic [31:0] top_10_7_out;
    logic top_10_7_done;
    logic [31:0] left_10_7_in;
    logic left_10_7_write_en;
    logic left_10_7_clk;
    logic [31:0] left_10_7_out;
    logic left_10_7_done;
    logic [31:0] pe_10_8_top;
    logic [31:0] pe_10_8_left;
    logic [31:0] pe_10_8_out;
    logic pe_10_8_go;
    logic pe_10_8_clk;
    logic pe_10_8_done;
    logic [31:0] top_10_8_in;
    logic top_10_8_write_en;
    logic top_10_8_clk;
    logic [31:0] top_10_8_out;
    logic top_10_8_done;
    logic [31:0] left_10_8_in;
    logic left_10_8_write_en;
    logic left_10_8_clk;
    logic [31:0] left_10_8_out;
    logic left_10_8_done;
    logic [31:0] pe_10_9_top;
    logic [31:0] pe_10_9_left;
    logic [31:0] pe_10_9_out;
    logic pe_10_9_go;
    logic pe_10_9_clk;
    logic pe_10_9_done;
    logic [31:0] top_10_9_in;
    logic top_10_9_write_en;
    logic top_10_9_clk;
    logic [31:0] top_10_9_out;
    logic top_10_9_done;
    logic [31:0] left_10_9_in;
    logic left_10_9_write_en;
    logic left_10_9_clk;
    logic [31:0] left_10_9_out;
    logic left_10_9_done;
    logic [31:0] pe_10_10_top;
    logic [31:0] pe_10_10_left;
    logic [31:0] pe_10_10_out;
    logic pe_10_10_go;
    logic pe_10_10_clk;
    logic pe_10_10_done;
    logic [31:0] top_10_10_in;
    logic top_10_10_write_en;
    logic top_10_10_clk;
    logic [31:0] top_10_10_out;
    logic top_10_10_done;
    logic [31:0] left_10_10_in;
    logic left_10_10_write_en;
    logic left_10_10_clk;
    logic [31:0] left_10_10_out;
    logic left_10_10_done;
    logic [31:0] pe_10_11_top;
    logic [31:0] pe_10_11_left;
    logic [31:0] pe_10_11_out;
    logic pe_10_11_go;
    logic pe_10_11_clk;
    logic pe_10_11_done;
    logic [31:0] top_10_11_in;
    logic top_10_11_write_en;
    logic top_10_11_clk;
    logic [31:0] top_10_11_out;
    logic top_10_11_done;
    logic [31:0] left_10_11_in;
    logic left_10_11_write_en;
    logic left_10_11_clk;
    logic [31:0] left_10_11_out;
    logic left_10_11_done;
    logic [31:0] pe_10_12_top;
    logic [31:0] pe_10_12_left;
    logic [31:0] pe_10_12_out;
    logic pe_10_12_go;
    logic pe_10_12_clk;
    logic pe_10_12_done;
    logic [31:0] top_10_12_in;
    logic top_10_12_write_en;
    logic top_10_12_clk;
    logic [31:0] top_10_12_out;
    logic top_10_12_done;
    logic [31:0] left_10_12_in;
    logic left_10_12_write_en;
    logic left_10_12_clk;
    logic [31:0] left_10_12_out;
    logic left_10_12_done;
    logic [31:0] pe_10_13_top;
    logic [31:0] pe_10_13_left;
    logic [31:0] pe_10_13_out;
    logic pe_10_13_go;
    logic pe_10_13_clk;
    logic pe_10_13_done;
    logic [31:0] top_10_13_in;
    logic top_10_13_write_en;
    logic top_10_13_clk;
    logic [31:0] top_10_13_out;
    logic top_10_13_done;
    logic [31:0] left_10_13_in;
    logic left_10_13_write_en;
    logic left_10_13_clk;
    logic [31:0] left_10_13_out;
    logic left_10_13_done;
    logic [31:0] pe_10_14_top;
    logic [31:0] pe_10_14_left;
    logic [31:0] pe_10_14_out;
    logic pe_10_14_go;
    logic pe_10_14_clk;
    logic pe_10_14_done;
    logic [31:0] top_10_14_in;
    logic top_10_14_write_en;
    logic top_10_14_clk;
    logic [31:0] top_10_14_out;
    logic top_10_14_done;
    logic [31:0] left_10_14_in;
    logic left_10_14_write_en;
    logic left_10_14_clk;
    logic [31:0] left_10_14_out;
    logic left_10_14_done;
    logic [31:0] pe_10_15_top;
    logic [31:0] pe_10_15_left;
    logic [31:0] pe_10_15_out;
    logic pe_10_15_go;
    logic pe_10_15_clk;
    logic pe_10_15_done;
    logic [31:0] top_10_15_in;
    logic top_10_15_write_en;
    logic top_10_15_clk;
    logic [31:0] top_10_15_out;
    logic top_10_15_done;
    logic [31:0] left_10_15_in;
    logic left_10_15_write_en;
    logic left_10_15_clk;
    logic [31:0] left_10_15_out;
    logic left_10_15_done;
    logic [31:0] pe_11_0_top;
    logic [31:0] pe_11_0_left;
    logic [31:0] pe_11_0_out;
    logic pe_11_0_go;
    logic pe_11_0_clk;
    logic pe_11_0_done;
    logic [31:0] top_11_0_in;
    logic top_11_0_write_en;
    logic top_11_0_clk;
    logic [31:0] top_11_0_out;
    logic top_11_0_done;
    logic [31:0] left_11_0_in;
    logic left_11_0_write_en;
    logic left_11_0_clk;
    logic [31:0] left_11_0_out;
    logic left_11_0_done;
    logic [31:0] pe_11_1_top;
    logic [31:0] pe_11_1_left;
    logic [31:0] pe_11_1_out;
    logic pe_11_1_go;
    logic pe_11_1_clk;
    logic pe_11_1_done;
    logic [31:0] top_11_1_in;
    logic top_11_1_write_en;
    logic top_11_1_clk;
    logic [31:0] top_11_1_out;
    logic top_11_1_done;
    logic [31:0] left_11_1_in;
    logic left_11_1_write_en;
    logic left_11_1_clk;
    logic [31:0] left_11_1_out;
    logic left_11_1_done;
    logic [31:0] pe_11_2_top;
    logic [31:0] pe_11_2_left;
    logic [31:0] pe_11_2_out;
    logic pe_11_2_go;
    logic pe_11_2_clk;
    logic pe_11_2_done;
    logic [31:0] top_11_2_in;
    logic top_11_2_write_en;
    logic top_11_2_clk;
    logic [31:0] top_11_2_out;
    logic top_11_2_done;
    logic [31:0] left_11_2_in;
    logic left_11_2_write_en;
    logic left_11_2_clk;
    logic [31:0] left_11_2_out;
    logic left_11_2_done;
    logic [31:0] pe_11_3_top;
    logic [31:0] pe_11_3_left;
    logic [31:0] pe_11_3_out;
    logic pe_11_3_go;
    logic pe_11_3_clk;
    logic pe_11_3_done;
    logic [31:0] top_11_3_in;
    logic top_11_3_write_en;
    logic top_11_3_clk;
    logic [31:0] top_11_3_out;
    logic top_11_3_done;
    logic [31:0] left_11_3_in;
    logic left_11_3_write_en;
    logic left_11_3_clk;
    logic [31:0] left_11_3_out;
    logic left_11_3_done;
    logic [31:0] pe_11_4_top;
    logic [31:0] pe_11_4_left;
    logic [31:0] pe_11_4_out;
    logic pe_11_4_go;
    logic pe_11_4_clk;
    logic pe_11_4_done;
    logic [31:0] top_11_4_in;
    logic top_11_4_write_en;
    logic top_11_4_clk;
    logic [31:0] top_11_4_out;
    logic top_11_4_done;
    logic [31:0] left_11_4_in;
    logic left_11_4_write_en;
    logic left_11_4_clk;
    logic [31:0] left_11_4_out;
    logic left_11_4_done;
    logic [31:0] pe_11_5_top;
    logic [31:0] pe_11_5_left;
    logic [31:0] pe_11_5_out;
    logic pe_11_5_go;
    logic pe_11_5_clk;
    logic pe_11_5_done;
    logic [31:0] top_11_5_in;
    logic top_11_5_write_en;
    logic top_11_5_clk;
    logic [31:0] top_11_5_out;
    logic top_11_5_done;
    logic [31:0] left_11_5_in;
    logic left_11_5_write_en;
    logic left_11_5_clk;
    logic [31:0] left_11_5_out;
    logic left_11_5_done;
    logic [31:0] pe_11_6_top;
    logic [31:0] pe_11_6_left;
    logic [31:0] pe_11_6_out;
    logic pe_11_6_go;
    logic pe_11_6_clk;
    logic pe_11_6_done;
    logic [31:0] top_11_6_in;
    logic top_11_6_write_en;
    logic top_11_6_clk;
    logic [31:0] top_11_6_out;
    logic top_11_6_done;
    logic [31:0] left_11_6_in;
    logic left_11_6_write_en;
    logic left_11_6_clk;
    logic [31:0] left_11_6_out;
    logic left_11_6_done;
    logic [31:0] pe_11_7_top;
    logic [31:0] pe_11_7_left;
    logic [31:0] pe_11_7_out;
    logic pe_11_7_go;
    logic pe_11_7_clk;
    logic pe_11_7_done;
    logic [31:0] top_11_7_in;
    logic top_11_7_write_en;
    logic top_11_7_clk;
    logic [31:0] top_11_7_out;
    logic top_11_7_done;
    logic [31:0] left_11_7_in;
    logic left_11_7_write_en;
    logic left_11_7_clk;
    logic [31:0] left_11_7_out;
    logic left_11_7_done;
    logic [31:0] pe_11_8_top;
    logic [31:0] pe_11_8_left;
    logic [31:0] pe_11_8_out;
    logic pe_11_8_go;
    logic pe_11_8_clk;
    logic pe_11_8_done;
    logic [31:0] top_11_8_in;
    logic top_11_8_write_en;
    logic top_11_8_clk;
    logic [31:0] top_11_8_out;
    logic top_11_8_done;
    logic [31:0] left_11_8_in;
    logic left_11_8_write_en;
    logic left_11_8_clk;
    logic [31:0] left_11_8_out;
    logic left_11_8_done;
    logic [31:0] pe_11_9_top;
    logic [31:0] pe_11_9_left;
    logic [31:0] pe_11_9_out;
    logic pe_11_9_go;
    logic pe_11_9_clk;
    logic pe_11_9_done;
    logic [31:0] top_11_9_in;
    logic top_11_9_write_en;
    logic top_11_9_clk;
    logic [31:0] top_11_9_out;
    logic top_11_9_done;
    logic [31:0] left_11_9_in;
    logic left_11_9_write_en;
    logic left_11_9_clk;
    logic [31:0] left_11_9_out;
    logic left_11_9_done;
    logic [31:0] pe_11_10_top;
    logic [31:0] pe_11_10_left;
    logic [31:0] pe_11_10_out;
    logic pe_11_10_go;
    logic pe_11_10_clk;
    logic pe_11_10_done;
    logic [31:0] top_11_10_in;
    logic top_11_10_write_en;
    logic top_11_10_clk;
    logic [31:0] top_11_10_out;
    logic top_11_10_done;
    logic [31:0] left_11_10_in;
    logic left_11_10_write_en;
    logic left_11_10_clk;
    logic [31:0] left_11_10_out;
    logic left_11_10_done;
    logic [31:0] pe_11_11_top;
    logic [31:0] pe_11_11_left;
    logic [31:0] pe_11_11_out;
    logic pe_11_11_go;
    logic pe_11_11_clk;
    logic pe_11_11_done;
    logic [31:0] top_11_11_in;
    logic top_11_11_write_en;
    logic top_11_11_clk;
    logic [31:0] top_11_11_out;
    logic top_11_11_done;
    logic [31:0] left_11_11_in;
    logic left_11_11_write_en;
    logic left_11_11_clk;
    logic [31:0] left_11_11_out;
    logic left_11_11_done;
    logic [31:0] pe_11_12_top;
    logic [31:0] pe_11_12_left;
    logic [31:0] pe_11_12_out;
    logic pe_11_12_go;
    logic pe_11_12_clk;
    logic pe_11_12_done;
    logic [31:0] top_11_12_in;
    logic top_11_12_write_en;
    logic top_11_12_clk;
    logic [31:0] top_11_12_out;
    logic top_11_12_done;
    logic [31:0] left_11_12_in;
    logic left_11_12_write_en;
    logic left_11_12_clk;
    logic [31:0] left_11_12_out;
    logic left_11_12_done;
    logic [31:0] pe_11_13_top;
    logic [31:0] pe_11_13_left;
    logic [31:0] pe_11_13_out;
    logic pe_11_13_go;
    logic pe_11_13_clk;
    logic pe_11_13_done;
    logic [31:0] top_11_13_in;
    logic top_11_13_write_en;
    logic top_11_13_clk;
    logic [31:0] top_11_13_out;
    logic top_11_13_done;
    logic [31:0] left_11_13_in;
    logic left_11_13_write_en;
    logic left_11_13_clk;
    logic [31:0] left_11_13_out;
    logic left_11_13_done;
    logic [31:0] pe_11_14_top;
    logic [31:0] pe_11_14_left;
    logic [31:0] pe_11_14_out;
    logic pe_11_14_go;
    logic pe_11_14_clk;
    logic pe_11_14_done;
    logic [31:0] top_11_14_in;
    logic top_11_14_write_en;
    logic top_11_14_clk;
    logic [31:0] top_11_14_out;
    logic top_11_14_done;
    logic [31:0] left_11_14_in;
    logic left_11_14_write_en;
    logic left_11_14_clk;
    logic [31:0] left_11_14_out;
    logic left_11_14_done;
    logic [31:0] pe_11_15_top;
    logic [31:0] pe_11_15_left;
    logic [31:0] pe_11_15_out;
    logic pe_11_15_go;
    logic pe_11_15_clk;
    logic pe_11_15_done;
    logic [31:0] top_11_15_in;
    logic top_11_15_write_en;
    logic top_11_15_clk;
    logic [31:0] top_11_15_out;
    logic top_11_15_done;
    logic [31:0] left_11_15_in;
    logic left_11_15_write_en;
    logic left_11_15_clk;
    logic [31:0] left_11_15_out;
    logic left_11_15_done;
    logic [31:0] pe_12_0_top;
    logic [31:0] pe_12_0_left;
    logic [31:0] pe_12_0_out;
    logic pe_12_0_go;
    logic pe_12_0_clk;
    logic pe_12_0_done;
    logic [31:0] top_12_0_in;
    logic top_12_0_write_en;
    logic top_12_0_clk;
    logic [31:0] top_12_0_out;
    logic top_12_0_done;
    logic [31:0] left_12_0_in;
    logic left_12_0_write_en;
    logic left_12_0_clk;
    logic [31:0] left_12_0_out;
    logic left_12_0_done;
    logic [31:0] pe_12_1_top;
    logic [31:0] pe_12_1_left;
    logic [31:0] pe_12_1_out;
    logic pe_12_1_go;
    logic pe_12_1_clk;
    logic pe_12_1_done;
    logic [31:0] top_12_1_in;
    logic top_12_1_write_en;
    logic top_12_1_clk;
    logic [31:0] top_12_1_out;
    logic top_12_1_done;
    logic [31:0] left_12_1_in;
    logic left_12_1_write_en;
    logic left_12_1_clk;
    logic [31:0] left_12_1_out;
    logic left_12_1_done;
    logic [31:0] pe_12_2_top;
    logic [31:0] pe_12_2_left;
    logic [31:0] pe_12_2_out;
    logic pe_12_2_go;
    logic pe_12_2_clk;
    logic pe_12_2_done;
    logic [31:0] top_12_2_in;
    logic top_12_2_write_en;
    logic top_12_2_clk;
    logic [31:0] top_12_2_out;
    logic top_12_2_done;
    logic [31:0] left_12_2_in;
    logic left_12_2_write_en;
    logic left_12_2_clk;
    logic [31:0] left_12_2_out;
    logic left_12_2_done;
    logic [31:0] pe_12_3_top;
    logic [31:0] pe_12_3_left;
    logic [31:0] pe_12_3_out;
    logic pe_12_3_go;
    logic pe_12_3_clk;
    logic pe_12_3_done;
    logic [31:0] top_12_3_in;
    logic top_12_3_write_en;
    logic top_12_3_clk;
    logic [31:0] top_12_3_out;
    logic top_12_3_done;
    logic [31:0] left_12_3_in;
    logic left_12_3_write_en;
    logic left_12_3_clk;
    logic [31:0] left_12_3_out;
    logic left_12_3_done;
    logic [31:0] pe_12_4_top;
    logic [31:0] pe_12_4_left;
    logic [31:0] pe_12_4_out;
    logic pe_12_4_go;
    logic pe_12_4_clk;
    logic pe_12_4_done;
    logic [31:0] top_12_4_in;
    logic top_12_4_write_en;
    logic top_12_4_clk;
    logic [31:0] top_12_4_out;
    logic top_12_4_done;
    logic [31:0] left_12_4_in;
    logic left_12_4_write_en;
    logic left_12_4_clk;
    logic [31:0] left_12_4_out;
    logic left_12_4_done;
    logic [31:0] pe_12_5_top;
    logic [31:0] pe_12_5_left;
    logic [31:0] pe_12_5_out;
    logic pe_12_5_go;
    logic pe_12_5_clk;
    logic pe_12_5_done;
    logic [31:0] top_12_5_in;
    logic top_12_5_write_en;
    logic top_12_5_clk;
    logic [31:0] top_12_5_out;
    logic top_12_5_done;
    logic [31:0] left_12_5_in;
    logic left_12_5_write_en;
    logic left_12_5_clk;
    logic [31:0] left_12_5_out;
    logic left_12_5_done;
    logic [31:0] pe_12_6_top;
    logic [31:0] pe_12_6_left;
    logic [31:0] pe_12_6_out;
    logic pe_12_6_go;
    logic pe_12_6_clk;
    logic pe_12_6_done;
    logic [31:0] top_12_6_in;
    logic top_12_6_write_en;
    logic top_12_6_clk;
    logic [31:0] top_12_6_out;
    logic top_12_6_done;
    logic [31:0] left_12_6_in;
    logic left_12_6_write_en;
    logic left_12_6_clk;
    logic [31:0] left_12_6_out;
    logic left_12_6_done;
    logic [31:0] pe_12_7_top;
    logic [31:0] pe_12_7_left;
    logic [31:0] pe_12_7_out;
    logic pe_12_7_go;
    logic pe_12_7_clk;
    logic pe_12_7_done;
    logic [31:0] top_12_7_in;
    logic top_12_7_write_en;
    logic top_12_7_clk;
    logic [31:0] top_12_7_out;
    logic top_12_7_done;
    logic [31:0] left_12_7_in;
    logic left_12_7_write_en;
    logic left_12_7_clk;
    logic [31:0] left_12_7_out;
    logic left_12_7_done;
    logic [31:0] pe_12_8_top;
    logic [31:0] pe_12_8_left;
    logic [31:0] pe_12_8_out;
    logic pe_12_8_go;
    logic pe_12_8_clk;
    logic pe_12_8_done;
    logic [31:0] top_12_8_in;
    logic top_12_8_write_en;
    logic top_12_8_clk;
    logic [31:0] top_12_8_out;
    logic top_12_8_done;
    logic [31:0] left_12_8_in;
    logic left_12_8_write_en;
    logic left_12_8_clk;
    logic [31:0] left_12_8_out;
    logic left_12_8_done;
    logic [31:0] pe_12_9_top;
    logic [31:0] pe_12_9_left;
    logic [31:0] pe_12_9_out;
    logic pe_12_9_go;
    logic pe_12_9_clk;
    logic pe_12_9_done;
    logic [31:0] top_12_9_in;
    logic top_12_9_write_en;
    logic top_12_9_clk;
    logic [31:0] top_12_9_out;
    logic top_12_9_done;
    logic [31:0] left_12_9_in;
    logic left_12_9_write_en;
    logic left_12_9_clk;
    logic [31:0] left_12_9_out;
    logic left_12_9_done;
    logic [31:0] pe_12_10_top;
    logic [31:0] pe_12_10_left;
    logic [31:0] pe_12_10_out;
    logic pe_12_10_go;
    logic pe_12_10_clk;
    logic pe_12_10_done;
    logic [31:0] top_12_10_in;
    logic top_12_10_write_en;
    logic top_12_10_clk;
    logic [31:0] top_12_10_out;
    logic top_12_10_done;
    logic [31:0] left_12_10_in;
    logic left_12_10_write_en;
    logic left_12_10_clk;
    logic [31:0] left_12_10_out;
    logic left_12_10_done;
    logic [31:0] pe_12_11_top;
    logic [31:0] pe_12_11_left;
    logic [31:0] pe_12_11_out;
    logic pe_12_11_go;
    logic pe_12_11_clk;
    logic pe_12_11_done;
    logic [31:0] top_12_11_in;
    logic top_12_11_write_en;
    logic top_12_11_clk;
    logic [31:0] top_12_11_out;
    logic top_12_11_done;
    logic [31:0] left_12_11_in;
    logic left_12_11_write_en;
    logic left_12_11_clk;
    logic [31:0] left_12_11_out;
    logic left_12_11_done;
    logic [31:0] pe_12_12_top;
    logic [31:0] pe_12_12_left;
    logic [31:0] pe_12_12_out;
    logic pe_12_12_go;
    logic pe_12_12_clk;
    logic pe_12_12_done;
    logic [31:0] top_12_12_in;
    logic top_12_12_write_en;
    logic top_12_12_clk;
    logic [31:0] top_12_12_out;
    logic top_12_12_done;
    logic [31:0] left_12_12_in;
    logic left_12_12_write_en;
    logic left_12_12_clk;
    logic [31:0] left_12_12_out;
    logic left_12_12_done;
    logic [31:0] pe_12_13_top;
    logic [31:0] pe_12_13_left;
    logic [31:0] pe_12_13_out;
    logic pe_12_13_go;
    logic pe_12_13_clk;
    logic pe_12_13_done;
    logic [31:0] top_12_13_in;
    logic top_12_13_write_en;
    logic top_12_13_clk;
    logic [31:0] top_12_13_out;
    logic top_12_13_done;
    logic [31:0] left_12_13_in;
    logic left_12_13_write_en;
    logic left_12_13_clk;
    logic [31:0] left_12_13_out;
    logic left_12_13_done;
    logic [31:0] pe_12_14_top;
    logic [31:0] pe_12_14_left;
    logic [31:0] pe_12_14_out;
    logic pe_12_14_go;
    logic pe_12_14_clk;
    logic pe_12_14_done;
    logic [31:0] top_12_14_in;
    logic top_12_14_write_en;
    logic top_12_14_clk;
    logic [31:0] top_12_14_out;
    logic top_12_14_done;
    logic [31:0] left_12_14_in;
    logic left_12_14_write_en;
    logic left_12_14_clk;
    logic [31:0] left_12_14_out;
    logic left_12_14_done;
    logic [31:0] pe_12_15_top;
    logic [31:0] pe_12_15_left;
    logic [31:0] pe_12_15_out;
    logic pe_12_15_go;
    logic pe_12_15_clk;
    logic pe_12_15_done;
    logic [31:0] top_12_15_in;
    logic top_12_15_write_en;
    logic top_12_15_clk;
    logic [31:0] top_12_15_out;
    logic top_12_15_done;
    logic [31:0] left_12_15_in;
    logic left_12_15_write_en;
    logic left_12_15_clk;
    logic [31:0] left_12_15_out;
    logic left_12_15_done;
    logic [31:0] pe_13_0_top;
    logic [31:0] pe_13_0_left;
    logic [31:0] pe_13_0_out;
    logic pe_13_0_go;
    logic pe_13_0_clk;
    logic pe_13_0_done;
    logic [31:0] top_13_0_in;
    logic top_13_0_write_en;
    logic top_13_0_clk;
    logic [31:0] top_13_0_out;
    logic top_13_0_done;
    logic [31:0] left_13_0_in;
    logic left_13_0_write_en;
    logic left_13_0_clk;
    logic [31:0] left_13_0_out;
    logic left_13_0_done;
    logic [31:0] pe_13_1_top;
    logic [31:0] pe_13_1_left;
    logic [31:0] pe_13_1_out;
    logic pe_13_1_go;
    logic pe_13_1_clk;
    logic pe_13_1_done;
    logic [31:0] top_13_1_in;
    logic top_13_1_write_en;
    logic top_13_1_clk;
    logic [31:0] top_13_1_out;
    logic top_13_1_done;
    logic [31:0] left_13_1_in;
    logic left_13_1_write_en;
    logic left_13_1_clk;
    logic [31:0] left_13_1_out;
    logic left_13_1_done;
    logic [31:0] pe_13_2_top;
    logic [31:0] pe_13_2_left;
    logic [31:0] pe_13_2_out;
    logic pe_13_2_go;
    logic pe_13_2_clk;
    logic pe_13_2_done;
    logic [31:0] top_13_2_in;
    logic top_13_2_write_en;
    logic top_13_2_clk;
    logic [31:0] top_13_2_out;
    logic top_13_2_done;
    logic [31:0] left_13_2_in;
    logic left_13_2_write_en;
    logic left_13_2_clk;
    logic [31:0] left_13_2_out;
    logic left_13_2_done;
    logic [31:0] pe_13_3_top;
    logic [31:0] pe_13_3_left;
    logic [31:0] pe_13_3_out;
    logic pe_13_3_go;
    logic pe_13_3_clk;
    logic pe_13_3_done;
    logic [31:0] top_13_3_in;
    logic top_13_3_write_en;
    logic top_13_3_clk;
    logic [31:0] top_13_3_out;
    logic top_13_3_done;
    logic [31:0] left_13_3_in;
    logic left_13_3_write_en;
    logic left_13_3_clk;
    logic [31:0] left_13_3_out;
    logic left_13_3_done;
    logic [31:0] pe_13_4_top;
    logic [31:0] pe_13_4_left;
    logic [31:0] pe_13_4_out;
    logic pe_13_4_go;
    logic pe_13_4_clk;
    logic pe_13_4_done;
    logic [31:0] top_13_4_in;
    logic top_13_4_write_en;
    logic top_13_4_clk;
    logic [31:0] top_13_4_out;
    logic top_13_4_done;
    logic [31:0] left_13_4_in;
    logic left_13_4_write_en;
    logic left_13_4_clk;
    logic [31:0] left_13_4_out;
    logic left_13_4_done;
    logic [31:0] pe_13_5_top;
    logic [31:0] pe_13_5_left;
    logic [31:0] pe_13_5_out;
    logic pe_13_5_go;
    logic pe_13_5_clk;
    logic pe_13_5_done;
    logic [31:0] top_13_5_in;
    logic top_13_5_write_en;
    logic top_13_5_clk;
    logic [31:0] top_13_5_out;
    logic top_13_5_done;
    logic [31:0] left_13_5_in;
    logic left_13_5_write_en;
    logic left_13_5_clk;
    logic [31:0] left_13_5_out;
    logic left_13_5_done;
    logic [31:0] pe_13_6_top;
    logic [31:0] pe_13_6_left;
    logic [31:0] pe_13_6_out;
    logic pe_13_6_go;
    logic pe_13_6_clk;
    logic pe_13_6_done;
    logic [31:0] top_13_6_in;
    logic top_13_6_write_en;
    logic top_13_6_clk;
    logic [31:0] top_13_6_out;
    logic top_13_6_done;
    logic [31:0] left_13_6_in;
    logic left_13_6_write_en;
    logic left_13_6_clk;
    logic [31:0] left_13_6_out;
    logic left_13_6_done;
    logic [31:0] pe_13_7_top;
    logic [31:0] pe_13_7_left;
    logic [31:0] pe_13_7_out;
    logic pe_13_7_go;
    logic pe_13_7_clk;
    logic pe_13_7_done;
    logic [31:0] top_13_7_in;
    logic top_13_7_write_en;
    logic top_13_7_clk;
    logic [31:0] top_13_7_out;
    logic top_13_7_done;
    logic [31:0] left_13_7_in;
    logic left_13_7_write_en;
    logic left_13_7_clk;
    logic [31:0] left_13_7_out;
    logic left_13_7_done;
    logic [31:0] pe_13_8_top;
    logic [31:0] pe_13_8_left;
    logic [31:0] pe_13_8_out;
    logic pe_13_8_go;
    logic pe_13_8_clk;
    logic pe_13_8_done;
    logic [31:0] top_13_8_in;
    logic top_13_8_write_en;
    logic top_13_8_clk;
    logic [31:0] top_13_8_out;
    logic top_13_8_done;
    logic [31:0] left_13_8_in;
    logic left_13_8_write_en;
    logic left_13_8_clk;
    logic [31:0] left_13_8_out;
    logic left_13_8_done;
    logic [31:0] pe_13_9_top;
    logic [31:0] pe_13_9_left;
    logic [31:0] pe_13_9_out;
    logic pe_13_9_go;
    logic pe_13_9_clk;
    logic pe_13_9_done;
    logic [31:0] top_13_9_in;
    logic top_13_9_write_en;
    logic top_13_9_clk;
    logic [31:0] top_13_9_out;
    logic top_13_9_done;
    logic [31:0] left_13_9_in;
    logic left_13_9_write_en;
    logic left_13_9_clk;
    logic [31:0] left_13_9_out;
    logic left_13_9_done;
    logic [31:0] pe_13_10_top;
    logic [31:0] pe_13_10_left;
    logic [31:0] pe_13_10_out;
    logic pe_13_10_go;
    logic pe_13_10_clk;
    logic pe_13_10_done;
    logic [31:0] top_13_10_in;
    logic top_13_10_write_en;
    logic top_13_10_clk;
    logic [31:0] top_13_10_out;
    logic top_13_10_done;
    logic [31:0] left_13_10_in;
    logic left_13_10_write_en;
    logic left_13_10_clk;
    logic [31:0] left_13_10_out;
    logic left_13_10_done;
    logic [31:0] pe_13_11_top;
    logic [31:0] pe_13_11_left;
    logic [31:0] pe_13_11_out;
    logic pe_13_11_go;
    logic pe_13_11_clk;
    logic pe_13_11_done;
    logic [31:0] top_13_11_in;
    logic top_13_11_write_en;
    logic top_13_11_clk;
    logic [31:0] top_13_11_out;
    logic top_13_11_done;
    logic [31:0] left_13_11_in;
    logic left_13_11_write_en;
    logic left_13_11_clk;
    logic [31:0] left_13_11_out;
    logic left_13_11_done;
    logic [31:0] pe_13_12_top;
    logic [31:0] pe_13_12_left;
    logic [31:0] pe_13_12_out;
    logic pe_13_12_go;
    logic pe_13_12_clk;
    logic pe_13_12_done;
    logic [31:0] top_13_12_in;
    logic top_13_12_write_en;
    logic top_13_12_clk;
    logic [31:0] top_13_12_out;
    logic top_13_12_done;
    logic [31:0] left_13_12_in;
    logic left_13_12_write_en;
    logic left_13_12_clk;
    logic [31:0] left_13_12_out;
    logic left_13_12_done;
    logic [31:0] pe_13_13_top;
    logic [31:0] pe_13_13_left;
    logic [31:0] pe_13_13_out;
    logic pe_13_13_go;
    logic pe_13_13_clk;
    logic pe_13_13_done;
    logic [31:0] top_13_13_in;
    logic top_13_13_write_en;
    logic top_13_13_clk;
    logic [31:0] top_13_13_out;
    logic top_13_13_done;
    logic [31:0] left_13_13_in;
    logic left_13_13_write_en;
    logic left_13_13_clk;
    logic [31:0] left_13_13_out;
    logic left_13_13_done;
    logic [31:0] pe_13_14_top;
    logic [31:0] pe_13_14_left;
    logic [31:0] pe_13_14_out;
    logic pe_13_14_go;
    logic pe_13_14_clk;
    logic pe_13_14_done;
    logic [31:0] top_13_14_in;
    logic top_13_14_write_en;
    logic top_13_14_clk;
    logic [31:0] top_13_14_out;
    logic top_13_14_done;
    logic [31:0] left_13_14_in;
    logic left_13_14_write_en;
    logic left_13_14_clk;
    logic [31:0] left_13_14_out;
    logic left_13_14_done;
    logic [31:0] pe_13_15_top;
    logic [31:0] pe_13_15_left;
    logic [31:0] pe_13_15_out;
    logic pe_13_15_go;
    logic pe_13_15_clk;
    logic pe_13_15_done;
    logic [31:0] top_13_15_in;
    logic top_13_15_write_en;
    logic top_13_15_clk;
    logic [31:0] top_13_15_out;
    logic top_13_15_done;
    logic [31:0] left_13_15_in;
    logic left_13_15_write_en;
    logic left_13_15_clk;
    logic [31:0] left_13_15_out;
    logic left_13_15_done;
    logic [31:0] pe_14_0_top;
    logic [31:0] pe_14_0_left;
    logic [31:0] pe_14_0_out;
    logic pe_14_0_go;
    logic pe_14_0_clk;
    logic pe_14_0_done;
    logic [31:0] top_14_0_in;
    logic top_14_0_write_en;
    logic top_14_0_clk;
    logic [31:0] top_14_0_out;
    logic top_14_0_done;
    logic [31:0] left_14_0_in;
    logic left_14_0_write_en;
    logic left_14_0_clk;
    logic [31:0] left_14_0_out;
    logic left_14_0_done;
    logic [31:0] pe_14_1_top;
    logic [31:0] pe_14_1_left;
    logic [31:0] pe_14_1_out;
    logic pe_14_1_go;
    logic pe_14_1_clk;
    logic pe_14_1_done;
    logic [31:0] top_14_1_in;
    logic top_14_1_write_en;
    logic top_14_1_clk;
    logic [31:0] top_14_1_out;
    logic top_14_1_done;
    logic [31:0] left_14_1_in;
    logic left_14_1_write_en;
    logic left_14_1_clk;
    logic [31:0] left_14_1_out;
    logic left_14_1_done;
    logic [31:0] pe_14_2_top;
    logic [31:0] pe_14_2_left;
    logic [31:0] pe_14_2_out;
    logic pe_14_2_go;
    logic pe_14_2_clk;
    logic pe_14_2_done;
    logic [31:0] top_14_2_in;
    logic top_14_2_write_en;
    logic top_14_2_clk;
    logic [31:0] top_14_2_out;
    logic top_14_2_done;
    logic [31:0] left_14_2_in;
    logic left_14_2_write_en;
    logic left_14_2_clk;
    logic [31:0] left_14_2_out;
    logic left_14_2_done;
    logic [31:0] pe_14_3_top;
    logic [31:0] pe_14_3_left;
    logic [31:0] pe_14_3_out;
    logic pe_14_3_go;
    logic pe_14_3_clk;
    logic pe_14_3_done;
    logic [31:0] top_14_3_in;
    logic top_14_3_write_en;
    logic top_14_3_clk;
    logic [31:0] top_14_3_out;
    logic top_14_3_done;
    logic [31:0] left_14_3_in;
    logic left_14_3_write_en;
    logic left_14_3_clk;
    logic [31:0] left_14_3_out;
    logic left_14_3_done;
    logic [31:0] pe_14_4_top;
    logic [31:0] pe_14_4_left;
    logic [31:0] pe_14_4_out;
    logic pe_14_4_go;
    logic pe_14_4_clk;
    logic pe_14_4_done;
    logic [31:0] top_14_4_in;
    logic top_14_4_write_en;
    logic top_14_4_clk;
    logic [31:0] top_14_4_out;
    logic top_14_4_done;
    logic [31:0] left_14_4_in;
    logic left_14_4_write_en;
    logic left_14_4_clk;
    logic [31:0] left_14_4_out;
    logic left_14_4_done;
    logic [31:0] pe_14_5_top;
    logic [31:0] pe_14_5_left;
    logic [31:0] pe_14_5_out;
    logic pe_14_5_go;
    logic pe_14_5_clk;
    logic pe_14_5_done;
    logic [31:0] top_14_5_in;
    logic top_14_5_write_en;
    logic top_14_5_clk;
    logic [31:0] top_14_5_out;
    logic top_14_5_done;
    logic [31:0] left_14_5_in;
    logic left_14_5_write_en;
    logic left_14_5_clk;
    logic [31:0] left_14_5_out;
    logic left_14_5_done;
    logic [31:0] pe_14_6_top;
    logic [31:0] pe_14_6_left;
    logic [31:0] pe_14_6_out;
    logic pe_14_6_go;
    logic pe_14_6_clk;
    logic pe_14_6_done;
    logic [31:0] top_14_6_in;
    logic top_14_6_write_en;
    logic top_14_6_clk;
    logic [31:0] top_14_6_out;
    logic top_14_6_done;
    logic [31:0] left_14_6_in;
    logic left_14_6_write_en;
    logic left_14_6_clk;
    logic [31:0] left_14_6_out;
    logic left_14_6_done;
    logic [31:0] pe_14_7_top;
    logic [31:0] pe_14_7_left;
    logic [31:0] pe_14_7_out;
    logic pe_14_7_go;
    logic pe_14_7_clk;
    logic pe_14_7_done;
    logic [31:0] top_14_7_in;
    logic top_14_7_write_en;
    logic top_14_7_clk;
    logic [31:0] top_14_7_out;
    logic top_14_7_done;
    logic [31:0] left_14_7_in;
    logic left_14_7_write_en;
    logic left_14_7_clk;
    logic [31:0] left_14_7_out;
    logic left_14_7_done;
    logic [31:0] pe_14_8_top;
    logic [31:0] pe_14_8_left;
    logic [31:0] pe_14_8_out;
    logic pe_14_8_go;
    logic pe_14_8_clk;
    logic pe_14_8_done;
    logic [31:0] top_14_8_in;
    logic top_14_8_write_en;
    logic top_14_8_clk;
    logic [31:0] top_14_8_out;
    logic top_14_8_done;
    logic [31:0] left_14_8_in;
    logic left_14_8_write_en;
    logic left_14_8_clk;
    logic [31:0] left_14_8_out;
    logic left_14_8_done;
    logic [31:0] pe_14_9_top;
    logic [31:0] pe_14_9_left;
    logic [31:0] pe_14_9_out;
    logic pe_14_9_go;
    logic pe_14_9_clk;
    logic pe_14_9_done;
    logic [31:0] top_14_9_in;
    logic top_14_9_write_en;
    logic top_14_9_clk;
    logic [31:0] top_14_9_out;
    logic top_14_9_done;
    logic [31:0] left_14_9_in;
    logic left_14_9_write_en;
    logic left_14_9_clk;
    logic [31:0] left_14_9_out;
    logic left_14_9_done;
    logic [31:0] pe_14_10_top;
    logic [31:0] pe_14_10_left;
    logic [31:0] pe_14_10_out;
    logic pe_14_10_go;
    logic pe_14_10_clk;
    logic pe_14_10_done;
    logic [31:0] top_14_10_in;
    logic top_14_10_write_en;
    logic top_14_10_clk;
    logic [31:0] top_14_10_out;
    logic top_14_10_done;
    logic [31:0] left_14_10_in;
    logic left_14_10_write_en;
    logic left_14_10_clk;
    logic [31:0] left_14_10_out;
    logic left_14_10_done;
    logic [31:0] pe_14_11_top;
    logic [31:0] pe_14_11_left;
    logic [31:0] pe_14_11_out;
    logic pe_14_11_go;
    logic pe_14_11_clk;
    logic pe_14_11_done;
    logic [31:0] top_14_11_in;
    logic top_14_11_write_en;
    logic top_14_11_clk;
    logic [31:0] top_14_11_out;
    logic top_14_11_done;
    logic [31:0] left_14_11_in;
    logic left_14_11_write_en;
    logic left_14_11_clk;
    logic [31:0] left_14_11_out;
    logic left_14_11_done;
    logic [31:0] pe_14_12_top;
    logic [31:0] pe_14_12_left;
    logic [31:0] pe_14_12_out;
    logic pe_14_12_go;
    logic pe_14_12_clk;
    logic pe_14_12_done;
    logic [31:0] top_14_12_in;
    logic top_14_12_write_en;
    logic top_14_12_clk;
    logic [31:0] top_14_12_out;
    logic top_14_12_done;
    logic [31:0] left_14_12_in;
    logic left_14_12_write_en;
    logic left_14_12_clk;
    logic [31:0] left_14_12_out;
    logic left_14_12_done;
    logic [31:0] pe_14_13_top;
    logic [31:0] pe_14_13_left;
    logic [31:0] pe_14_13_out;
    logic pe_14_13_go;
    logic pe_14_13_clk;
    logic pe_14_13_done;
    logic [31:0] top_14_13_in;
    logic top_14_13_write_en;
    logic top_14_13_clk;
    logic [31:0] top_14_13_out;
    logic top_14_13_done;
    logic [31:0] left_14_13_in;
    logic left_14_13_write_en;
    logic left_14_13_clk;
    logic [31:0] left_14_13_out;
    logic left_14_13_done;
    logic [31:0] pe_14_14_top;
    logic [31:0] pe_14_14_left;
    logic [31:0] pe_14_14_out;
    logic pe_14_14_go;
    logic pe_14_14_clk;
    logic pe_14_14_done;
    logic [31:0] top_14_14_in;
    logic top_14_14_write_en;
    logic top_14_14_clk;
    logic [31:0] top_14_14_out;
    logic top_14_14_done;
    logic [31:0] left_14_14_in;
    logic left_14_14_write_en;
    logic left_14_14_clk;
    logic [31:0] left_14_14_out;
    logic left_14_14_done;
    logic [31:0] pe_14_15_top;
    logic [31:0] pe_14_15_left;
    logic [31:0] pe_14_15_out;
    logic pe_14_15_go;
    logic pe_14_15_clk;
    logic pe_14_15_done;
    logic [31:0] top_14_15_in;
    logic top_14_15_write_en;
    logic top_14_15_clk;
    logic [31:0] top_14_15_out;
    logic top_14_15_done;
    logic [31:0] left_14_15_in;
    logic left_14_15_write_en;
    logic left_14_15_clk;
    logic [31:0] left_14_15_out;
    logic left_14_15_done;
    logic [31:0] pe_15_0_top;
    logic [31:0] pe_15_0_left;
    logic [31:0] pe_15_0_out;
    logic pe_15_0_go;
    logic pe_15_0_clk;
    logic pe_15_0_done;
    logic [31:0] top_15_0_in;
    logic top_15_0_write_en;
    logic top_15_0_clk;
    logic [31:0] top_15_0_out;
    logic top_15_0_done;
    logic [31:0] left_15_0_in;
    logic left_15_0_write_en;
    logic left_15_0_clk;
    logic [31:0] left_15_0_out;
    logic left_15_0_done;
    logic [31:0] pe_15_1_top;
    logic [31:0] pe_15_1_left;
    logic [31:0] pe_15_1_out;
    logic pe_15_1_go;
    logic pe_15_1_clk;
    logic pe_15_1_done;
    logic [31:0] top_15_1_in;
    logic top_15_1_write_en;
    logic top_15_1_clk;
    logic [31:0] top_15_1_out;
    logic top_15_1_done;
    logic [31:0] left_15_1_in;
    logic left_15_1_write_en;
    logic left_15_1_clk;
    logic [31:0] left_15_1_out;
    logic left_15_1_done;
    logic [31:0] pe_15_2_top;
    logic [31:0] pe_15_2_left;
    logic [31:0] pe_15_2_out;
    logic pe_15_2_go;
    logic pe_15_2_clk;
    logic pe_15_2_done;
    logic [31:0] top_15_2_in;
    logic top_15_2_write_en;
    logic top_15_2_clk;
    logic [31:0] top_15_2_out;
    logic top_15_2_done;
    logic [31:0] left_15_2_in;
    logic left_15_2_write_en;
    logic left_15_2_clk;
    logic [31:0] left_15_2_out;
    logic left_15_2_done;
    logic [31:0] pe_15_3_top;
    logic [31:0] pe_15_3_left;
    logic [31:0] pe_15_3_out;
    logic pe_15_3_go;
    logic pe_15_3_clk;
    logic pe_15_3_done;
    logic [31:0] top_15_3_in;
    logic top_15_3_write_en;
    logic top_15_3_clk;
    logic [31:0] top_15_3_out;
    logic top_15_3_done;
    logic [31:0] left_15_3_in;
    logic left_15_3_write_en;
    logic left_15_3_clk;
    logic [31:0] left_15_3_out;
    logic left_15_3_done;
    logic [31:0] pe_15_4_top;
    logic [31:0] pe_15_4_left;
    logic [31:0] pe_15_4_out;
    logic pe_15_4_go;
    logic pe_15_4_clk;
    logic pe_15_4_done;
    logic [31:0] top_15_4_in;
    logic top_15_4_write_en;
    logic top_15_4_clk;
    logic [31:0] top_15_4_out;
    logic top_15_4_done;
    logic [31:0] left_15_4_in;
    logic left_15_4_write_en;
    logic left_15_4_clk;
    logic [31:0] left_15_4_out;
    logic left_15_4_done;
    logic [31:0] pe_15_5_top;
    logic [31:0] pe_15_5_left;
    logic [31:0] pe_15_5_out;
    logic pe_15_5_go;
    logic pe_15_5_clk;
    logic pe_15_5_done;
    logic [31:0] top_15_5_in;
    logic top_15_5_write_en;
    logic top_15_5_clk;
    logic [31:0] top_15_5_out;
    logic top_15_5_done;
    logic [31:0] left_15_5_in;
    logic left_15_5_write_en;
    logic left_15_5_clk;
    logic [31:0] left_15_5_out;
    logic left_15_5_done;
    logic [31:0] pe_15_6_top;
    logic [31:0] pe_15_6_left;
    logic [31:0] pe_15_6_out;
    logic pe_15_6_go;
    logic pe_15_6_clk;
    logic pe_15_6_done;
    logic [31:0] top_15_6_in;
    logic top_15_6_write_en;
    logic top_15_6_clk;
    logic [31:0] top_15_6_out;
    logic top_15_6_done;
    logic [31:0] left_15_6_in;
    logic left_15_6_write_en;
    logic left_15_6_clk;
    logic [31:0] left_15_6_out;
    logic left_15_6_done;
    logic [31:0] pe_15_7_top;
    logic [31:0] pe_15_7_left;
    logic [31:0] pe_15_7_out;
    logic pe_15_7_go;
    logic pe_15_7_clk;
    logic pe_15_7_done;
    logic [31:0] top_15_7_in;
    logic top_15_7_write_en;
    logic top_15_7_clk;
    logic [31:0] top_15_7_out;
    logic top_15_7_done;
    logic [31:0] left_15_7_in;
    logic left_15_7_write_en;
    logic left_15_7_clk;
    logic [31:0] left_15_7_out;
    logic left_15_7_done;
    logic [31:0] pe_15_8_top;
    logic [31:0] pe_15_8_left;
    logic [31:0] pe_15_8_out;
    logic pe_15_8_go;
    logic pe_15_8_clk;
    logic pe_15_8_done;
    logic [31:0] top_15_8_in;
    logic top_15_8_write_en;
    logic top_15_8_clk;
    logic [31:0] top_15_8_out;
    logic top_15_8_done;
    logic [31:0] left_15_8_in;
    logic left_15_8_write_en;
    logic left_15_8_clk;
    logic [31:0] left_15_8_out;
    logic left_15_8_done;
    logic [31:0] pe_15_9_top;
    logic [31:0] pe_15_9_left;
    logic [31:0] pe_15_9_out;
    logic pe_15_9_go;
    logic pe_15_9_clk;
    logic pe_15_9_done;
    logic [31:0] top_15_9_in;
    logic top_15_9_write_en;
    logic top_15_9_clk;
    logic [31:0] top_15_9_out;
    logic top_15_9_done;
    logic [31:0] left_15_9_in;
    logic left_15_9_write_en;
    logic left_15_9_clk;
    logic [31:0] left_15_9_out;
    logic left_15_9_done;
    logic [31:0] pe_15_10_top;
    logic [31:0] pe_15_10_left;
    logic [31:0] pe_15_10_out;
    logic pe_15_10_go;
    logic pe_15_10_clk;
    logic pe_15_10_done;
    logic [31:0] top_15_10_in;
    logic top_15_10_write_en;
    logic top_15_10_clk;
    logic [31:0] top_15_10_out;
    logic top_15_10_done;
    logic [31:0] left_15_10_in;
    logic left_15_10_write_en;
    logic left_15_10_clk;
    logic [31:0] left_15_10_out;
    logic left_15_10_done;
    logic [31:0] pe_15_11_top;
    logic [31:0] pe_15_11_left;
    logic [31:0] pe_15_11_out;
    logic pe_15_11_go;
    logic pe_15_11_clk;
    logic pe_15_11_done;
    logic [31:0] top_15_11_in;
    logic top_15_11_write_en;
    logic top_15_11_clk;
    logic [31:0] top_15_11_out;
    logic top_15_11_done;
    logic [31:0] left_15_11_in;
    logic left_15_11_write_en;
    logic left_15_11_clk;
    logic [31:0] left_15_11_out;
    logic left_15_11_done;
    logic [31:0] pe_15_12_top;
    logic [31:0] pe_15_12_left;
    logic [31:0] pe_15_12_out;
    logic pe_15_12_go;
    logic pe_15_12_clk;
    logic pe_15_12_done;
    logic [31:0] top_15_12_in;
    logic top_15_12_write_en;
    logic top_15_12_clk;
    logic [31:0] top_15_12_out;
    logic top_15_12_done;
    logic [31:0] left_15_12_in;
    logic left_15_12_write_en;
    logic left_15_12_clk;
    logic [31:0] left_15_12_out;
    logic left_15_12_done;
    logic [31:0] pe_15_13_top;
    logic [31:0] pe_15_13_left;
    logic [31:0] pe_15_13_out;
    logic pe_15_13_go;
    logic pe_15_13_clk;
    logic pe_15_13_done;
    logic [31:0] top_15_13_in;
    logic top_15_13_write_en;
    logic top_15_13_clk;
    logic [31:0] top_15_13_out;
    logic top_15_13_done;
    logic [31:0] left_15_13_in;
    logic left_15_13_write_en;
    logic left_15_13_clk;
    logic [31:0] left_15_13_out;
    logic left_15_13_done;
    logic [31:0] pe_15_14_top;
    logic [31:0] pe_15_14_left;
    logic [31:0] pe_15_14_out;
    logic pe_15_14_go;
    logic pe_15_14_clk;
    logic pe_15_14_done;
    logic [31:0] top_15_14_in;
    logic top_15_14_write_en;
    logic top_15_14_clk;
    logic [31:0] top_15_14_out;
    logic top_15_14_done;
    logic [31:0] left_15_14_in;
    logic left_15_14_write_en;
    logic left_15_14_clk;
    logic [31:0] left_15_14_out;
    logic left_15_14_done;
    logic [31:0] pe_15_15_top;
    logic [31:0] pe_15_15_left;
    logic [31:0] pe_15_15_out;
    logic pe_15_15_go;
    logic pe_15_15_clk;
    logic pe_15_15_done;
    logic [31:0] top_15_15_in;
    logic top_15_15_write_en;
    logic top_15_15_clk;
    logic [31:0] top_15_15_out;
    logic top_15_15_done;
    logic [31:0] left_15_15_in;
    logic left_15_15_write_en;
    logic left_15_15_clk;
    logic [31:0] left_15_15_out;
    logic left_15_15_done;
    logic fsm_in;
    logic fsm_write_en;
    logic fsm_clk;
    logic fsm_out;
    logic fsm_done;
    logic incr_left;
    logic incr_right;
    logic incr_out;
    logic fsm0_in;
    logic fsm0_write_en;
    logic fsm0_clk;
    logic fsm0_out;
    logic fsm0_done;
    logic incr0_left;
    logic incr0_right;
    logic incr0_out;
    logic fsm1_in;
    logic fsm1_write_en;
    logic fsm1_clk;
    logic fsm1_out;
    logic fsm1_done;
    logic incr1_left;
    logic incr1_right;
    logic incr1_out;
    logic [2:0] fsm2_in;
    logic fsm2_write_en;
    logic fsm2_clk;
    logic [2:0] fsm2_out;
    logic fsm2_done;
    logic [2:0] incr2_left;
    logic [2:0] incr2_right;
    logic [2:0] incr2_out;
    logic fsm3_in;
    logic fsm3_write_en;
    logic fsm3_clk;
    logic fsm3_out;
    logic fsm3_done;
    logic incr3_left;
    logic incr3_right;
    logic incr3_out;
    logic [2:0] fsm4_in;
    logic fsm4_write_en;
    logic fsm4_clk;
    logic [2:0] fsm4_out;
    logic fsm4_done;
    logic [2:0] incr4_left;
    logic [2:0] incr4_right;
    logic [2:0] incr4_out;
    logic fsm5_in;
    logic fsm5_write_en;
    logic fsm5_clk;
    logic fsm5_out;
    logic fsm5_done;
    logic incr5_left;
    logic incr5_right;
    logic incr5_out;
    logic [2:0] fsm6_in;
    logic fsm6_write_en;
    logic fsm6_clk;
    logic [2:0] fsm6_out;
    logic fsm6_done;
    logic [2:0] incr6_left;
    logic [2:0] incr6_right;
    logic [2:0] incr6_out;
    logic fsm7_in;
    logic fsm7_write_en;
    logic fsm7_clk;
    logic fsm7_out;
    logic fsm7_done;
    logic incr7_left;
    logic incr7_right;
    logic incr7_out;
    logic [2:0] fsm8_in;
    logic fsm8_write_en;
    logic fsm8_clk;
    logic [2:0] fsm8_out;
    logic fsm8_done;
    logic [2:0] incr8_left;
    logic [2:0] incr8_right;
    logic [2:0] incr8_out;
    logic fsm9_in;
    logic fsm9_write_en;
    logic fsm9_clk;
    logic fsm9_out;
    logic fsm9_done;
    logic incr9_left;
    logic incr9_right;
    logic incr9_out;
    logic [2:0] fsm10_in;
    logic fsm10_write_en;
    logic fsm10_clk;
    logic [2:0] fsm10_out;
    logic fsm10_done;
    logic [2:0] incr10_left;
    logic [2:0] incr10_right;
    logic [2:0] incr10_out;
    logic fsm11_in;
    logic fsm11_write_en;
    logic fsm11_clk;
    logic fsm11_out;
    logic fsm11_done;
    logic incr11_left;
    logic incr11_right;
    logic incr11_out;
    logic [2:0] fsm12_in;
    logic fsm12_write_en;
    logic fsm12_clk;
    logic [2:0] fsm12_out;
    logic fsm12_done;
    logic [2:0] incr12_left;
    logic [2:0] incr12_right;
    logic [2:0] incr12_out;
    logic fsm13_in;
    logic fsm13_write_en;
    logic fsm13_clk;
    logic fsm13_out;
    logic fsm13_done;
    logic incr13_left;
    logic incr13_right;
    logic incr13_out;
    logic [2:0] fsm14_in;
    logic fsm14_write_en;
    logic fsm14_clk;
    logic [2:0] fsm14_out;
    logic fsm14_done;
    logic [2:0] incr14_left;
    logic [2:0] incr14_right;
    logic [2:0] incr14_out;
    logic fsm15_in;
    logic fsm15_write_en;
    logic fsm15_clk;
    logic fsm15_out;
    logic fsm15_done;
    logic incr15_left;
    logic incr15_right;
    logic incr15_out;
    logic [2:0] fsm16_in;
    logic fsm16_write_en;
    logic fsm16_clk;
    logic [2:0] fsm16_out;
    logic fsm16_done;
    logic [2:0] incr16_left;
    logic [2:0] incr16_right;
    logic [2:0] incr16_out;
    logic fsm17_in;
    logic fsm17_write_en;
    logic fsm17_clk;
    logic fsm17_out;
    logic fsm17_done;
    logic incr17_left;
    logic incr17_right;
    logic incr17_out;
    logic [2:0] fsm18_in;
    logic fsm18_write_en;
    logic fsm18_clk;
    logic [2:0] fsm18_out;
    logic fsm18_done;
    logic [2:0] incr18_left;
    logic [2:0] incr18_right;
    logic [2:0] incr18_out;
    logic fsm19_in;
    logic fsm19_write_en;
    logic fsm19_clk;
    logic fsm19_out;
    logic fsm19_done;
    logic incr19_left;
    logic incr19_right;
    logic incr19_out;
    logic [2:0] fsm20_in;
    logic fsm20_write_en;
    logic fsm20_clk;
    logic [2:0] fsm20_out;
    logic fsm20_done;
    logic [2:0] incr20_left;
    logic [2:0] incr20_right;
    logic [2:0] incr20_out;
    logic fsm21_in;
    logic fsm21_write_en;
    logic fsm21_clk;
    logic fsm21_out;
    logic fsm21_done;
    logic incr21_left;
    logic incr21_right;
    logic incr21_out;
    logic [2:0] fsm22_in;
    logic fsm22_write_en;
    logic fsm22_clk;
    logic [2:0] fsm22_out;
    logic fsm22_done;
    logic [2:0] incr22_left;
    logic [2:0] incr22_right;
    logic [2:0] incr22_out;
    logic fsm23_in;
    logic fsm23_write_en;
    logic fsm23_clk;
    logic fsm23_out;
    logic fsm23_done;
    logic incr23_left;
    logic incr23_right;
    logic incr23_out;
    logic [2:0] fsm24_in;
    logic fsm24_write_en;
    logic fsm24_clk;
    logic [2:0] fsm24_out;
    logic fsm24_done;
    logic [2:0] incr24_left;
    logic [2:0] incr24_right;
    logic [2:0] incr24_out;
    logic fsm25_in;
    logic fsm25_write_en;
    logic fsm25_clk;
    logic fsm25_out;
    logic fsm25_done;
    logic incr25_left;
    logic incr25_right;
    logic incr25_out;
    logic [2:0] fsm26_in;
    logic fsm26_write_en;
    logic fsm26_clk;
    logic [2:0] fsm26_out;
    logic fsm26_done;
    logic [2:0] incr26_left;
    logic [2:0] incr26_right;
    logic [2:0] incr26_out;
    logic fsm27_in;
    logic fsm27_write_en;
    logic fsm27_clk;
    logic fsm27_out;
    logic fsm27_done;
    logic incr27_left;
    logic incr27_right;
    logic incr27_out;
    logic [2:0] fsm28_in;
    logic fsm28_write_en;
    logic fsm28_clk;
    logic [2:0] fsm28_out;
    logic fsm28_done;
    logic [2:0] incr28_left;
    logic [2:0] incr28_right;
    logic [2:0] incr28_out;
    logic fsm29_in;
    logic fsm29_write_en;
    logic fsm29_clk;
    logic fsm29_out;
    logic fsm29_done;
    logic incr29_left;
    logic incr29_right;
    logic incr29_out;
    logic [2:0] fsm30_in;
    logic fsm30_write_en;
    logic fsm30_clk;
    logic [2:0] fsm30_out;
    logic fsm30_done;
    logic [2:0] incr30_left;
    logic [2:0] incr30_right;
    logic [2:0] incr30_out;
    logic fsm31_in;
    logic fsm31_write_en;
    logic fsm31_clk;
    logic fsm31_out;
    logic fsm31_done;
    logic incr31_left;
    logic incr31_right;
    logic incr31_out;
    logic [2:0] fsm32_in;
    logic fsm32_write_en;
    logic fsm32_clk;
    logic [2:0] fsm32_out;
    logic fsm32_done;
    logic [2:0] incr32_left;
    logic [2:0] incr32_right;
    logic [2:0] incr32_out;
    logic fsm33_in;
    logic fsm33_write_en;
    logic fsm33_clk;
    logic fsm33_out;
    logic fsm33_done;
    logic incr33_left;
    logic incr33_right;
    logic incr33_out;
    logic [2:0] fsm34_in;
    logic fsm34_write_en;
    logic fsm34_clk;
    logic [2:0] fsm34_out;
    logic fsm34_done;
    logic [2:0] incr34_left;
    logic [2:0] incr34_right;
    logic [2:0] incr34_out;
    logic fsm35_in;
    logic fsm35_write_en;
    logic fsm35_clk;
    logic fsm35_out;
    logic fsm35_done;
    logic incr35_left;
    logic incr35_right;
    logic incr35_out;
    logic [2:0] fsm36_in;
    logic fsm36_write_en;
    logic fsm36_clk;
    logic [2:0] fsm36_out;
    logic fsm36_done;
    logic [2:0] incr36_left;
    logic [2:0] incr36_right;
    logic [2:0] incr36_out;
    logic fsm37_in;
    logic fsm37_write_en;
    logic fsm37_clk;
    logic fsm37_out;
    logic fsm37_done;
    logic incr37_left;
    logic incr37_right;
    logic incr37_out;
    logic [2:0] fsm38_in;
    logic fsm38_write_en;
    logic fsm38_clk;
    logic [2:0] fsm38_out;
    logic fsm38_done;
    logic [2:0] incr38_left;
    logic [2:0] incr38_right;
    logic [2:0] incr38_out;
    logic fsm39_in;
    logic fsm39_write_en;
    logic fsm39_clk;
    logic fsm39_out;
    logic fsm39_done;
    logic incr39_left;
    logic incr39_right;
    logic incr39_out;
    logic [2:0] fsm40_in;
    logic fsm40_write_en;
    logic fsm40_clk;
    logic [2:0] fsm40_out;
    logic fsm40_done;
    logic [2:0] incr40_left;
    logic [2:0] incr40_right;
    logic [2:0] incr40_out;
    logic fsm41_in;
    logic fsm41_write_en;
    logic fsm41_clk;
    logic fsm41_out;
    logic fsm41_done;
    logic incr41_left;
    logic incr41_right;
    logic incr41_out;
    logic [2:0] fsm42_in;
    logic fsm42_write_en;
    logic fsm42_clk;
    logic [2:0] fsm42_out;
    logic fsm42_done;
    logic [2:0] incr42_left;
    logic [2:0] incr42_right;
    logic [2:0] incr42_out;
    logic fsm43_in;
    logic fsm43_write_en;
    logic fsm43_clk;
    logic fsm43_out;
    logic fsm43_done;
    logic incr43_left;
    logic incr43_right;
    logic incr43_out;
    logic [2:0] fsm44_in;
    logic fsm44_write_en;
    logic fsm44_clk;
    logic [2:0] fsm44_out;
    logic fsm44_done;
    logic [2:0] incr44_left;
    logic [2:0] incr44_right;
    logic [2:0] incr44_out;
    logic fsm45_in;
    logic fsm45_write_en;
    logic fsm45_clk;
    logic fsm45_out;
    logic fsm45_done;
    logic incr45_left;
    logic incr45_right;
    logic incr45_out;
    logic [2:0] fsm46_in;
    logic fsm46_write_en;
    logic fsm46_clk;
    logic [2:0] fsm46_out;
    logic fsm46_done;
    logic [2:0] incr46_left;
    logic [2:0] incr46_right;
    logic [2:0] incr46_out;
    logic fsm47_in;
    logic fsm47_write_en;
    logic fsm47_clk;
    logic fsm47_out;
    logic fsm47_done;
    logic incr47_left;
    logic incr47_right;
    logic incr47_out;
    logic [2:0] fsm48_in;
    logic fsm48_write_en;
    logic fsm48_clk;
    logic [2:0] fsm48_out;
    logic fsm48_done;
    logic [2:0] incr48_left;
    logic [2:0] incr48_right;
    logic [2:0] incr48_out;
    logic fsm49_in;
    logic fsm49_write_en;
    logic fsm49_clk;
    logic fsm49_out;
    logic fsm49_done;
    logic incr49_left;
    logic incr49_right;
    logic incr49_out;
    logic [2:0] fsm50_in;
    logic fsm50_write_en;
    logic fsm50_clk;
    logic [2:0] fsm50_out;
    logic fsm50_done;
    logic [2:0] incr50_left;
    logic [2:0] incr50_right;
    logic [2:0] incr50_out;
    logic fsm51_in;
    logic fsm51_write_en;
    logic fsm51_clk;
    logic fsm51_out;
    logic fsm51_done;
    logic incr51_left;
    logic incr51_right;
    logic incr51_out;
    logic [2:0] fsm52_in;
    logic fsm52_write_en;
    logic fsm52_clk;
    logic [2:0] fsm52_out;
    logic fsm52_done;
    logic [2:0] incr52_left;
    logic [2:0] incr52_right;
    logic [2:0] incr52_out;
    logic fsm53_in;
    logic fsm53_write_en;
    logic fsm53_clk;
    logic fsm53_out;
    logic fsm53_done;
    logic incr53_left;
    logic incr53_right;
    logic incr53_out;
    logic [2:0] fsm54_in;
    logic fsm54_write_en;
    logic fsm54_clk;
    logic [2:0] fsm54_out;
    logic fsm54_done;
    logic [2:0] incr54_left;
    logic [2:0] incr54_right;
    logic [2:0] incr54_out;
    logic fsm55_in;
    logic fsm55_write_en;
    logic fsm55_clk;
    logic fsm55_out;
    logic fsm55_done;
    logic incr55_left;
    logic incr55_right;
    logic incr55_out;
    logic [2:0] fsm56_in;
    logic fsm56_write_en;
    logic fsm56_clk;
    logic [2:0] fsm56_out;
    logic fsm56_done;
    logic [2:0] incr56_left;
    logic [2:0] incr56_right;
    logic [2:0] incr56_out;
    logic fsm57_in;
    logic fsm57_write_en;
    logic fsm57_clk;
    logic fsm57_out;
    logic fsm57_done;
    logic incr57_left;
    logic incr57_right;
    logic incr57_out;
    logic [2:0] fsm58_in;
    logic fsm58_write_en;
    logic fsm58_clk;
    logic [2:0] fsm58_out;
    logic fsm58_done;
    logic [2:0] incr58_left;
    logic [2:0] incr58_right;
    logic [2:0] incr58_out;
    logic fsm59_in;
    logic fsm59_write_en;
    logic fsm59_clk;
    logic fsm59_out;
    logic fsm59_done;
    logic incr59_left;
    logic incr59_right;
    logic incr59_out;
    logic [2:0] fsm60_in;
    logic fsm60_write_en;
    logic fsm60_clk;
    logic [2:0] fsm60_out;
    logic fsm60_done;
    logic [2:0] incr60_left;
    logic [2:0] incr60_right;
    logic [2:0] incr60_out;
    logic fsm61_in;
    logic fsm61_write_en;
    logic fsm61_clk;
    logic fsm61_out;
    logic fsm61_done;
    logic incr61_left;
    logic incr61_right;
    logic incr61_out;
    logic [2:0] fsm62_in;
    logic fsm62_write_en;
    logic fsm62_clk;
    logic [2:0] fsm62_out;
    logic fsm62_done;
    logic [2:0] incr62_left;
    logic [2:0] incr62_right;
    logic [2:0] incr62_out;
    logic fsm63_in;
    logic fsm63_write_en;
    logic fsm63_clk;
    logic fsm63_out;
    logic fsm63_done;
    logic incr63_left;
    logic incr63_right;
    logic incr63_out;
    logic [2:0] fsm64_in;
    logic fsm64_write_en;
    logic fsm64_clk;
    logic [2:0] fsm64_out;
    logic fsm64_done;
    logic [2:0] incr64_left;
    logic [2:0] incr64_right;
    logic [2:0] incr64_out;
    logic fsm65_in;
    logic fsm65_write_en;
    logic fsm65_clk;
    logic fsm65_out;
    logic fsm65_done;
    logic incr65_left;
    logic incr65_right;
    logic incr65_out;
    logic [2:0] fsm66_in;
    logic fsm66_write_en;
    logic fsm66_clk;
    logic [2:0] fsm66_out;
    logic fsm66_done;
    logic [2:0] incr66_left;
    logic [2:0] incr66_right;
    logic [2:0] incr66_out;
    logic fsm67_in;
    logic fsm67_write_en;
    logic fsm67_clk;
    logic fsm67_out;
    logic fsm67_done;
    logic incr67_left;
    logic incr67_right;
    logic incr67_out;
    logic [2:0] fsm68_in;
    logic fsm68_write_en;
    logic fsm68_clk;
    logic [2:0] fsm68_out;
    logic fsm68_done;
    logic [2:0] incr68_left;
    logic [2:0] incr68_right;
    logic [2:0] incr68_out;
    logic fsm69_in;
    logic fsm69_write_en;
    logic fsm69_clk;
    logic fsm69_out;
    logic fsm69_done;
    logic incr69_left;
    logic incr69_right;
    logic incr69_out;
    logic [2:0] fsm70_in;
    logic fsm70_write_en;
    logic fsm70_clk;
    logic [2:0] fsm70_out;
    logic fsm70_done;
    logic [2:0] incr70_left;
    logic [2:0] incr70_right;
    logic [2:0] incr70_out;
    logic fsm71_in;
    logic fsm71_write_en;
    logic fsm71_clk;
    logic fsm71_out;
    logic fsm71_done;
    logic incr71_left;
    logic incr71_right;
    logic incr71_out;
    logic [2:0] fsm72_in;
    logic fsm72_write_en;
    logic fsm72_clk;
    logic [2:0] fsm72_out;
    logic fsm72_done;
    logic [2:0] incr72_left;
    logic [2:0] incr72_right;
    logic [2:0] incr72_out;
    logic fsm73_in;
    logic fsm73_write_en;
    logic fsm73_clk;
    logic fsm73_out;
    logic fsm73_done;
    logic incr73_left;
    logic incr73_right;
    logic incr73_out;
    logic [2:0] fsm74_in;
    logic fsm74_write_en;
    logic fsm74_clk;
    logic [2:0] fsm74_out;
    logic fsm74_done;
    logic [2:0] incr74_left;
    logic [2:0] incr74_right;
    logic [2:0] incr74_out;
    logic fsm75_in;
    logic fsm75_write_en;
    logic fsm75_clk;
    logic fsm75_out;
    logic fsm75_done;
    logic incr75_left;
    logic incr75_right;
    logic incr75_out;
    logic [2:0] fsm76_in;
    logic fsm76_write_en;
    logic fsm76_clk;
    logic [2:0] fsm76_out;
    logic fsm76_done;
    logic [2:0] incr76_left;
    logic [2:0] incr76_right;
    logic [2:0] incr76_out;
    logic fsm77_in;
    logic fsm77_write_en;
    logic fsm77_clk;
    logic fsm77_out;
    logic fsm77_done;
    logic incr77_left;
    logic incr77_right;
    logic incr77_out;
    logic [2:0] fsm78_in;
    logic fsm78_write_en;
    logic fsm78_clk;
    logic [2:0] fsm78_out;
    logic fsm78_done;
    logic [2:0] incr78_left;
    logic [2:0] incr78_right;
    logic [2:0] incr78_out;
    logic fsm79_in;
    logic fsm79_write_en;
    logic fsm79_clk;
    logic fsm79_out;
    logic fsm79_done;
    logic incr79_left;
    logic incr79_right;
    logic incr79_out;
    logic [2:0] fsm80_in;
    logic fsm80_write_en;
    logic fsm80_clk;
    logic [2:0] fsm80_out;
    logic fsm80_done;
    logic [2:0] incr80_left;
    logic [2:0] incr80_right;
    logic [2:0] incr80_out;
    logic fsm81_in;
    logic fsm81_write_en;
    logic fsm81_clk;
    logic fsm81_out;
    logic fsm81_done;
    logic incr81_left;
    logic incr81_right;
    logic incr81_out;
    logic [2:0] fsm82_in;
    logic fsm82_write_en;
    logic fsm82_clk;
    logic [2:0] fsm82_out;
    logic fsm82_done;
    logic [2:0] incr82_left;
    logic [2:0] incr82_right;
    logic [2:0] incr82_out;
    logic fsm83_in;
    logic fsm83_write_en;
    logic fsm83_clk;
    logic fsm83_out;
    logic fsm83_done;
    logic incr83_left;
    logic incr83_right;
    logic incr83_out;
    logic [2:0] fsm84_in;
    logic fsm84_write_en;
    logic fsm84_clk;
    logic [2:0] fsm84_out;
    logic fsm84_done;
    logic [2:0] incr84_left;
    logic [2:0] incr84_right;
    logic [2:0] incr84_out;
    logic fsm85_in;
    logic fsm85_write_en;
    logic fsm85_clk;
    logic fsm85_out;
    logic fsm85_done;
    logic incr85_left;
    logic incr85_right;
    logic incr85_out;
    logic [2:0] fsm86_in;
    logic fsm86_write_en;
    logic fsm86_clk;
    logic [2:0] fsm86_out;
    logic fsm86_done;
    logic [2:0] incr86_left;
    logic [2:0] incr86_right;
    logic [2:0] incr86_out;
    logic fsm87_in;
    logic fsm87_write_en;
    logic fsm87_clk;
    logic fsm87_out;
    logic fsm87_done;
    logic incr87_left;
    logic incr87_right;
    logic incr87_out;
    logic [2:0] fsm88_in;
    logic fsm88_write_en;
    logic fsm88_clk;
    logic [2:0] fsm88_out;
    logic fsm88_done;
    logic [2:0] incr88_left;
    logic [2:0] incr88_right;
    logic [2:0] incr88_out;
    logic fsm89_in;
    logic fsm89_write_en;
    logic fsm89_clk;
    logic fsm89_out;
    logic fsm89_done;
    logic incr89_left;
    logic incr89_right;
    logic incr89_out;
    logic [2:0] fsm90_in;
    logic fsm90_write_en;
    logic fsm90_clk;
    logic [2:0] fsm90_out;
    logic fsm90_done;
    logic [2:0] incr90_left;
    logic [2:0] incr90_right;
    logic [2:0] incr90_out;
    logic fsm91_in;
    logic fsm91_write_en;
    logic fsm91_clk;
    logic fsm91_out;
    logic fsm91_done;
    logic incr91_left;
    logic incr91_right;
    logic incr91_out;
    logic [9:0] fsm92_in;
    logic fsm92_write_en;
    logic fsm92_clk;
    logic [9:0] fsm92_out;
    logic fsm92_done;
    logic [9:0] incr92_left;
    logic [9:0] incr92_right;
    logic [9:0] incr92_out;
    initial begin
        t0_idx_in = 5'd0;
        t0_idx_write_en = 1'd0;
        t0_idx_clk = 1'd0;
        t0_add_left = 5'd0;
        t0_add_right = 5'd0;
        t1_idx_in = 5'd0;
        t1_idx_write_en = 1'd0;
        t1_idx_clk = 1'd0;
        t1_add_left = 5'd0;
        t1_add_right = 5'd0;
        t2_idx_in = 5'd0;
        t2_idx_write_en = 1'd0;
        t2_idx_clk = 1'd0;
        t2_add_left = 5'd0;
        t2_add_right = 5'd0;
        t3_idx_in = 5'd0;
        t3_idx_write_en = 1'd0;
        t3_idx_clk = 1'd0;
        t3_add_left = 5'd0;
        t3_add_right = 5'd0;
        t4_idx_in = 5'd0;
        t4_idx_write_en = 1'd0;
        t4_idx_clk = 1'd0;
        t4_add_left = 5'd0;
        t4_add_right = 5'd0;
        t5_idx_in = 5'd0;
        t5_idx_write_en = 1'd0;
        t5_idx_clk = 1'd0;
        t5_add_left = 5'd0;
        t5_add_right = 5'd0;
        t6_idx_in = 5'd0;
        t6_idx_write_en = 1'd0;
        t6_idx_clk = 1'd0;
        t6_add_left = 5'd0;
        t6_add_right = 5'd0;
        t7_idx_in = 5'd0;
        t7_idx_write_en = 1'd0;
        t7_idx_clk = 1'd0;
        t7_add_left = 5'd0;
        t7_add_right = 5'd0;
        t8_idx_in = 5'd0;
        t8_idx_write_en = 1'd0;
        t8_idx_clk = 1'd0;
        t8_add_left = 5'd0;
        t8_add_right = 5'd0;
        t9_idx_in = 5'd0;
        t9_idx_write_en = 1'd0;
        t9_idx_clk = 1'd0;
        t9_add_left = 5'd0;
        t9_add_right = 5'd0;
        t10_idx_in = 5'd0;
        t10_idx_write_en = 1'd0;
        t10_idx_clk = 1'd0;
        t10_add_left = 5'd0;
        t10_add_right = 5'd0;
        t11_idx_in = 5'd0;
        t11_idx_write_en = 1'd0;
        t11_idx_clk = 1'd0;
        t11_add_left = 5'd0;
        t11_add_right = 5'd0;
        t12_idx_in = 5'd0;
        t12_idx_write_en = 1'd0;
        t12_idx_clk = 1'd0;
        t12_add_left = 5'd0;
        t12_add_right = 5'd0;
        t13_idx_in = 5'd0;
        t13_idx_write_en = 1'd0;
        t13_idx_clk = 1'd0;
        t13_add_left = 5'd0;
        t13_add_right = 5'd0;
        t14_idx_in = 5'd0;
        t14_idx_write_en = 1'd0;
        t14_idx_clk = 1'd0;
        t14_add_left = 5'd0;
        t14_add_right = 5'd0;
        t15_idx_in = 5'd0;
        t15_idx_write_en = 1'd0;
        t15_idx_clk = 1'd0;
        t15_add_left = 5'd0;
        t15_add_right = 5'd0;
        l0_idx_in = 5'd0;
        l0_idx_write_en = 1'd0;
        l0_idx_clk = 1'd0;
        l0_add_left = 5'd0;
        l0_add_right = 5'd0;
        l1_idx_in = 5'd0;
        l1_idx_write_en = 1'd0;
        l1_idx_clk = 1'd0;
        l1_add_left = 5'd0;
        l1_add_right = 5'd0;
        l2_idx_in = 5'd0;
        l2_idx_write_en = 1'd0;
        l2_idx_clk = 1'd0;
        l2_add_left = 5'd0;
        l2_add_right = 5'd0;
        l3_idx_in = 5'd0;
        l3_idx_write_en = 1'd0;
        l3_idx_clk = 1'd0;
        l3_add_left = 5'd0;
        l3_add_right = 5'd0;
        l4_idx_in = 5'd0;
        l4_idx_write_en = 1'd0;
        l4_idx_clk = 1'd0;
        l4_add_left = 5'd0;
        l4_add_right = 5'd0;
        l5_idx_in = 5'd0;
        l5_idx_write_en = 1'd0;
        l5_idx_clk = 1'd0;
        l5_add_left = 5'd0;
        l5_add_right = 5'd0;
        l6_idx_in = 5'd0;
        l6_idx_write_en = 1'd0;
        l6_idx_clk = 1'd0;
        l6_add_left = 5'd0;
        l6_add_right = 5'd0;
        l7_idx_in = 5'd0;
        l7_idx_write_en = 1'd0;
        l7_idx_clk = 1'd0;
        l7_add_left = 5'd0;
        l7_add_right = 5'd0;
        l8_idx_in = 5'd0;
        l8_idx_write_en = 1'd0;
        l8_idx_clk = 1'd0;
        l8_add_left = 5'd0;
        l8_add_right = 5'd0;
        l9_idx_in = 5'd0;
        l9_idx_write_en = 1'd0;
        l9_idx_clk = 1'd0;
        l9_add_left = 5'd0;
        l9_add_right = 5'd0;
        l10_idx_in = 5'd0;
        l10_idx_write_en = 1'd0;
        l10_idx_clk = 1'd0;
        l10_add_left = 5'd0;
        l10_add_right = 5'd0;
        l11_idx_in = 5'd0;
        l11_idx_write_en = 1'd0;
        l11_idx_clk = 1'd0;
        l11_add_left = 5'd0;
        l11_add_right = 5'd0;
        l12_idx_in = 5'd0;
        l12_idx_write_en = 1'd0;
        l12_idx_clk = 1'd0;
        l12_add_left = 5'd0;
        l12_add_right = 5'd0;
        l13_idx_in = 5'd0;
        l13_idx_write_en = 1'd0;
        l13_idx_clk = 1'd0;
        l13_add_left = 5'd0;
        l13_add_right = 5'd0;
        l14_idx_in = 5'd0;
        l14_idx_write_en = 1'd0;
        l14_idx_clk = 1'd0;
        l14_add_left = 5'd0;
        l14_add_right = 5'd0;
        l15_idx_in = 5'd0;
        l15_idx_write_en = 1'd0;
        l15_idx_clk = 1'd0;
        l15_add_left = 5'd0;
        l15_add_right = 5'd0;
        pe_0_0_top = 32'd0;
        pe_0_0_left = 32'd0;
        pe_0_0_go = 1'd0;
        pe_0_0_clk = 1'd0;
        top_0_0_in = 32'd0;
        top_0_0_write_en = 1'd0;
        top_0_0_clk = 1'd0;
        left_0_0_in = 32'd0;
        left_0_0_write_en = 1'd0;
        left_0_0_clk = 1'd0;
        pe_0_1_top = 32'd0;
        pe_0_1_left = 32'd0;
        pe_0_1_go = 1'd0;
        pe_0_1_clk = 1'd0;
        top_0_1_in = 32'd0;
        top_0_1_write_en = 1'd0;
        top_0_1_clk = 1'd0;
        left_0_1_in = 32'd0;
        left_0_1_write_en = 1'd0;
        left_0_1_clk = 1'd0;
        pe_0_2_top = 32'd0;
        pe_0_2_left = 32'd0;
        pe_0_2_go = 1'd0;
        pe_0_2_clk = 1'd0;
        top_0_2_in = 32'd0;
        top_0_2_write_en = 1'd0;
        top_0_2_clk = 1'd0;
        left_0_2_in = 32'd0;
        left_0_2_write_en = 1'd0;
        left_0_2_clk = 1'd0;
        pe_0_3_top = 32'd0;
        pe_0_3_left = 32'd0;
        pe_0_3_go = 1'd0;
        pe_0_3_clk = 1'd0;
        top_0_3_in = 32'd0;
        top_0_3_write_en = 1'd0;
        top_0_3_clk = 1'd0;
        left_0_3_in = 32'd0;
        left_0_3_write_en = 1'd0;
        left_0_3_clk = 1'd0;
        pe_0_4_top = 32'd0;
        pe_0_4_left = 32'd0;
        pe_0_4_go = 1'd0;
        pe_0_4_clk = 1'd0;
        top_0_4_in = 32'd0;
        top_0_4_write_en = 1'd0;
        top_0_4_clk = 1'd0;
        left_0_4_in = 32'd0;
        left_0_4_write_en = 1'd0;
        left_0_4_clk = 1'd0;
        pe_0_5_top = 32'd0;
        pe_0_5_left = 32'd0;
        pe_0_5_go = 1'd0;
        pe_0_5_clk = 1'd0;
        top_0_5_in = 32'd0;
        top_0_5_write_en = 1'd0;
        top_0_5_clk = 1'd0;
        left_0_5_in = 32'd0;
        left_0_5_write_en = 1'd0;
        left_0_5_clk = 1'd0;
        pe_0_6_top = 32'd0;
        pe_0_6_left = 32'd0;
        pe_0_6_go = 1'd0;
        pe_0_6_clk = 1'd0;
        top_0_6_in = 32'd0;
        top_0_6_write_en = 1'd0;
        top_0_6_clk = 1'd0;
        left_0_6_in = 32'd0;
        left_0_6_write_en = 1'd0;
        left_0_6_clk = 1'd0;
        pe_0_7_top = 32'd0;
        pe_0_7_left = 32'd0;
        pe_0_7_go = 1'd0;
        pe_0_7_clk = 1'd0;
        top_0_7_in = 32'd0;
        top_0_7_write_en = 1'd0;
        top_0_7_clk = 1'd0;
        left_0_7_in = 32'd0;
        left_0_7_write_en = 1'd0;
        left_0_7_clk = 1'd0;
        pe_0_8_top = 32'd0;
        pe_0_8_left = 32'd0;
        pe_0_8_go = 1'd0;
        pe_0_8_clk = 1'd0;
        top_0_8_in = 32'd0;
        top_0_8_write_en = 1'd0;
        top_0_8_clk = 1'd0;
        left_0_8_in = 32'd0;
        left_0_8_write_en = 1'd0;
        left_0_8_clk = 1'd0;
        pe_0_9_top = 32'd0;
        pe_0_9_left = 32'd0;
        pe_0_9_go = 1'd0;
        pe_0_9_clk = 1'd0;
        top_0_9_in = 32'd0;
        top_0_9_write_en = 1'd0;
        top_0_9_clk = 1'd0;
        left_0_9_in = 32'd0;
        left_0_9_write_en = 1'd0;
        left_0_9_clk = 1'd0;
        pe_0_10_top = 32'd0;
        pe_0_10_left = 32'd0;
        pe_0_10_go = 1'd0;
        pe_0_10_clk = 1'd0;
        top_0_10_in = 32'd0;
        top_0_10_write_en = 1'd0;
        top_0_10_clk = 1'd0;
        left_0_10_in = 32'd0;
        left_0_10_write_en = 1'd0;
        left_0_10_clk = 1'd0;
        pe_0_11_top = 32'd0;
        pe_0_11_left = 32'd0;
        pe_0_11_go = 1'd0;
        pe_0_11_clk = 1'd0;
        top_0_11_in = 32'd0;
        top_0_11_write_en = 1'd0;
        top_0_11_clk = 1'd0;
        left_0_11_in = 32'd0;
        left_0_11_write_en = 1'd0;
        left_0_11_clk = 1'd0;
        pe_0_12_top = 32'd0;
        pe_0_12_left = 32'd0;
        pe_0_12_go = 1'd0;
        pe_0_12_clk = 1'd0;
        top_0_12_in = 32'd0;
        top_0_12_write_en = 1'd0;
        top_0_12_clk = 1'd0;
        left_0_12_in = 32'd0;
        left_0_12_write_en = 1'd0;
        left_0_12_clk = 1'd0;
        pe_0_13_top = 32'd0;
        pe_0_13_left = 32'd0;
        pe_0_13_go = 1'd0;
        pe_0_13_clk = 1'd0;
        top_0_13_in = 32'd0;
        top_0_13_write_en = 1'd0;
        top_0_13_clk = 1'd0;
        left_0_13_in = 32'd0;
        left_0_13_write_en = 1'd0;
        left_0_13_clk = 1'd0;
        pe_0_14_top = 32'd0;
        pe_0_14_left = 32'd0;
        pe_0_14_go = 1'd0;
        pe_0_14_clk = 1'd0;
        top_0_14_in = 32'd0;
        top_0_14_write_en = 1'd0;
        top_0_14_clk = 1'd0;
        left_0_14_in = 32'd0;
        left_0_14_write_en = 1'd0;
        left_0_14_clk = 1'd0;
        pe_0_15_top = 32'd0;
        pe_0_15_left = 32'd0;
        pe_0_15_go = 1'd0;
        pe_0_15_clk = 1'd0;
        top_0_15_in = 32'd0;
        top_0_15_write_en = 1'd0;
        top_0_15_clk = 1'd0;
        left_0_15_in = 32'd0;
        left_0_15_write_en = 1'd0;
        left_0_15_clk = 1'd0;
        pe_1_0_top = 32'd0;
        pe_1_0_left = 32'd0;
        pe_1_0_go = 1'd0;
        pe_1_0_clk = 1'd0;
        top_1_0_in = 32'd0;
        top_1_0_write_en = 1'd0;
        top_1_0_clk = 1'd0;
        left_1_0_in = 32'd0;
        left_1_0_write_en = 1'd0;
        left_1_0_clk = 1'd0;
        pe_1_1_top = 32'd0;
        pe_1_1_left = 32'd0;
        pe_1_1_go = 1'd0;
        pe_1_1_clk = 1'd0;
        top_1_1_in = 32'd0;
        top_1_1_write_en = 1'd0;
        top_1_1_clk = 1'd0;
        left_1_1_in = 32'd0;
        left_1_1_write_en = 1'd0;
        left_1_1_clk = 1'd0;
        pe_1_2_top = 32'd0;
        pe_1_2_left = 32'd0;
        pe_1_2_go = 1'd0;
        pe_1_2_clk = 1'd0;
        top_1_2_in = 32'd0;
        top_1_2_write_en = 1'd0;
        top_1_2_clk = 1'd0;
        left_1_2_in = 32'd0;
        left_1_2_write_en = 1'd0;
        left_1_2_clk = 1'd0;
        pe_1_3_top = 32'd0;
        pe_1_3_left = 32'd0;
        pe_1_3_go = 1'd0;
        pe_1_3_clk = 1'd0;
        top_1_3_in = 32'd0;
        top_1_3_write_en = 1'd0;
        top_1_3_clk = 1'd0;
        left_1_3_in = 32'd0;
        left_1_3_write_en = 1'd0;
        left_1_3_clk = 1'd0;
        pe_1_4_top = 32'd0;
        pe_1_4_left = 32'd0;
        pe_1_4_go = 1'd0;
        pe_1_4_clk = 1'd0;
        top_1_4_in = 32'd0;
        top_1_4_write_en = 1'd0;
        top_1_4_clk = 1'd0;
        left_1_4_in = 32'd0;
        left_1_4_write_en = 1'd0;
        left_1_4_clk = 1'd0;
        pe_1_5_top = 32'd0;
        pe_1_5_left = 32'd0;
        pe_1_5_go = 1'd0;
        pe_1_5_clk = 1'd0;
        top_1_5_in = 32'd0;
        top_1_5_write_en = 1'd0;
        top_1_5_clk = 1'd0;
        left_1_5_in = 32'd0;
        left_1_5_write_en = 1'd0;
        left_1_5_clk = 1'd0;
        pe_1_6_top = 32'd0;
        pe_1_6_left = 32'd0;
        pe_1_6_go = 1'd0;
        pe_1_6_clk = 1'd0;
        top_1_6_in = 32'd0;
        top_1_6_write_en = 1'd0;
        top_1_6_clk = 1'd0;
        left_1_6_in = 32'd0;
        left_1_6_write_en = 1'd0;
        left_1_6_clk = 1'd0;
        pe_1_7_top = 32'd0;
        pe_1_7_left = 32'd0;
        pe_1_7_go = 1'd0;
        pe_1_7_clk = 1'd0;
        top_1_7_in = 32'd0;
        top_1_7_write_en = 1'd0;
        top_1_7_clk = 1'd0;
        left_1_7_in = 32'd0;
        left_1_7_write_en = 1'd0;
        left_1_7_clk = 1'd0;
        pe_1_8_top = 32'd0;
        pe_1_8_left = 32'd0;
        pe_1_8_go = 1'd0;
        pe_1_8_clk = 1'd0;
        top_1_8_in = 32'd0;
        top_1_8_write_en = 1'd0;
        top_1_8_clk = 1'd0;
        left_1_8_in = 32'd0;
        left_1_8_write_en = 1'd0;
        left_1_8_clk = 1'd0;
        pe_1_9_top = 32'd0;
        pe_1_9_left = 32'd0;
        pe_1_9_go = 1'd0;
        pe_1_9_clk = 1'd0;
        top_1_9_in = 32'd0;
        top_1_9_write_en = 1'd0;
        top_1_9_clk = 1'd0;
        left_1_9_in = 32'd0;
        left_1_9_write_en = 1'd0;
        left_1_9_clk = 1'd0;
        pe_1_10_top = 32'd0;
        pe_1_10_left = 32'd0;
        pe_1_10_go = 1'd0;
        pe_1_10_clk = 1'd0;
        top_1_10_in = 32'd0;
        top_1_10_write_en = 1'd0;
        top_1_10_clk = 1'd0;
        left_1_10_in = 32'd0;
        left_1_10_write_en = 1'd0;
        left_1_10_clk = 1'd0;
        pe_1_11_top = 32'd0;
        pe_1_11_left = 32'd0;
        pe_1_11_go = 1'd0;
        pe_1_11_clk = 1'd0;
        top_1_11_in = 32'd0;
        top_1_11_write_en = 1'd0;
        top_1_11_clk = 1'd0;
        left_1_11_in = 32'd0;
        left_1_11_write_en = 1'd0;
        left_1_11_clk = 1'd0;
        pe_1_12_top = 32'd0;
        pe_1_12_left = 32'd0;
        pe_1_12_go = 1'd0;
        pe_1_12_clk = 1'd0;
        top_1_12_in = 32'd0;
        top_1_12_write_en = 1'd0;
        top_1_12_clk = 1'd0;
        left_1_12_in = 32'd0;
        left_1_12_write_en = 1'd0;
        left_1_12_clk = 1'd0;
        pe_1_13_top = 32'd0;
        pe_1_13_left = 32'd0;
        pe_1_13_go = 1'd0;
        pe_1_13_clk = 1'd0;
        top_1_13_in = 32'd0;
        top_1_13_write_en = 1'd0;
        top_1_13_clk = 1'd0;
        left_1_13_in = 32'd0;
        left_1_13_write_en = 1'd0;
        left_1_13_clk = 1'd0;
        pe_1_14_top = 32'd0;
        pe_1_14_left = 32'd0;
        pe_1_14_go = 1'd0;
        pe_1_14_clk = 1'd0;
        top_1_14_in = 32'd0;
        top_1_14_write_en = 1'd0;
        top_1_14_clk = 1'd0;
        left_1_14_in = 32'd0;
        left_1_14_write_en = 1'd0;
        left_1_14_clk = 1'd0;
        pe_1_15_top = 32'd0;
        pe_1_15_left = 32'd0;
        pe_1_15_go = 1'd0;
        pe_1_15_clk = 1'd0;
        top_1_15_in = 32'd0;
        top_1_15_write_en = 1'd0;
        top_1_15_clk = 1'd0;
        left_1_15_in = 32'd0;
        left_1_15_write_en = 1'd0;
        left_1_15_clk = 1'd0;
        pe_2_0_top = 32'd0;
        pe_2_0_left = 32'd0;
        pe_2_0_go = 1'd0;
        pe_2_0_clk = 1'd0;
        top_2_0_in = 32'd0;
        top_2_0_write_en = 1'd0;
        top_2_0_clk = 1'd0;
        left_2_0_in = 32'd0;
        left_2_0_write_en = 1'd0;
        left_2_0_clk = 1'd0;
        pe_2_1_top = 32'd0;
        pe_2_1_left = 32'd0;
        pe_2_1_go = 1'd0;
        pe_2_1_clk = 1'd0;
        top_2_1_in = 32'd0;
        top_2_1_write_en = 1'd0;
        top_2_1_clk = 1'd0;
        left_2_1_in = 32'd0;
        left_2_1_write_en = 1'd0;
        left_2_1_clk = 1'd0;
        pe_2_2_top = 32'd0;
        pe_2_2_left = 32'd0;
        pe_2_2_go = 1'd0;
        pe_2_2_clk = 1'd0;
        top_2_2_in = 32'd0;
        top_2_2_write_en = 1'd0;
        top_2_2_clk = 1'd0;
        left_2_2_in = 32'd0;
        left_2_2_write_en = 1'd0;
        left_2_2_clk = 1'd0;
        pe_2_3_top = 32'd0;
        pe_2_3_left = 32'd0;
        pe_2_3_go = 1'd0;
        pe_2_3_clk = 1'd0;
        top_2_3_in = 32'd0;
        top_2_3_write_en = 1'd0;
        top_2_3_clk = 1'd0;
        left_2_3_in = 32'd0;
        left_2_3_write_en = 1'd0;
        left_2_3_clk = 1'd0;
        pe_2_4_top = 32'd0;
        pe_2_4_left = 32'd0;
        pe_2_4_go = 1'd0;
        pe_2_4_clk = 1'd0;
        top_2_4_in = 32'd0;
        top_2_4_write_en = 1'd0;
        top_2_4_clk = 1'd0;
        left_2_4_in = 32'd0;
        left_2_4_write_en = 1'd0;
        left_2_4_clk = 1'd0;
        pe_2_5_top = 32'd0;
        pe_2_5_left = 32'd0;
        pe_2_5_go = 1'd0;
        pe_2_5_clk = 1'd0;
        top_2_5_in = 32'd0;
        top_2_5_write_en = 1'd0;
        top_2_5_clk = 1'd0;
        left_2_5_in = 32'd0;
        left_2_5_write_en = 1'd0;
        left_2_5_clk = 1'd0;
        pe_2_6_top = 32'd0;
        pe_2_6_left = 32'd0;
        pe_2_6_go = 1'd0;
        pe_2_6_clk = 1'd0;
        top_2_6_in = 32'd0;
        top_2_6_write_en = 1'd0;
        top_2_6_clk = 1'd0;
        left_2_6_in = 32'd0;
        left_2_6_write_en = 1'd0;
        left_2_6_clk = 1'd0;
        pe_2_7_top = 32'd0;
        pe_2_7_left = 32'd0;
        pe_2_7_go = 1'd0;
        pe_2_7_clk = 1'd0;
        top_2_7_in = 32'd0;
        top_2_7_write_en = 1'd0;
        top_2_7_clk = 1'd0;
        left_2_7_in = 32'd0;
        left_2_7_write_en = 1'd0;
        left_2_7_clk = 1'd0;
        pe_2_8_top = 32'd0;
        pe_2_8_left = 32'd0;
        pe_2_8_go = 1'd0;
        pe_2_8_clk = 1'd0;
        top_2_8_in = 32'd0;
        top_2_8_write_en = 1'd0;
        top_2_8_clk = 1'd0;
        left_2_8_in = 32'd0;
        left_2_8_write_en = 1'd0;
        left_2_8_clk = 1'd0;
        pe_2_9_top = 32'd0;
        pe_2_9_left = 32'd0;
        pe_2_9_go = 1'd0;
        pe_2_9_clk = 1'd0;
        top_2_9_in = 32'd0;
        top_2_9_write_en = 1'd0;
        top_2_9_clk = 1'd0;
        left_2_9_in = 32'd0;
        left_2_9_write_en = 1'd0;
        left_2_9_clk = 1'd0;
        pe_2_10_top = 32'd0;
        pe_2_10_left = 32'd0;
        pe_2_10_go = 1'd0;
        pe_2_10_clk = 1'd0;
        top_2_10_in = 32'd0;
        top_2_10_write_en = 1'd0;
        top_2_10_clk = 1'd0;
        left_2_10_in = 32'd0;
        left_2_10_write_en = 1'd0;
        left_2_10_clk = 1'd0;
        pe_2_11_top = 32'd0;
        pe_2_11_left = 32'd0;
        pe_2_11_go = 1'd0;
        pe_2_11_clk = 1'd0;
        top_2_11_in = 32'd0;
        top_2_11_write_en = 1'd0;
        top_2_11_clk = 1'd0;
        left_2_11_in = 32'd0;
        left_2_11_write_en = 1'd0;
        left_2_11_clk = 1'd0;
        pe_2_12_top = 32'd0;
        pe_2_12_left = 32'd0;
        pe_2_12_go = 1'd0;
        pe_2_12_clk = 1'd0;
        top_2_12_in = 32'd0;
        top_2_12_write_en = 1'd0;
        top_2_12_clk = 1'd0;
        left_2_12_in = 32'd0;
        left_2_12_write_en = 1'd0;
        left_2_12_clk = 1'd0;
        pe_2_13_top = 32'd0;
        pe_2_13_left = 32'd0;
        pe_2_13_go = 1'd0;
        pe_2_13_clk = 1'd0;
        top_2_13_in = 32'd0;
        top_2_13_write_en = 1'd0;
        top_2_13_clk = 1'd0;
        left_2_13_in = 32'd0;
        left_2_13_write_en = 1'd0;
        left_2_13_clk = 1'd0;
        pe_2_14_top = 32'd0;
        pe_2_14_left = 32'd0;
        pe_2_14_go = 1'd0;
        pe_2_14_clk = 1'd0;
        top_2_14_in = 32'd0;
        top_2_14_write_en = 1'd0;
        top_2_14_clk = 1'd0;
        left_2_14_in = 32'd0;
        left_2_14_write_en = 1'd0;
        left_2_14_clk = 1'd0;
        pe_2_15_top = 32'd0;
        pe_2_15_left = 32'd0;
        pe_2_15_go = 1'd0;
        pe_2_15_clk = 1'd0;
        top_2_15_in = 32'd0;
        top_2_15_write_en = 1'd0;
        top_2_15_clk = 1'd0;
        left_2_15_in = 32'd0;
        left_2_15_write_en = 1'd0;
        left_2_15_clk = 1'd0;
        pe_3_0_top = 32'd0;
        pe_3_0_left = 32'd0;
        pe_3_0_go = 1'd0;
        pe_3_0_clk = 1'd0;
        top_3_0_in = 32'd0;
        top_3_0_write_en = 1'd0;
        top_3_0_clk = 1'd0;
        left_3_0_in = 32'd0;
        left_3_0_write_en = 1'd0;
        left_3_0_clk = 1'd0;
        pe_3_1_top = 32'd0;
        pe_3_1_left = 32'd0;
        pe_3_1_go = 1'd0;
        pe_3_1_clk = 1'd0;
        top_3_1_in = 32'd0;
        top_3_1_write_en = 1'd0;
        top_3_1_clk = 1'd0;
        left_3_1_in = 32'd0;
        left_3_1_write_en = 1'd0;
        left_3_1_clk = 1'd0;
        pe_3_2_top = 32'd0;
        pe_3_2_left = 32'd0;
        pe_3_2_go = 1'd0;
        pe_3_2_clk = 1'd0;
        top_3_2_in = 32'd0;
        top_3_2_write_en = 1'd0;
        top_3_2_clk = 1'd0;
        left_3_2_in = 32'd0;
        left_3_2_write_en = 1'd0;
        left_3_2_clk = 1'd0;
        pe_3_3_top = 32'd0;
        pe_3_3_left = 32'd0;
        pe_3_3_go = 1'd0;
        pe_3_3_clk = 1'd0;
        top_3_3_in = 32'd0;
        top_3_3_write_en = 1'd0;
        top_3_3_clk = 1'd0;
        left_3_3_in = 32'd0;
        left_3_3_write_en = 1'd0;
        left_3_3_clk = 1'd0;
        pe_3_4_top = 32'd0;
        pe_3_4_left = 32'd0;
        pe_3_4_go = 1'd0;
        pe_3_4_clk = 1'd0;
        top_3_4_in = 32'd0;
        top_3_4_write_en = 1'd0;
        top_3_4_clk = 1'd0;
        left_3_4_in = 32'd0;
        left_3_4_write_en = 1'd0;
        left_3_4_clk = 1'd0;
        pe_3_5_top = 32'd0;
        pe_3_5_left = 32'd0;
        pe_3_5_go = 1'd0;
        pe_3_5_clk = 1'd0;
        top_3_5_in = 32'd0;
        top_3_5_write_en = 1'd0;
        top_3_5_clk = 1'd0;
        left_3_5_in = 32'd0;
        left_3_5_write_en = 1'd0;
        left_3_5_clk = 1'd0;
        pe_3_6_top = 32'd0;
        pe_3_6_left = 32'd0;
        pe_3_6_go = 1'd0;
        pe_3_6_clk = 1'd0;
        top_3_6_in = 32'd0;
        top_3_6_write_en = 1'd0;
        top_3_6_clk = 1'd0;
        left_3_6_in = 32'd0;
        left_3_6_write_en = 1'd0;
        left_3_6_clk = 1'd0;
        pe_3_7_top = 32'd0;
        pe_3_7_left = 32'd0;
        pe_3_7_go = 1'd0;
        pe_3_7_clk = 1'd0;
        top_3_7_in = 32'd0;
        top_3_7_write_en = 1'd0;
        top_3_7_clk = 1'd0;
        left_3_7_in = 32'd0;
        left_3_7_write_en = 1'd0;
        left_3_7_clk = 1'd0;
        pe_3_8_top = 32'd0;
        pe_3_8_left = 32'd0;
        pe_3_8_go = 1'd0;
        pe_3_8_clk = 1'd0;
        top_3_8_in = 32'd0;
        top_3_8_write_en = 1'd0;
        top_3_8_clk = 1'd0;
        left_3_8_in = 32'd0;
        left_3_8_write_en = 1'd0;
        left_3_8_clk = 1'd0;
        pe_3_9_top = 32'd0;
        pe_3_9_left = 32'd0;
        pe_3_9_go = 1'd0;
        pe_3_9_clk = 1'd0;
        top_3_9_in = 32'd0;
        top_3_9_write_en = 1'd0;
        top_3_9_clk = 1'd0;
        left_3_9_in = 32'd0;
        left_3_9_write_en = 1'd0;
        left_3_9_clk = 1'd0;
        pe_3_10_top = 32'd0;
        pe_3_10_left = 32'd0;
        pe_3_10_go = 1'd0;
        pe_3_10_clk = 1'd0;
        top_3_10_in = 32'd0;
        top_3_10_write_en = 1'd0;
        top_3_10_clk = 1'd0;
        left_3_10_in = 32'd0;
        left_3_10_write_en = 1'd0;
        left_3_10_clk = 1'd0;
        pe_3_11_top = 32'd0;
        pe_3_11_left = 32'd0;
        pe_3_11_go = 1'd0;
        pe_3_11_clk = 1'd0;
        top_3_11_in = 32'd0;
        top_3_11_write_en = 1'd0;
        top_3_11_clk = 1'd0;
        left_3_11_in = 32'd0;
        left_3_11_write_en = 1'd0;
        left_3_11_clk = 1'd0;
        pe_3_12_top = 32'd0;
        pe_3_12_left = 32'd0;
        pe_3_12_go = 1'd0;
        pe_3_12_clk = 1'd0;
        top_3_12_in = 32'd0;
        top_3_12_write_en = 1'd0;
        top_3_12_clk = 1'd0;
        left_3_12_in = 32'd0;
        left_3_12_write_en = 1'd0;
        left_3_12_clk = 1'd0;
        pe_3_13_top = 32'd0;
        pe_3_13_left = 32'd0;
        pe_3_13_go = 1'd0;
        pe_3_13_clk = 1'd0;
        top_3_13_in = 32'd0;
        top_3_13_write_en = 1'd0;
        top_3_13_clk = 1'd0;
        left_3_13_in = 32'd0;
        left_3_13_write_en = 1'd0;
        left_3_13_clk = 1'd0;
        pe_3_14_top = 32'd0;
        pe_3_14_left = 32'd0;
        pe_3_14_go = 1'd0;
        pe_3_14_clk = 1'd0;
        top_3_14_in = 32'd0;
        top_3_14_write_en = 1'd0;
        top_3_14_clk = 1'd0;
        left_3_14_in = 32'd0;
        left_3_14_write_en = 1'd0;
        left_3_14_clk = 1'd0;
        pe_3_15_top = 32'd0;
        pe_3_15_left = 32'd0;
        pe_3_15_go = 1'd0;
        pe_3_15_clk = 1'd0;
        top_3_15_in = 32'd0;
        top_3_15_write_en = 1'd0;
        top_3_15_clk = 1'd0;
        left_3_15_in = 32'd0;
        left_3_15_write_en = 1'd0;
        left_3_15_clk = 1'd0;
        pe_4_0_top = 32'd0;
        pe_4_0_left = 32'd0;
        pe_4_0_go = 1'd0;
        pe_4_0_clk = 1'd0;
        top_4_0_in = 32'd0;
        top_4_0_write_en = 1'd0;
        top_4_0_clk = 1'd0;
        left_4_0_in = 32'd0;
        left_4_0_write_en = 1'd0;
        left_4_0_clk = 1'd0;
        pe_4_1_top = 32'd0;
        pe_4_1_left = 32'd0;
        pe_4_1_go = 1'd0;
        pe_4_1_clk = 1'd0;
        top_4_1_in = 32'd0;
        top_4_1_write_en = 1'd0;
        top_4_1_clk = 1'd0;
        left_4_1_in = 32'd0;
        left_4_1_write_en = 1'd0;
        left_4_1_clk = 1'd0;
        pe_4_2_top = 32'd0;
        pe_4_2_left = 32'd0;
        pe_4_2_go = 1'd0;
        pe_4_2_clk = 1'd0;
        top_4_2_in = 32'd0;
        top_4_2_write_en = 1'd0;
        top_4_2_clk = 1'd0;
        left_4_2_in = 32'd0;
        left_4_2_write_en = 1'd0;
        left_4_2_clk = 1'd0;
        pe_4_3_top = 32'd0;
        pe_4_3_left = 32'd0;
        pe_4_3_go = 1'd0;
        pe_4_3_clk = 1'd0;
        top_4_3_in = 32'd0;
        top_4_3_write_en = 1'd0;
        top_4_3_clk = 1'd0;
        left_4_3_in = 32'd0;
        left_4_3_write_en = 1'd0;
        left_4_3_clk = 1'd0;
        pe_4_4_top = 32'd0;
        pe_4_4_left = 32'd0;
        pe_4_4_go = 1'd0;
        pe_4_4_clk = 1'd0;
        top_4_4_in = 32'd0;
        top_4_4_write_en = 1'd0;
        top_4_4_clk = 1'd0;
        left_4_4_in = 32'd0;
        left_4_4_write_en = 1'd0;
        left_4_4_clk = 1'd0;
        pe_4_5_top = 32'd0;
        pe_4_5_left = 32'd0;
        pe_4_5_go = 1'd0;
        pe_4_5_clk = 1'd0;
        top_4_5_in = 32'd0;
        top_4_5_write_en = 1'd0;
        top_4_5_clk = 1'd0;
        left_4_5_in = 32'd0;
        left_4_5_write_en = 1'd0;
        left_4_5_clk = 1'd0;
        pe_4_6_top = 32'd0;
        pe_4_6_left = 32'd0;
        pe_4_6_go = 1'd0;
        pe_4_6_clk = 1'd0;
        top_4_6_in = 32'd0;
        top_4_6_write_en = 1'd0;
        top_4_6_clk = 1'd0;
        left_4_6_in = 32'd0;
        left_4_6_write_en = 1'd0;
        left_4_6_clk = 1'd0;
        pe_4_7_top = 32'd0;
        pe_4_7_left = 32'd0;
        pe_4_7_go = 1'd0;
        pe_4_7_clk = 1'd0;
        top_4_7_in = 32'd0;
        top_4_7_write_en = 1'd0;
        top_4_7_clk = 1'd0;
        left_4_7_in = 32'd0;
        left_4_7_write_en = 1'd0;
        left_4_7_clk = 1'd0;
        pe_4_8_top = 32'd0;
        pe_4_8_left = 32'd0;
        pe_4_8_go = 1'd0;
        pe_4_8_clk = 1'd0;
        top_4_8_in = 32'd0;
        top_4_8_write_en = 1'd0;
        top_4_8_clk = 1'd0;
        left_4_8_in = 32'd0;
        left_4_8_write_en = 1'd0;
        left_4_8_clk = 1'd0;
        pe_4_9_top = 32'd0;
        pe_4_9_left = 32'd0;
        pe_4_9_go = 1'd0;
        pe_4_9_clk = 1'd0;
        top_4_9_in = 32'd0;
        top_4_9_write_en = 1'd0;
        top_4_9_clk = 1'd0;
        left_4_9_in = 32'd0;
        left_4_9_write_en = 1'd0;
        left_4_9_clk = 1'd0;
        pe_4_10_top = 32'd0;
        pe_4_10_left = 32'd0;
        pe_4_10_go = 1'd0;
        pe_4_10_clk = 1'd0;
        top_4_10_in = 32'd0;
        top_4_10_write_en = 1'd0;
        top_4_10_clk = 1'd0;
        left_4_10_in = 32'd0;
        left_4_10_write_en = 1'd0;
        left_4_10_clk = 1'd0;
        pe_4_11_top = 32'd0;
        pe_4_11_left = 32'd0;
        pe_4_11_go = 1'd0;
        pe_4_11_clk = 1'd0;
        top_4_11_in = 32'd0;
        top_4_11_write_en = 1'd0;
        top_4_11_clk = 1'd0;
        left_4_11_in = 32'd0;
        left_4_11_write_en = 1'd0;
        left_4_11_clk = 1'd0;
        pe_4_12_top = 32'd0;
        pe_4_12_left = 32'd0;
        pe_4_12_go = 1'd0;
        pe_4_12_clk = 1'd0;
        top_4_12_in = 32'd0;
        top_4_12_write_en = 1'd0;
        top_4_12_clk = 1'd0;
        left_4_12_in = 32'd0;
        left_4_12_write_en = 1'd0;
        left_4_12_clk = 1'd0;
        pe_4_13_top = 32'd0;
        pe_4_13_left = 32'd0;
        pe_4_13_go = 1'd0;
        pe_4_13_clk = 1'd0;
        top_4_13_in = 32'd0;
        top_4_13_write_en = 1'd0;
        top_4_13_clk = 1'd0;
        left_4_13_in = 32'd0;
        left_4_13_write_en = 1'd0;
        left_4_13_clk = 1'd0;
        pe_4_14_top = 32'd0;
        pe_4_14_left = 32'd0;
        pe_4_14_go = 1'd0;
        pe_4_14_clk = 1'd0;
        top_4_14_in = 32'd0;
        top_4_14_write_en = 1'd0;
        top_4_14_clk = 1'd0;
        left_4_14_in = 32'd0;
        left_4_14_write_en = 1'd0;
        left_4_14_clk = 1'd0;
        pe_4_15_top = 32'd0;
        pe_4_15_left = 32'd0;
        pe_4_15_go = 1'd0;
        pe_4_15_clk = 1'd0;
        top_4_15_in = 32'd0;
        top_4_15_write_en = 1'd0;
        top_4_15_clk = 1'd0;
        left_4_15_in = 32'd0;
        left_4_15_write_en = 1'd0;
        left_4_15_clk = 1'd0;
        pe_5_0_top = 32'd0;
        pe_5_0_left = 32'd0;
        pe_5_0_go = 1'd0;
        pe_5_0_clk = 1'd0;
        top_5_0_in = 32'd0;
        top_5_0_write_en = 1'd0;
        top_5_0_clk = 1'd0;
        left_5_0_in = 32'd0;
        left_5_0_write_en = 1'd0;
        left_5_0_clk = 1'd0;
        pe_5_1_top = 32'd0;
        pe_5_1_left = 32'd0;
        pe_5_1_go = 1'd0;
        pe_5_1_clk = 1'd0;
        top_5_1_in = 32'd0;
        top_5_1_write_en = 1'd0;
        top_5_1_clk = 1'd0;
        left_5_1_in = 32'd0;
        left_5_1_write_en = 1'd0;
        left_5_1_clk = 1'd0;
        pe_5_2_top = 32'd0;
        pe_5_2_left = 32'd0;
        pe_5_2_go = 1'd0;
        pe_5_2_clk = 1'd0;
        top_5_2_in = 32'd0;
        top_5_2_write_en = 1'd0;
        top_5_2_clk = 1'd0;
        left_5_2_in = 32'd0;
        left_5_2_write_en = 1'd0;
        left_5_2_clk = 1'd0;
        pe_5_3_top = 32'd0;
        pe_5_3_left = 32'd0;
        pe_5_3_go = 1'd0;
        pe_5_3_clk = 1'd0;
        top_5_3_in = 32'd0;
        top_5_3_write_en = 1'd0;
        top_5_3_clk = 1'd0;
        left_5_3_in = 32'd0;
        left_5_3_write_en = 1'd0;
        left_5_3_clk = 1'd0;
        pe_5_4_top = 32'd0;
        pe_5_4_left = 32'd0;
        pe_5_4_go = 1'd0;
        pe_5_4_clk = 1'd0;
        top_5_4_in = 32'd0;
        top_5_4_write_en = 1'd0;
        top_5_4_clk = 1'd0;
        left_5_4_in = 32'd0;
        left_5_4_write_en = 1'd0;
        left_5_4_clk = 1'd0;
        pe_5_5_top = 32'd0;
        pe_5_5_left = 32'd0;
        pe_5_5_go = 1'd0;
        pe_5_5_clk = 1'd0;
        top_5_5_in = 32'd0;
        top_5_5_write_en = 1'd0;
        top_5_5_clk = 1'd0;
        left_5_5_in = 32'd0;
        left_5_5_write_en = 1'd0;
        left_5_5_clk = 1'd0;
        pe_5_6_top = 32'd0;
        pe_5_6_left = 32'd0;
        pe_5_6_go = 1'd0;
        pe_5_6_clk = 1'd0;
        top_5_6_in = 32'd0;
        top_5_6_write_en = 1'd0;
        top_5_6_clk = 1'd0;
        left_5_6_in = 32'd0;
        left_5_6_write_en = 1'd0;
        left_5_6_clk = 1'd0;
        pe_5_7_top = 32'd0;
        pe_5_7_left = 32'd0;
        pe_5_7_go = 1'd0;
        pe_5_7_clk = 1'd0;
        top_5_7_in = 32'd0;
        top_5_7_write_en = 1'd0;
        top_5_7_clk = 1'd0;
        left_5_7_in = 32'd0;
        left_5_7_write_en = 1'd0;
        left_5_7_clk = 1'd0;
        pe_5_8_top = 32'd0;
        pe_5_8_left = 32'd0;
        pe_5_8_go = 1'd0;
        pe_5_8_clk = 1'd0;
        top_5_8_in = 32'd0;
        top_5_8_write_en = 1'd0;
        top_5_8_clk = 1'd0;
        left_5_8_in = 32'd0;
        left_5_8_write_en = 1'd0;
        left_5_8_clk = 1'd0;
        pe_5_9_top = 32'd0;
        pe_5_9_left = 32'd0;
        pe_5_9_go = 1'd0;
        pe_5_9_clk = 1'd0;
        top_5_9_in = 32'd0;
        top_5_9_write_en = 1'd0;
        top_5_9_clk = 1'd0;
        left_5_9_in = 32'd0;
        left_5_9_write_en = 1'd0;
        left_5_9_clk = 1'd0;
        pe_5_10_top = 32'd0;
        pe_5_10_left = 32'd0;
        pe_5_10_go = 1'd0;
        pe_5_10_clk = 1'd0;
        top_5_10_in = 32'd0;
        top_5_10_write_en = 1'd0;
        top_5_10_clk = 1'd0;
        left_5_10_in = 32'd0;
        left_5_10_write_en = 1'd0;
        left_5_10_clk = 1'd0;
        pe_5_11_top = 32'd0;
        pe_5_11_left = 32'd0;
        pe_5_11_go = 1'd0;
        pe_5_11_clk = 1'd0;
        top_5_11_in = 32'd0;
        top_5_11_write_en = 1'd0;
        top_5_11_clk = 1'd0;
        left_5_11_in = 32'd0;
        left_5_11_write_en = 1'd0;
        left_5_11_clk = 1'd0;
        pe_5_12_top = 32'd0;
        pe_5_12_left = 32'd0;
        pe_5_12_go = 1'd0;
        pe_5_12_clk = 1'd0;
        top_5_12_in = 32'd0;
        top_5_12_write_en = 1'd0;
        top_5_12_clk = 1'd0;
        left_5_12_in = 32'd0;
        left_5_12_write_en = 1'd0;
        left_5_12_clk = 1'd0;
        pe_5_13_top = 32'd0;
        pe_5_13_left = 32'd0;
        pe_5_13_go = 1'd0;
        pe_5_13_clk = 1'd0;
        top_5_13_in = 32'd0;
        top_5_13_write_en = 1'd0;
        top_5_13_clk = 1'd0;
        left_5_13_in = 32'd0;
        left_5_13_write_en = 1'd0;
        left_5_13_clk = 1'd0;
        pe_5_14_top = 32'd0;
        pe_5_14_left = 32'd0;
        pe_5_14_go = 1'd0;
        pe_5_14_clk = 1'd0;
        top_5_14_in = 32'd0;
        top_5_14_write_en = 1'd0;
        top_5_14_clk = 1'd0;
        left_5_14_in = 32'd0;
        left_5_14_write_en = 1'd0;
        left_5_14_clk = 1'd0;
        pe_5_15_top = 32'd0;
        pe_5_15_left = 32'd0;
        pe_5_15_go = 1'd0;
        pe_5_15_clk = 1'd0;
        top_5_15_in = 32'd0;
        top_5_15_write_en = 1'd0;
        top_5_15_clk = 1'd0;
        left_5_15_in = 32'd0;
        left_5_15_write_en = 1'd0;
        left_5_15_clk = 1'd0;
        pe_6_0_top = 32'd0;
        pe_6_0_left = 32'd0;
        pe_6_0_go = 1'd0;
        pe_6_0_clk = 1'd0;
        top_6_0_in = 32'd0;
        top_6_0_write_en = 1'd0;
        top_6_0_clk = 1'd0;
        left_6_0_in = 32'd0;
        left_6_0_write_en = 1'd0;
        left_6_0_clk = 1'd0;
        pe_6_1_top = 32'd0;
        pe_6_1_left = 32'd0;
        pe_6_1_go = 1'd0;
        pe_6_1_clk = 1'd0;
        top_6_1_in = 32'd0;
        top_6_1_write_en = 1'd0;
        top_6_1_clk = 1'd0;
        left_6_1_in = 32'd0;
        left_6_1_write_en = 1'd0;
        left_6_1_clk = 1'd0;
        pe_6_2_top = 32'd0;
        pe_6_2_left = 32'd0;
        pe_6_2_go = 1'd0;
        pe_6_2_clk = 1'd0;
        top_6_2_in = 32'd0;
        top_6_2_write_en = 1'd0;
        top_6_2_clk = 1'd0;
        left_6_2_in = 32'd0;
        left_6_2_write_en = 1'd0;
        left_6_2_clk = 1'd0;
        pe_6_3_top = 32'd0;
        pe_6_3_left = 32'd0;
        pe_6_3_go = 1'd0;
        pe_6_3_clk = 1'd0;
        top_6_3_in = 32'd0;
        top_6_3_write_en = 1'd0;
        top_6_3_clk = 1'd0;
        left_6_3_in = 32'd0;
        left_6_3_write_en = 1'd0;
        left_6_3_clk = 1'd0;
        pe_6_4_top = 32'd0;
        pe_6_4_left = 32'd0;
        pe_6_4_go = 1'd0;
        pe_6_4_clk = 1'd0;
        top_6_4_in = 32'd0;
        top_6_4_write_en = 1'd0;
        top_6_4_clk = 1'd0;
        left_6_4_in = 32'd0;
        left_6_4_write_en = 1'd0;
        left_6_4_clk = 1'd0;
        pe_6_5_top = 32'd0;
        pe_6_5_left = 32'd0;
        pe_6_5_go = 1'd0;
        pe_6_5_clk = 1'd0;
        top_6_5_in = 32'd0;
        top_6_5_write_en = 1'd0;
        top_6_5_clk = 1'd0;
        left_6_5_in = 32'd0;
        left_6_5_write_en = 1'd0;
        left_6_5_clk = 1'd0;
        pe_6_6_top = 32'd0;
        pe_6_6_left = 32'd0;
        pe_6_6_go = 1'd0;
        pe_6_6_clk = 1'd0;
        top_6_6_in = 32'd0;
        top_6_6_write_en = 1'd0;
        top_6_6_clk = 1'd0;
        left_6_6_in = 32'd0;
        left_6_6_write_en = 1'd0;
        left_6_6_clk = 1'd0;
        pe_6_7_top = 32'd0;
        pe_6_7_left = 32'd0;
        pe_6_7_go = 1'd0;
        pe_6_7_clk = 1'd0;
        top_6_7_in = 32'd0;
        top_6_7_write_en = 1'd0;
        top_6_7_clk = 1'd0;
        left_6_7_in = 32'd0;
        left_6_7_write_en = 1'd0;
        left_6_7_clk = 1'd0;
        pe_6_8_top = 32'd0;
        pe_6_8_left = 32'd0;
        pe_6_8_go = 1'd0;
        pe_6_8_clk = 1'd0;
        top_6_8_in = 32'd0;
        top_6_8_write_en = 1'd0;
        top_6_8_clk = 1'd0;
        left_6_8_in = 32'd0;
        left_6_8_write_en = 1'd0;
        left_6_8_clk = 1'd0;
        pe_6_9_top = 32'd0;
        pe_6_9_left = 32'd0;
        pe_6_9_go = 1'd0;
        pe_6_9_clk = 1'd0;
        top_6_9_in = 32'd0;
        top_6_9_write_en = 1'd0;
        top_6_9_clk = 1'd0;
        left_6_9_in = 32'd0;
        left_6_9_write_en = 1'd0;
        left_6_9_clk = 1'd0;
        pe_6_10_top = 32'd0;
        pe_6_10_left = 32'd0;
        pe_6_10_go = 1'd0;
        pe_6_10_clk = 1'd0;
        top_6_10_in = 32'd0;
        top_6_10_write_en = 1'd0;
        top_6_10_clk = 1'd0;
        left_6_10_in = 32'd0;
        left_6_10_write_en = 1'd0;
        left_6_10_clk = 1'd0;
        pe_6_11_top = 32'd0;
        pe_6_11_left = 32'd0;
        pe_6_11_go = 1'd0;
        pe_6_11_clk = 1'd0;
        top_6_11_in = 32'd0;
        top_6_11_write_en = 1'd0;
        top_6_11_clk = 1'd0;
        left_6_11_in = 32'd0;
        left_6_11_write_en = 1'd0;
        left_6_11_clk = 1'd0;
        pe_6_12_top = 32'd0;
        pe_6_12_left = 32'd0;
        pe_6_12_go = 1'd0;
        pe_6_12_clk = 1'd0;
        top_6_12_in = 32'd0;
        top_6_12_write_en = 1'd0;
        top_6_12_clk = 1'd0;
        left_6_12_in = 32'd0;
        left_6_12_write_en = 1'd0;
        left_6_12_clk = 1'd0;
        pe_6_13_top = 32'd0;
        pe_6_13_left = 32'd0;
        pe_6_13_go = 1'd0;
        pe_6_13_clk = 1'd0;
        top_6_13_in = 32'd0;
        top_6_13_write_en = 1'd0;
        top_6_13_clk = 1'd0;
        left_6_13_in = 32'd0;
        left_6_13_write_en = 1'd0;
        left_6_13_clk = 1'd0;
        pe_6_14_top = 32'd0;
        pe_6_14_left = 32'd0;
        pe_6_14_go = 1'd0;
        pe_6_14_clk = 1'd0;
        top_6_14_in = 32'd0;
        top_6_14_write_en = 1'd0;
        top_6_14_clk = 1'd0;
        left_6_14_in = 32'd0;
        left_6_14_write_en = 1'd0;
        left_6_14_clk = 1'd0;
        pe_6_15_top = 32'd0;
        pe_6_15_left = 32'd0;
        pe_6_15_go = 1'd0;
        pe_6_15_clk = 1'd0;
        top_6_15_in = 32'd0;
        top_6_15_write_en = 1'd0;
        top_6_15_clk = 1'd0;
        left_6_15_in = 32'd0;
        left_6_15_write_en = 1'd0;
        left_6_15_clk = 1'd0;
        pe_7_0_top = 32'd0;
        pe_7_0_left = 32'd0;
        pe_7_0_go = 1'd0;
        pe_7_0_clk = 1'd0;
        top_7_0_in = 32'd0;
        top_7_0_write_en = 1'd0;
        top_7_0_clk = 1'd0;
        left_7_0_in = 32'd0;
        left_7_0_write_en = 1'd0;
        left_7_0_clk = 1'd0;
        pe_7_1_top = 32'd0;
        pe_7_1_left = 32'd0;
        pe_7_1_go = 1'd0;
        pe_7_1_clk = 1'd0;
        top_7_1_in = 32'd0;
        top_7_1_write_en = 1'd0;
        top_7_1_clk = 1'd0;
        left_7_1_in = 32'd0;
        left_7_1_write_en = 1'd0;
        left_7_1_clk = 1'd0;
        pe_7_2_top = 32'd0;
        pe_7_2_left = 32'd0;
        pe_7_2_go = 1'd0;
        pe_7_2_clk = 1'd0;
        top_7_2_in = 32'd0;
        top_7_2_write_en = 1'd0;
        top_7_2_clk = 1'd0;
        left_7_2_in = 32'd0;
        left_7_2_write_en = 1'd0;
        left_7_2_clk = 1'd0;
        pe_7_3_top = 32'd0;
        pe_7_3_left = 32'd0;
        pe_7_3_go = 1'd0;
        pe_7_3_clk = 1'd0;
        top_7_3_in = 32'd0;
        top_7_3_write_en = 1'd0;
        top_7_3_clk = 1'd0;
        left_7_3_in = 32'd0;
        left_7_3_write_en = 1'd0;
        left_7_3_clk = 1'd0;
        pe_7_4_top = 32'd0;
        pe_7_4_left = 32'd0;
        pe_7_4_go = 1'd0;
        pe_7_4_clk = 1'd0;
        top_7_4_in = 32'd0;
        top_7_4_write_en = 1'd0;
        top_7_4_clk = 1'd0;
        left_7_4_in = 32'd0;
        left_7_4_write_en = 1'd0;
        left_7_4_clk = 1'd0;
        pe_7_5_top = 32'd0;
        pe_7_5_left = 32'd0;
        pe_7_5_go = 1'd0;
        pe_7_5_clk = 1'd0;
        top_7_5_in = 32'd0;
        top_7_5_write_en = 1'd0;
        top_7_5_clk = 1'd0;
        left_7_5_in = 32'd0;
        left_7_5_write_en = 1'd0;
        left_7_5_clk = 1'd0;
        pe_7_6_top = 32'd0;
        pe_7_6_left = 32'd0;
        pe_7_6_go = 1'd0;
        pe_7_6_clk = 1'd0;
        top_7_6_in = 32'd0;
        top_7_6_write_en = 1'd0;
        top_7_6_clk = 1'd0;
        left_7_6_in = 32'd0;
        left_7_6_write_en = 1'd0;
        left_7_6_clk = 1'd0;
        pe_7_7_top = 32'd0;
        pe_7_7_left = 32'd0;
        pe_7_7_go = 1'd0;
        pe_7_7_clk = 1'd0;
        top_7_7_in = 32'd0;
        top_7_7_write_en = 1'd0;
        top_7_7_clk = 1'd0;
        left_7_7_in = 32'd0;
        left_7_7_write_en = 1'd0;
        left_7_7_clk = 1'd0;
        pe_7_8_top = 32'd0;
        pe_7_8_left = 32'd0;
        pe_7_8_go = 1'd0;
        pe_7_8_clk = 1'd0;
        top_7_8_in = 32'd0;
        top_7_8_write_en = 1'd0;
        top_7_8_clk = 1'd0;
        left_7_8_in = 32'd0;
        left_7_8_write_en = 1'd0;
        left_7_8_clk = 1'd0;
        pe_7_9_top = 32'd0;
        pe_7_9_left = 32'd0;
        pe_7_9_go = 1'd0;
        pe_7_9_clk = 1'd0;
        top_7_9_in = 32'd0;
        top_7_9_write_en = 1'd0;
        top_7_9_clk = 1'd0;
        left_7_9_in = 32'd0;
        left_7_9_write_en = 1'd0;
        left_7_9_clk = 1'd0;
        pe_7_10_top = 32'd0;
        pe_7_10_left = 32'd0;
        pe_7_10_go = 1'd0;
        pe_7_10_clk = 1'd0;
        top_7_10_in = 32'd0;
        top_7_10_write_en = 1'd0;
        top_7_10_clk = 1'd0;
        left_7_10_in = 32'd0;
        left_7_10_write_en = 1'd0;
        left_7_10_clk = 1'd0;
        pe_7_11_top = 32'd0;
        pe_7_11_left = 32'd0;
        pe_7_11_go = 1'd0;
        pe_7_11_clk = 1'd0;
        top_7_11_in = 32'd0;
        top_7_11_write_en = 1'd0;
        top_7_11_clk = 1'd0;
        left_7_11_in = 32'd0;
        left_7_11_write_en = 1'd0;
        left_7_11_clk = 1'd0;
        pe_7_12_top = 32'd0;
        pe_7_12_left = 32'd0;
        pe_7_12_go = 1'd0;
        pe_7_12_clk = 1'd0;
        top_7_12_in = 32'd0;
        top_7_12_write_en = 1'd0;
        top_7_12_clk = 1'd0;
        left_7_12_in = 32'd0;
        left_7_12_write_en = 1'd0;
        left_7_12_clk = 1'd0;
        pe_7_13_top = 32'd0;
        pe_7_13_left = 32'd0;
        pe_7_13_go = 1'd0;
        pe_7_13_clk = 1'd0;
        top_7_13_in = 32'd0;
        top_7_13_write_en = 1'd0;
        top_7_13_clk = 1'd0;
        left_7_13_in = 32'd0;
        left_7_13_write_en = 1'd0;
        left_7_13_clk = 1'd0;
        pe_7_14_top = 32'd0;
        pe_7_14_left = 32'd0;
        pe_7_14_go = 1'd0;
        pe_7_14_clk = 1'd0;
        top_7_14_in = 32'd0;
        top_7_14_write_en = 1'd0;
        top_7_14_clk = 1'd0;
        left_7_14_in = 32'd0;
        left_7_14_write_en = 1'd0;
        left_7_14_clk = 1'd0;
        pe_7_15_top = 32'd0;
        pe_7_15_left = 32'd0;
        pe_7_15_go = 1'd0;
        pe_7_15_clk = 1'd0;
        top_7_15_in = 32'd0;
        top_7_15_write_en = 1'd0;
        top_7_15_clk = 1'd0;
        left_7_15_in = 32'd0;
        left_7_15_write_en = 1'd0;
        left_7_15_clk = 1'd0;
        pe_8_0_top = 32'd0;
        pe_8_0_left = 32'd0;
        pe_8_0_go = 1'd0;
        pe_8_0_clk = 1'd0;
        top_8_0_in = 32'd0;
        top_8_0_write_en = 1'd0;
        top_8_0_clk = 1'd0;
        left_8_0_in = 32'd0;
        left_8_0_write_en = 1'd0;
        left_8_0_clk = 1'd0;
        pe_8_1_top = 32'd0;
        pe_8_1_left = 32'd0;
        pe_8_1_go = 1'd0;
        pe_8_1_clk = 1'd0;
        top_8_1_in = 32'd0;
        top_8_1_write_en = 1'd0;
        top_8_1_clk = 1'd0;
        left_8_1_in = 32'd0;
        left_8_1_write_en = 1'd0;
        left_8_1_clk = 1'd0;
        pe_8_2_top = 32'd0;
        pe_8_2_left = 32'd0;
        pe_8_2_go = 1'd0;
        pe_8_2_clk = 1'd0;
        top_8_2_in = 32'd0;
        top_8_2_write_en = 1'd0;
        top_8_2_clk = 1'd0;
        left_8_2_in = 32'd0;
        left_8_2_write_en = 1'd0;
        left_8_2_clk = 1'd0;
        pe_8_3_top = 32'd0;
        pe_8_3_left = 32'd0;
        pe_8_3_go = 1'd0;
        pe_8_3_clk = 1'd0;
        top_8_3_in = 32'd0;
        top_8_3_write_en = 1'd0;
        top_8_3_clk = 1'd0;
        left_8_3_in = 32'd0;
        left_8_3_write_en = 1'd0;
        left_8_3_clk = 1'd0;
        pe_8_4_top = 32'd0;
        pe_8_4_left = 32'd0;
        pe_8_4_go = 1'd0;
        pe_8_4_clk = 1'd0;
        top_8_4_in = 32'd0;
        top_8_4_write_en = 1'd0;
        top_8_4_clk = 1'd0;
        left_8_4_in = 32'd0;
        left_8_4_write_en = 1'd0;
        left_8_4_clk = 1'd0;
        pe_8_5_top = 32'd0;
        pe_8_5_left = 32'd0;
        pe_8_5_go = 1'd0;
        pe_8_5_clk = 1'd0;
        top_8_5_in = 32'd0;
        top_8_5_write_en = 1'd0;
        top_8_5_clk = 1'd0;
        left_8_5_in = 32'd0;
        left_8_5_write_en = 1'd0;
        left_8_5_clk = 1'd0;
        pe_8_6_top = 32'd0;
        pe_8_6_left = 32'd0;
        pe_8_6_go = 1'd0;
        pe_8_6_clk = 1'd0;
        top_8_6_in = 32'd0;
        top_8_6_write_en = 1'd0;
        top_8_6_clk = 1'd0;
        left_8_6_in = 32'd0;
        left_8_6_write_en = 1'd0;
        left_8_6_clk = 1'd0;
        pe_8_7_top = 32'd0;
        pe_8_7_left = 32'd0;
        pe_8_7_go = 1'd0;
        pe_8_7_clk = 1'd0;
        top_8_7_in = 32'd0;
        top_8_7_write_en = 1'd0;
        top_8_7_clk = 1'd0;
        left_8_7_in = 32'd0;
        left_8_7_write_en = 1'd0;
        left_8_7_clk = 1'd0;
        pe_8_8_top = 32'd0;
        pe_8_8_left = 32'd0;
        pe_8_8_go = 1'd0;
        pe_8_8_clk = 1'd0;
        top_8_8_in = 32'd0;
        top_8_8_write_en = 1'd0;
        top_8_8_clk = 1'd0;
        left_8_8_in = 32'd0;
        left_8_8_write_en = 1'd0;
        left_8_8_clk = 1'd0;
        pe_8_9_top = 32'd0;
        pe_8_9_left = 32'd0;
        pe_8_9_go = 1'd0;
        pe_8_9_clk = 1'd0;
        top_8_9_in = 32'd0;
        top_8_9_write_en = 1'd0;
        top_8_9_clk = 1'd0;
        left_8_9_in = 32'd0;
        left_8_9_write_en = 1'd0;
        left_8_9_clk = 1'd0;
        pe_8_10_top = 32'd0;
        pe_8_10_left = 32'd0;
        pe_8_10_go = 1'd0;
        pe_8_10_clk = 1'd0;
        top_8_10_in = 32'd0;
        top_8_10_write_en = 1'd0;
        top_8_10_clk = 1'd0;
        left_8_10_in = 32'd0;
        left_8_10_write_en = 1'd0;
        left_8_10_clk = 1'd0;
        pe_8_11_top = 32'd0;
        pe_8_11_left = 32'd0;
        pe_8_11_go = 1'd0;
        pe_8_11_clk = 1'd0;
        top_8_11_in = 32'd0;
        top_8_11_write_en = 1'd0;
        top_8_11_clk = 1'd0;
        left_8_11_in = 32'd0;
        left_8_11_write_en = 1'd0;
        left_8_11_clk = 1'd0;
        pe_8_12_top = 32'd0;
        pe_8_12_left = 32'd0;
        pe_8_12_go = 1'd0;
        pe_8_12_clk = 1'd0;
        top_8_12_in = 32'd0;
        top_8_12_write_en = 1'd0;
        top_8_12_clk = 1'd0;
        left_8_12_in = 32'd0;
        left_8_12_write_en = 1'd0;
        left_8_12_clk = 1'd0;
        pe_8_13_top = 32'd0;
        pe_8_13_left = 32'd0;
        pe_8_13_go = 1'd0;
        pe_8_13_clk = 1'd0;
        top_8_13_in = 32'd0;
        top_8_13_write_en = 1'd0;
        top_8_13_clk = 1'd0;
        left_8_13_in = 32'd0;
        left_8_13_write_en = 1'd0;
        left_8_13_clk = 1'd0;
        pe_8_14_top = 32'd0;
        pe_8_14_left = 32'd0;
        pe_8_14_go = 1'd0;
        pe_8_14_clk = 1'd0;
        top_8_14_in = 32'd0;
        top_8_14_write_en = 1'd0;
        top_8_14_clk = 1'd0;
        left_8_14_in = 32'd0;
        left_8_14_write_en = 1'd0;
        left_8_14_clk = 1'd0;
        pe_8_15_top = 32'd0;
        pe_8_15_left = 32'd0;
        pe_8_15_go = 1'd0;
        pe_8_15_clk = 1'd0;
        top_8_15_in = 32'd0;
        top_8_15_write_en = 1'd0;
        top_8_15_clk = 1'd0;
        left_8_15_in = 32'd0;
        left_8_15_write_en = 1'd0;
        left_8_15_clk = 1'd0;
        pe_9_0_top = 32'd0;
        pe_9_0_left = 32'd0;
        pe_9_0_go = 1'd0;
        pe_9_0_clk = 1'd0;
        top_9_0_in = 32'd0;
        top_9_0_write_en = 1'd0;
        top_9_0_clk = 1'd0;
        left_9_0_in = 32'd0;
        left_9_0_write_en = 1'd0;
        left_9_0_clk = 1'd0;
        pe_9_1_top = 32'd0;
        pe_9_1_left = 32'd0;
        pe_9_1_go = 1'd0;
        pe_9_1_clk = 1'd0;
        top_9_1_in = 32'd0;
        top_9_1_write_en = 1'd0;
        top_9_1_clk = 1'd0;
        left_9_1_in = 32'd0;
        left_9_1_write_en = 1'd0;
        left_9_1_clk = 1'd0;
        pe_9_2_top = 32'd0;
        pe_9_2_left = 32'd0;
        pe_9_2_go = 1'd0;
        pe_9_2_clk = 1'd0;
        top_9_2_in = 32'd0;
        top_9_2_write_en = 1'd0;
        top_9_2_clk = 1'd0;
        left_9_2_in = 32'd0;
        left_9_2_write_en = 1'd0;
        left_9_2_clk = 1'd0;
        pe_9_3_top = 32'd0;
        pe_9_3_left = 32'd0;
        pe_9_3_go = 1'd0;
        pe_9_3_clk = 1'd0;
        top_9_3_in = 32'd0;
        top_9_3_write_en = 1'd0;
        top_9_3_clk = 1'd0;
        left_9_3_in = 32'd0;
        left_9_3_write_en = 1'd0;
        left_9_3_clk = 1'd0;
        pe_9_4_top = 32'd0;
        pe_9_4_left = 32'd0;
        pe_9_4_go = 1'd0;
        pe_9_4_clk = 1'd0;
        top_9_4_in = 32'd0;
        top_9_4_write_en = 1'd0;
        top_9_4_clk = 1'd0;
        left_9_4_in = 32'd0;
        left_9_4_write_en = 1'd0;
        left_9_4_clk = 1'd0;
        pe_9_5_top = 32'd0;
        pe_9_5_left = 32'd0;
        pe_9_5_go = 1'd0;
        pe_9_5_clk = 1'd0;
        top_9_5_in = 32'd0;
        top_9_5_write_en = 1'd0;
        top_9_5_clk = 1'd0;
        left_9_5_in = 32'd0;
        left_9_5_write_en = 1'd0;
        left_9_5_clk = 1'd0;
        pe_9_6_top = 32'd0;
        pe_9_6_left = 32'd0;
        pe_9_6_go = 1'd0;
        pe_9_6_clk = 1'd0;
        top_9_6_in = 32'd0;
        top_9_6_write_en = 1'd0;
        top_9_6_clk = 1'd0;
        left_9_6_in = 32'd0;
        left_9_6_write_en = 1'd0;
        left_9_6_clk = 1'd0;
        pe_9_7_top = 32'd0;
        pe_9_7_left = 32'd0;
        pe_9_7_go = 1'd0;
        pe_9_7_clk = 1'd0;
        top_9_7_in = 32'd0;
        top_9_7_write_en = 1'd0;
        top_9_7_clk = 1'd0;
        left_9_7_in = 32'd0;
        left_9_7_write_en = 1'd0;
        left_9_7_clk = 1'd0;
        pe_9_8_top = 32'd0;
        pe_9_8_left = 32'd0;
        pe_9_8_go = 1'd0;
        pe_9_8_clk = 1'd0;
        top_9_8_in = 32'd0;
        top_9_8_write_en = 1'd0;
        top_9_8_clk = 1'd0;
        left_9_8_in = 32'd0;
        left_9_8_write_en = 1'd0;
        left_9_8_clk = 1'd0;
        pe_9_9_top = 32'd0;
        pe_9_9_left = 32'd0;
        pe_9_9_go = 1'd0;
        pe_9_9_clk = 1'd0;
        top_9_9_in = 32'd0;
        top_9_9_write_en = 1'd0;
        top_9_9_clk = 1'd0;
        left_9_9_in = 32'd0;
        left_9_9_write_en = 1'd0;
        left_9_9_clk = 1'd0;
        pe_9_10_top = 32'd0;
        pe_9_10_left = 32'd0;
        pe_9_10_go = 1'd0;
        pe_9_10_clk = 1'd0;
        top_9_10_in = 32'd0;
        top_9_10_write_en = 1'd0;
        top_9_10_clk = 1'd0;
        left_9_10_in = 32'd0;
        left_9_10_write_en = 1'd0;
        left_9_10_clk = 1'd0;
        pe_9_11_top = 32'd0;
        pe_9_11_left = 32'd0;
        pe_9_11_go = 1'd0;
        pe_9_11_clk = 1'd0;
        top_9_11_in = 32'd0;
        top_9_11_write_en = 1'd0;
        top_9_11_clk = 1'd0;
        left_9_11_in = 32'd0;
        left_9_11_write_en = 1'd0;
        left_9_11_clk = 1'd0;
        pe_9_12_top = 32'd0;
        pe_9_12_left = 32'd0;
        pe_9_12_go = 1'd0;
        pe_9_12_clk = 1'd0;
        top_9_12_in = 32'd0;
        top_9_12_write_en = 1'd0;
        top_9_12_clk = 1'd0;
        left_9_12_in = 32'd0;
        left_9_12_write_en = 1'd0;
        left_9_12_clk = 1'd0;
        pe_9_13_top = 32'd0;
        pe_9_13_left = 32'd0;
        pe_9_13_go = 1'd0;
        pe_9_13_clk = 1'd0;
        top_9_13_in = 32'd0;
        top_9_13_write_en = 1'd0;
        top_9_13_clk = 1'd0;
        left_9_13_in = 32'd0;
        left_9_13_write_en = 1'd0;
        left_9_13_clk = 1'd0;
        pe_9_14_top = 32'd0;
        pe_9_14_left = 32'd0;
        pe_9_14_go = 1'd0;
        pe_9_14_clk = 1'd0;
        top_9_14_in = 32'd0;
        top_9_14_write_en = 1'd0;
        top_9_14_clk = 1'd0;
        left_9_14_in = 32'd0;
        left_9_14_write_en = 1'd0;
        left_9_14_clk = 1'd0;
        pe_9_15_top = 32'd0;
        pe_9_15_left = 32'd0;
        pe_9_15_go = 1'd0;
        pe_9_15_clk = 1'd0;
        top_9_15_in = 32'd0;
        top_9_15_write_en = 1'd0;
        top_9_15_clk = 1'd0;
        left_9_15_in = 32'd0;
        left_9_15_write_en = 1'd0;
        left_9_15_clk = 1'd0;
        pe_10_0_top = 32'd0;
        pe_10_0_left = 32'd0;
        pe_10_0_go = 1'd0;
        pe_10_0_clk = 1'd0;
        top_10_0_in = 32'd0;
        top_10_0_write_en = 1'd0;
        top_10_0_clk = 1'd0;
        left_10_0_in = 32'd0;
        left_10_0_write_en = 1'd0;
        left_10_0_clk = 1'd0;
        pe_10_1_top = 32'd0;
        pe_10_1_left = 32'd0;
        pe_10_1_go = 1'd0;
        pe_10_1_clk = 1'd0;
        top_10_1_in = 32'd0;
        top_10_1_write_en = 1'd0;
        top_10_1_clk = 1'd0;
        left_10_1_in = 32'd0;
        left_10_1_write_en = 1'd0;
        left_10_1_clk = 1'd0;
        pe_10_2_top = 32'd0;
        pe_10_2_left = 32'd0;
        pe_10_2_go = 1'd0;
        pe_10_2_clk = 1'd0;
        top_10_2_in = 32'd0;
        top_10_2_write_en = 1'd0;
        top_10_2_clk = 1'd0;
        left_10_2_in = 32'd0;
        left_10_2_write_en = 1'd0;
        left_10_2_clk = 1'd0;
        pe_10_3_top = 32'd0;
        pe_10_3_left = 32'd0;
        pe_10_3_go = 1'd0;
        pe_10_3_clk = 1'd0;
        top_10_3_in = 32'd0;
        top_10_3_write_en = 1'd0;
        top_10_3_clk = 1'd0;
        left_10_3_in = 32'd0;
        left_10_3_write_en = 1'd0;
        left_10_3_clk = 1'd0;
        pe_10_4_top = 32'd0;
        pe_10_4_left = 32'd0;
        pe_10_4_go = 1'd0;
        pe_10_4_clk = 1'd0;
        top_10_4_in = 32'd0;
        top_10_4_write_en = 1'd0;
        top_10_4_clk = 1'd0;
        left_10_4_in = 32'd0;
        left_10_4_write_en = 1'd0;
        left_10_4_clk = 1'd0;
        pe_10_5_top = 32'd0;
        pe_10_5_left = 32'd0;
        pe_10_5_go = 1'd0;
        pe_10_5_clk = 1'd0;
        top_10_5_in = 32'd0;
        top_10_5_write_en = 1'd0;
        top_10_5_clk = 1'd0;
        left_10_5_in = 32'd0;
        left_10_5_write_en = 1'd0;
        left_10_5_clk = 1'd0;
        pe_10_6_top = 32'd0;
        pe_10_6_left = 32'd0;
        pe_10_6_go = 1'd0;
        pe_10_6_clk = 1'd0;
        top_10_6_in = 32'd0;
        top_10_6_write_en = 1'd0;
        top_10_6_clk = 1'd0;
        left_10_6_in = 32'd0;
        left_10_6_write_en = 1'd0;
        left_10_6_clk = 1'd0;
        pe_10_7_top = 32'd0;
        pe_10_7_left = 32'd0;
        pe_10_7_go = 1'd0;
        pe_10_7_clk = 1'd0;
        top_10_7_in = 32'd0;
        top_10_7_write_en = 1'd0;
        top_10_7_clk = 1'd0;
        left_10_7_in = 32'd0;
        left_10_7_write_en = 1'd0;
        left_10_7_clk = 1'd0;
        pe_10_8_top = 32'd0;
        pe_10_8_left = 32'd0;
        pe_10_8_go = 1'd0;
        pe_10_8_clk = 1'd0;
        top_10_8_in = 32'd0;
        top_10_8_write_en = 1'd0;
        top_10_8_clk = 1'd0;
        left_10_8_in = 32'd0;
        left_10_8_write_en = 1'd0;
        left_10_8_clk = 1'd0;
        pe_10_9_top = 32'd0;
        pe_10_9_left = 32'd0;
        pe_10_9_go = 1'd0;
        pe_10_9_clk = 1'd0;
        top_10_9_in = 32'd0;
        top_10_9_write_en = 1'd0;
        top_10_9_clk = 1'd0;
        left_10_9_in = 32'd0;
        left_10_9_write_en = 1'd0;
        left_10_9_clk = 1'd0;
        pe_10_10_top = 32'd0;
        pe_10_10_left = 32'd0;
        pe_10_10_go = 1'd0;
        pe_10_10_clk = 1'd0;
        top_10_10_in = 32'd0;
        top_10_10_write_en = 1'd0;
        top_10_10_clk = 1'd0;
        left_10_10_in = 32'd0;
        left_10_10_write_en = 1'd0;
        left_10_10_clk = 1'd0;
        pe_10_11_top = 32'd0;
        pe_10_11_left = 32'd0;
        pe_10_11_go = 1'd0;
        pe_10_11_clk = 1'd0;
        top_10_11_in = 32'd0;
        top_10_11_write_en = 1'd0;
        top_10_11_clk = 1'd0;
        left_10_11_in = 32'd0;
        left_10_11_write_en = 1'd0;
        left_10_11_clk = 1'd0;
        pe_10_12_top = 32'd0;
        pe_10_12_left = 32'd0;
        pe_10_12_go = 1'd0;
        pe_10_12_clk = 1'd0;
        top_10_12_in = 32'd0;
        top_10_12_write_en = 1'd0;
        top_10_12_clk = 1'd0;
        left_10_12_in = 32'd0;
        left_10_12_write_en = 1'd0;
        left_10_12_clk = 1'd0;
        pe_10_13_top = 32'd0;
        pe_10_13_left = 32'd0;
        pe_10_13_go = 1'd0;
        pe_10_13_clk = 1'd0;
        top_10_13_in = 32'd0;
        top_10_13_write_en = 1'd0;
        top_10_13_clk = 1'd0;
        left_10_13_in = 32'd0;
        left_10_13_write_en = 1'd0;
        left_10_13_clk = 1'd0;
        pe_10_14_top = 32'd0;
        pe_10_14_left = 32'd0;
        pe_10_14_go = 1'd0;
        pe_10_14_clk = 1'd0;
        top_10_14_in = 32'd0;
        top_10_14_write_en = 1'd0;
        top_10_14_clk = 1'd0;
        left_10_14_in = 32'd0;
        left_10_14_write_en = 1'd0;
        left_10_14_clk = 1'd0;
        pe_10_15_top = 32'd0;
        pe_10_15_left = 32'd0;
        pe_10_15_go = 1'd0;
        pe_10_15_clk = 1'd0;
        top_10_15_in = 32'd0;
        top_10_15_write_en = 1'd0;
        top_10_15_clk = 1'd0;
        left_10_15_in = 32'd0;
        left_10_15_write_en = 1'd0;
        left_10_15_clk = 1'd0;
        pe_11_0_top = 32'd0;
        pe_11_0_left = 32'd0;
        pe_11_0_go = 1'd0;
        pe_11_0_clk = 1'd0;
        top_11_0_in = 32'd0;
        top_11_0_write_en = 1'd0;
        top_11_0_clk = 1'd0;
        left_11_0_in = 32'd0;
        left_11_0_write_en = 1'd0;
        left_11_0_clk = 1'd0;
        pe_11_1_top = 32'd0;
        pe_11_1_left = 32'd0;
        pe_11_1_go = 1'd0;
        pe_11_1_clk = 1'd0;
        top_11_1_in = 32'd0;
        top_11_1_write_en = 1'd0;
        top_11_1_clk = 1'd0;
        left_11_1_in = 32'd0;
        left_11_1_write_en = 1'd0;
        left_11_1_clk = 1'd0;
        pe_11_2_top = 32'd0;
        pe_11_2_left = 32'd0;
        pe_11_2_go = 1'd0;
        pe_11_2_clk = 1'd0;
        top_11_2_in = 32'd0;
        top_11_2_write_en = 1'd0;
        top_11_2_clk = 1'd0;
        left_11_2_in = 32'd0;
        left_11_2_write_en = 1'd0;
        left_11_2_clk = 1'd0;
        pe_11_3_top = 32'd0;
        pe_11_3_left = 32'd0;
        pe_11_3_go = 1'd0;
        pe_11_3_clk = 1'd0;
        top_11_3_in = 32'd0;
        top_11_3_write_en = 1'd0;
        top_11_3_clk = 1'd0;
        left_11_3_in = 32'd0;
        left_11_3_write_en = 1'd0;
        left_11_3_clk = 1'd0;
        pe_11_4_top = 32'd0;
        pe_11_4_left = 32'd0;
        pe_11_4_go = 1'd0;
        pe_11_4_clk = 1'd0;
        top_11_4_in = 32'd0;
        top_11_4_write_en = 1'd0;
        top_11_4_clk = 1'd0;
        left_11_4_in = 32'd0;
        left_11_4_write_en = 1'd0;
        left_11_4_clk = 1'd0;
        pe_11_5_top = 32'd0;
        pe_11_5_left = 32'd0;
        pe_11_5_go = 1'd0;
        pe_11_5_clk = 1'd0;
        top_11_5_in = 32'd0;
        top_11_5_write_en = 1'd0;
        top_11_5_clk = 1'd0;
        left_11_5_in = 32'd0;
        left_11_5_write_en = 1'd0;
        left_11_5_clk = 1'd0;
        pe_11_6_top = 32'd0;
        pe_11_6_left = 32'd0;
        pe_11_6_go = 1'd0;
        pe_11_6_clk = 1'd0;
        top_11_6_in = 32'd0;
        top_11_6_write_en = 1'd0;
        top_11_6_clk = 1'd0;
        left_11_6_in = 32'd0;
        left_11_6_write_en = 1'd0;
        left_11_6_clk = 1'd0;
        pe_11_7_top = 32'd0;
        pe_11_7_left = 32'd0;
        pe_11_7_go = 1'd0;
        pe_11_7_clk = 1'd0;
        top_11_7_in = 32'd0;
        top_11_7_write_en = 1'd0;
        top_11_7_clk = 1'd0;
        left_11_7_in = 32'd0;
        left_11_7_write_en = 1'd0;
        left_11_7_clk = 1'd0;
        pe_11_8_top = 32'd0;
        pe_11_8_left = 32'd0;
        pe_11_8_go = 1'd0;
        pe_11_8_clk = 1'd0;
        top_11_8_in = 32'd0;
        top_11_8_write_en = 1'd0;
        top_11_8_clk = 1'd0;
        left_11_8_in = 32'd0;
        left_11_8_write_en = 1'd0;
        left_11_8_clk = 1'd0;
        pe_11_9_top = 32'd0;
        pe_11_9_left = 32'd0;
        pe_11_9_go = 1'd0;
        pe_11_9_clk = 1'd0;
        top_11_9_in = 32'd0;
        top_11_9_write_en = 1'd0;
        top_11_9_clk = 1'd0;
        left_11_9_in = 32'd0;
        left_11_9_write_en = 1'd0;
        left_11_9_clk = 1'd0;
        pe_11_10_top = 32'd0;
        pe_11_10_left = 32'd0;
        pe_11_10_go = 1'd0;
        pe_11_10_clk = 1'd0;
        top_11_10_in = 32'd0;
        top_11_10_write_en = 1'd0;
        top_11_10_clk = 1'd0;
        left_11_10_in = 32'd0;
        left_11_10_write_en = 1'd0;
        left_11_10_clk = 1'd0;
        pe_11_11_top = 32'd0;
        pe_11_11_left = 32'd0;
        pe_11_11_go = 1'd0;
        pe_11_11_clk = 1'd0;
        top_11_11_in = 32'd0;
        top_11_11_write_en = 1'd0;
        top_11_11_clk = 1'd0;
        left_11_11_in = 32'd0;
        left_11_11_write_en = 1'd0;
        left_11_11_clk = 1'd0;
        pe_11_12_top = 32'd0;
        pe_11_12_left = 32'd0;
        pe_11_12_go = 1'd0;
        pe_11_12_clk = 1'd0;
        top_11_12_in = 32'd0;
        top_11_12_write_en = 1'd0;
        top_11_12_clk = 1'd0;
        left_11_12_in = 32'd0;
        left_11_12_write_en = 1'd0;
        left_11_12_clk = 1'd0;
        pe_11_13_top = 32'd0;
        pe_11_13_left = 32'd0;
        pe_11_13_go = 1'd0;
        pe_11_13_clk = 1'd0;
        top_11_13_in = 32'd0;
        top_11_13_write_en = 1'd0;
        top_11_13_clk = 1'd0;
        left_11_13_in = 32'd0;
        left_11_13_write_en = 1'd0;
        left_11_13_clk = 1'd0;
        pe_11_14_top = 32'd0;
        pe_11_14_left = 32'd0;
        pe_11_14_go = 1'd0;
        pe_11_14_clk = 1'd0;
        top_11_14_in = 32'd0;
        top_11_14_write_en = 1'd0;
        top_11_14_clk = 1'd0;
        left_11_14_in = 32'd0;
        left_11_14_write_en = 1'd0;
        left_11_14_clk = 1'd0;
        pe_11_15_top = 32'd0;
        pe_11_15_left = 32'd0;
        pe_11_15_go = 1'd0;
        pe_11_15_clk = 1'd0;
        top_11_15_in = 32'd0;
        top_11_15_write_en = 1'd0;
        top_11_15_clk = 1'd0;
        left_11_15_in = 32'd0;
        left_11_15_write_en = 1'd0;
        left_11_15_clk = 1'd0;
        pe_12_0_top = 32'd0;
        pe_12_0_left = 32'd0;
        pe_12_0_go = 1'd0;
        pe_12_0_clk = 1'd0;
        top_12_0_in = 32'd0;
        top_12_0_write_en = 1'd0;
        top_12_0_clk = 1'd0;
        left_12_0_in = 32'd0;
        left_12_0_write_en = 1'd0;
        left_12_0_clk = 1'd0;
        pe_12_1_top = 32'd0;
        pe_12_1_left = 32'd0;
        pe_12_1_go = 1'd0;
        pe_12_1_clk = 1'd0;
        top_12_1_in = 32'd0;
        top_12_1_write_en = 1'd0;
        top_12_1_clk = 1'd0;
        left_12_1_in = 32'd0;
        left_12_1_write_en = 1'd0;
        left_12_1_clk = 1'd0;
        pe_12_2_top = 32'd0;
        pe_12_2_left = 32'd0;
        pe_12_2_go = 1'd0;
        pe_12_2_clk = 1'd0;
        top_12_2_in = 32'd0;
        top_12_2_write_en = 1'd0;
        top_12_2_clk = 1'd0;
        left_12_2_in = 32'd0;
        left_12_2_write_en = 1'd0;
        left_12_2_clk = 1'd0;
        pe_12_3_top = 32'd0;
        pe_12_3_left = 32'd0;
        pe_12_3_go = 1'd0;
        pe_12_3_clk = 1'd0;
        top_12_3_in = 32'd0;
        top_12_3_write_en = 1'd0;
        top_12_3_clk = 1'd0;
        left_12_3_in = 32'd0;
        left_12_3_write_en = 1'd0;
        left_12_3_clk = 1'd0;
        pe_12_4_top = 32'd0;
        pe_12_4_left = 32'd0;
        pe_12_4_go = 1'd0;
        pe_12_4_clk = 1'd0;
        top_12_4_in = 32'd0;
        top_12_4_write_en = 1'd0;
        top_12_4_clk = 1'd0;
        left_12_4_in = 32'd0;
        left_12_4_write_en = 1'd0;
        left_12_4_clk = 1'd0;
        pe_12_5_top = 32'd0;
        pe_12_5_left = 32'd0;
        pe_12_5_go = 1'd0;
        pe_12_5_clk = 1'd0;
        top_12_5_in = 32'd0;
        top_12_5_write_en = 1'd0;
        top_12_5_clk = 1'd0;
        left_12_5_in = 32'd0;
        left_12_5_write_en = 1'd0;
        left_12_5_clk = 1'd0;
        pe_12_6_top = 32'd0;
        pe_12_6_left = 32'd0;
        pe_12_6_go = 1'd0;
        pe_12_6_clk = 1'd0;
        top_12_6_in = 32'd0;
        top_12_6_write_en = 1'd0;
        top_12_6_clk = 1'd0;
        left_12_6_in = 32'd0;
        left_12_6_write_en = 1'd0;
        left_12_6_clk = 1'd0;
        pe_12_7_top = 32'd0;
        pe_12_7_left = 32'd0;
        pe_12_7_go = 1'd0;
        pe_12_7_clk = 1'd0;
        top_12_7_in = 32'd0;
        top_12_7_write_en = 1'd0;
        top_12_7_clk = 1'd0;
        left_12_7_in = 32'd0;
        left_12_7_write_en = 1'd0;
        left_12_7_clk = 1'd0;
        pe_12_8_top = 32'd0;
        pe_12_8_left = 32'd0;
        pe_12_8_go = 1'd0;
        pe_12_8_clk = 1'd0;
        top_12_8_in = 32'd0;
        top_12_8_write_en = 1'd0;
        top_12_8_clk = 1'd0;
        left_12_8_in = 32'd0;
        left_12_8_write_en = 1'd0;
        left_12_8_clk = 1'd0;
        pe_12_9_top = 32'd0;
        pe_12_9_left = 32'd0;
        pe_12_9_go = 1'd0;
        pe_12_9_clk = 1'd0;
        top_12_9_in = 32'd0;
        top_12_9_write_en = 1'd0;
        top_12_9_clk = 1'd0;
        left_12_9_in = 32'd0;
        left_12_9_write_en = 1'd0;
        left_12_9_clk = 1'd0;
        pe_12_10_top = 32'd0;
        pe_12_10_left = 32'd0;
        pe_12_10_go = 1'd0;
        pe_12_10_clk = 1'd0;
        top_12_10_in = 32'd0;
        top_12_10_write_en = 1'd0;
        top_12_10_clk = 1'd0;
        left_12_10_in = 32'd0;
        left_12_10_write_en = 1'd0;
        left_12_10_clk = 1'd0;
        pe_12_11_top = 32'd0;
        pe_12_11_left = 32'd0;
        pe_12_11_go = 1'd0;
        pe_12_11_clk = 1'd0;
        top_12_11_in = 32'd0;
        top_12_11_write_en = 1'd0;
        top_12_11_clk = 1'd0;
        left_12_11_in = 32'd0;
        left_12_11_write_en = 1'd0;
        left_12_11_clk = 1'd0;
        pe_12_12_top = 32'd0;
        pe_12_12_left = 32'd0;
        pe_12_12_go = 1'd0;
        pe_12_12_clk = 1'd0;
        top_12_12_in = 32'd0;
        top_12_12_write_en = 1'd0;
        top_12_12_clk = 1'd0;
        left_12_12_in = 32'd0;
        left_12_12_write_en = 1'd0;
        left_12_12_clk = 1'd0;
        pe_12_13_top = 32'd0;
        pe_12_13_left = 32'd0;
        pe_12_13_go = 1'd0;
        pe_12_13_clk = 1'd0;
        top_12_13_in = 32'd0;
        top_12_13_write_en = 1'd0;
        top_12_13_clk = 1'd0;
        left_12_13_in = 32'd0;
        left_12_13_write_en = 1'd0;
        left_12_13_clk = 1'd0;
        pe_12_14_top = 32'd0;
        pe_12_14_left = 32'd0;
        pe_12_14_go = 1'd0;
        pe_12_14_clk = 1'd0;
        top_12_14_in = 32'd0;
        top_12_14_write_en = 1'd0;
        top_12_14_clk = 1'd0;
        left_12_14_in = 32'd0;
        left_12_14_write_en = 1'd0;
        left_12_14_clk = 1'd0;
        pe_12_15_top = 32'd0;
        pe_12_15_left = 32'd0;
        pe_12_15_go = 1'd0;
        pe_12_15_clk = 1'd0;
        top_12_15_in = 32'd0;
        top_12_15_write_en = 1'd0;
        top_12_15_clk = 1'd0;
        left_12_15_in = 32'd0;
        left_12_15_write_en = 1'd0;
        left_12_15_clk = 1'd0;
        pe_13_0_top = 32'd0;
        pe_13_0_left = 32'd0;
        pe_13_0_go = 1'd0;
        pe_13_0_clk = 1'd0;
        top_13_0_in = 32'd0;
        top_13_0_write_en = 1'd0;
        top_13_0_clk = 1'd0;
        left_13_0_in = 32'd0;
        left_13_0_write_en = 1'd0;
        left_13_0_clk = 1'd0;
        pe_13_1_top = 32'd0;
        pe_13_1_left = 32'd0;
        pe_13_1_go = 1'd0;
        pe_13_1_clk = 1'd0;
        top_13_1_in = 32'd0;
        top_13_1_write_en = 1'd0;
        top_13_1_clk = 1'd0;
        left_13_1_in = 32'd0;
        left_13_1_write_en = 1'd0;
        left_13_1_clk = 1'd0;
        pe_13_2_top = 32'd0;
        pe_13_2_left = 32'd0;
        pe_13_2_go = 1'd0;
        pe_13_2_clk = 1'd0;
        top_13_2_in = 32'd0;
        top_13_2_write_en = 1'd0;
        top_13_2_clk = 1'd0;
        left_13_2_in = 32'd0;
        left_13_2_write_en = 1'd0;
        left_13_2_clk = 1'd0;
        pe_13_3_top = 32'd0;
        pe_13_3_left = 32'd0;
        pe_13_3_go = 1'd0;
        pe_13_3_clk = 1'd0;
        top_13_3_in = 32'd0;
        top_13_3_write_en = 1'd0;
        top_13_3_clk = 1'd0;
        left_13_3_in = 32'd0;
        left_13_3_write_en = 1'd0;
        left_13_3_clk = 1'd0;
        pe_13_4_top = 32'd0;
        pe_13_4_left = 32'd0;
        pe_13_4_go = 1'd0;
        pe_13_4_clk = 1'd0;
        top_13_4_in = 32'd0;
        top_13_4_write_en = 1'd0;
        top_13_4_clk = 1'd0;
        left_13_4_in = 32'd0;
        left_13_4_write_en = 1'd0;
        left_13_4_clk = 1'd0;
        pe_13_5_top = 32'd0;
        pe_13_5_left = 32'd0;
        pe_13_5_go = 1'd0;
        pe_13_5_clk = 1'd0;
        top_13_5_in = 32'd0;
        top_13_5_write_en = 1'd0;
        top_13_5_clk = 1'd0;
        left_13_5_in = 32'd0;
        left_13_5_write_en = 1'd0;
        left_13_5_clk = 1'd0;
        pe_13_6_top = 32'd0;
        pe_13_6_left = 32'd0;
        pe_13_6_go = 1'd0;
        pe_13_6_clk = 1'd0;
        top_13_6_in = 32'd0;
        top_13_6_write_en = 1'd0;
        top_13_6_clk = 1'd0;
        left_13_6_in = 32'd0;
        left_13_6_write_en = 1'd0;
        left_13_6_clk = 1'd0;
        pe_13_7_top = 32'd0;
        pe_13_7_left = 32'd0;
        pe_13_7_go = 1'd0;
        pe_13_7_clk = 1'd0;
        top_13_7_in = 32'd0;
        top_13_7_write_en = 1'd0;
        top_13_7_clk = 1'd0;
        left_13_7_in = 32'd0;
        left_13_7_write_en = 1'd0;
        left_13_7_clk = 1'd0;
        pe_13_8_top = 32'd0;
        pe_13_8_left = 32'd0;
        pe_13_8_go = 1'd0;
        pe_13_8_clk = 1'd0;
        top_13_8_in = 32'd0;
        top_13_8_write_en = 1'd0;
        top_13_8_clk = 1'd0;
        left_13_8_in = 32'd0;
        left_13_8_write_en = 1'd0;
        left_13_8_clk = 1'd0;
        pe_13_9_top = 32'd0;
        pe_13_9_left = 32'd0;
        pe_13_9_go = 1'd0;
        pe_13_9_clk = 1'd0;
        top_13_9_in = 32'd0;
        top_13_9_write_en = 1'd0;
        top_13_9_clk = 1'd0;
        left_13_9_in = 32'd0;
        left_13_9_write_en = 1'd0;
        left_13_9_clk = 1'd0;
        pe_13_10_top = 32'd0;
        pe_13_10_left = 32'd0;
        pe_13_10_go = 1'd0;
        pe_13_10_clk = 1'd0;
        top_13_10_in = 32'd0;
        top_13_10_write_en = 1'd0;
        top_13_10_clk = 1'd0;
        left_13_10_in = 32'd0;
        left_13_10_write_en = 1'd0;
        left_13_10_clk = 1'd0;
        pe_13_11_top = 32'd0;
        pe_13_11_left = 32'd0;
        pe_13_11_go = 1'd0;
        pe_13_11_clk = 1'd0;
        top_13_11_in = 32'd0;
        top_13_11_write_en = 1'd0;
        top_13_11_clk = 1'd0;
        left_13_11_in = 32'd0;
        left_13_11_write_en = 1'd0;
        left_13_11_clk = 1'd0;
        pe_13_12_top = 32'd0;
        pe_13_12_left = 32'd0;
        pe_13_12_go = 1'd0;
        pe_13_12_clk = 1'd0;
        top_13_12_in = 32'd0;
        top_13_12_write_en = 1'd0;
        top_13_12_clk = 1'd0;
        left_13_12_in = 32'd0;
        left_13_12_write_en = 1'd0;
        left_13_12_clk = 1'd0;
        pe_13_13_top = 32'd0;
        pe_13_13_left = 32'd0;
        pe_13_13_go = 1'd0;
        pe_13_13_clk = 1'd0;
        top_13_13_in = 32'd0;
        top_13_13_write_en = 1'd0;
        top_13_13_clk = 1'd0;
        left_13_13_in = 32'd0;
        left_13_13_write_en = 1'd0;
        left_13_13_clk = 1'd0;
        pe_13_14_top = 32'd0;
        pe_13_14_left = 32'd0;
        pe_13_14_go = 1'd0;
        pe_13_14_clk = 1'd0;
        top_13_14_in = 32'd0;
        top_13_14_write_en = 1'd0;
        top_13_14_clk = 1'd0;
        left_13_14_in = 32'd0;
        left_13_14_write_en = 1'd0;
        left_13_14_clk = 1'd0;
        pe_13_15_top = 32'd0;
        pe_13_15_left = 32'd0;
        pe_13_15_go = 1'd0;
        pe_13_15_clk = 1'd0;
        top_13_15_in = 32'd0;
        top_13_15_write_en = 1'd0;
        top_13_15_clk = 1'd0;
        left_13_15_in = 32'd0;
        left_13_15_write_en = 1'd0;
        left_13_15_clk = 1'd0;
        pe_14_0_top = 32'd0;
        pe_14_0_left = 32'd0;
        pe_14_0_go = 1'd0;
        pe_14_0_clk = 1'd0;
        top_14_0_in = 32'd0;
        top_14_0_write_en = 1'd0;
        top_14_0_clk = 1'd0;
        left_14_0_in = 32'd0;
        left_14_0_write_en = 1'd0;
        left_14_0_clk = 1'd0;
        pe_14_1_top = 32'd0;
        pe_14_1_left = 32'd0;
        pe_14_1_go = 1'd0;
        pe_14_1_clk = 1'd0;
        top_14_1_in = 32'd0;
        top_14_1_write_en = 1'd0;
        top_14_1_clk = 1'd0;
        left_14_1_in = 32'd0;
        left_14_1_write_en = 1'd0;
        left_14_1_clk = 1'd0;
        pe_14_2_top = 32'd0;
        pe_14_2_left = 32'd0;
        pe_14_2_go = 1'd0;
        pe_14_2_clk = 1'd0;
        top_14_2_in = 32'd0;
        top_14_2_write_en = 1'd0;
        top_14_2_clk = 1'd0;
        left_14_2_in = 32'd0;
        left_14_2_write_en = 1'd0;
        left_14_2_clk = 1'd0;
        pe_14_3_top = 32'd0;
        pe_14_3_left = 32'd0;
        pe_14_3_go = 1'd0;
        pe_14_3_clk = 1'd0;
        top_14_3_in = 32'd0;
        top_14_3_write_en = 1'd0;
        top_14_3_clk = 1'd0;
        left_14_3_in = 32'd0;
        left_14_3_write_en = 1'd0;
        left_14_3_clk = 1'd0;
        pe_14_4_top = 32'd0;
        pe_14_4_left = 32'd0;
        pe_14_4_go = 1'd0;
        pe_14_4_clk = 1'd0;
        top_14_4_in = 32'd0;
        top_14_4_write_en = 1'd0;
        top_14_4_clk = 1'd0;
        left_14_4_in = 32'd0;
        left_14_4_write_en = 1'd0;
        left_14_4_clk = 1'd0;
        pe_14_5_top = 32'd0;
        pe_14_5_left = 32'd0;
        pe_14_5_go = 1'd0;
        pe_14_5_clk = 1'd0;
        top_14_5_in = 32'd0;
        top_14_5_write_en = 1'd0;
        top_14_5_clk = 1'd0;
        left_14_5_in = 32'd0;
        left_14_5_write_en = 1'd0;
        left_14_5_clk = 1'd0;
        pe_14_6_top = 32'd0;
        pe_14_6_left = 32'd0;
        pe_14_6_go = 1'd0;
        pe_14_6_clk = 1'd0;
        top_14_6_in = 32'd0;
        top_14_6_write_en = 1'd0;
        top_14_6_clk = 1'd0;
        left_14_6_in = 32'd0;
        left_14_6_write_en = 1'd0;
        left_14_6_clk = 1'd0;
        pe_14_7_top = 32'd0;
        pe_14_7_left = 32'd0;
        pe_14_7_go = 1'd0;
        pe_14_7_clk = 1'd0;
        top_14_7_in = 32'd0;
        top_14_7_write_en = 1'd0;
        top_14_7_clk = 1'd0;
        left_14_7_in = 32'd0;
        left_14_7_write_en = 1'd0;
        left_14_7_clk = 1'd0;
        pe_14_8_top = 32'd0;
        pe_14_8_left = 32'd0;
        pe_14_8_go = 1'd0;
        pe_14_8_clk = 1'd0;
        top_14_8_in = 32'd0;
        top_14_8_write_en = 1'd0;
        top_14_8_clk = 1'd0;
        left_14_8_in = 32'd0;
        left_14_8_write_en = 1'd0;
        left_14_8_clk = 1'd0;
        pe_14_9_top = 32'd0;
        pe_14_9_left = 32'd0;
        pe_14_9_go = 1'd0;
        pe_14_9_clk = 1'd0;
        top_14_9_in = 32'd0;
        top_14_9_write_en = 1'd0;
        top_14_9_clk = 1'd0;
        left_14_9_in = 32'd0;
        left_14_9_write_en = 1'd0;
        left_14_9_clk = 1'd0;
        pe_14_10_top = 32'd0;
        pe_14_10_left = 32'd0;
        pe_14_10_go = 1'd0;
        pe_14_10_clk = 1'd0;
        top_14_10_in = 32'd0;
        top_14_10_write_en = 1'd0;
        top_14_10_clk = 1'd0;
        left_14_10_in = 32'd0;
        left_14_10_write_en = 1'd0;
        left_14_10_clk = 1'd0;
        pe_14_11_top = 32'd0;
        pe_14_11_left = 32'd0;
        pe_14_11_go = 1'd0;
        pe_14_11_clk = 1'd0;
        top_14_11_in = 32'd0;
        top_14_11_write_en = 1'd0;
        top_14_11_clk = 1'd0;
        left_14_11_in = 32'd0;
        left_14_11_write_en = 1'd0;
        left_14_11_clk = 1'd0;
        pe_14_12_top = 32'd0;
        pe_14_12_left = 32'd0;
        pe_14_12_go = 1'd0;
        pe_14_12_clk = 1'd0;
        top_14_12_in = 32'd0;
        top_14_12_write_en = 1'd0;
        top_14_12_clk = 1'd0;
        left_14_12_in = 32'd0;
        left_14_12_write_en = 1'd0;
        left_14_12_clk = 1'd0;
        pe_14_13_top = 32'd0;
        pe_14_13_left = 32'd0;
        pe_14_13_go = 1'd0;
        pe_14_13_clk = 1'd0;
        top_14_13_in = 32'd0;
        top_14_13_write_en = 1'd0;
        top_14_13_clk = 1'd0;
        left_14_13_in = 32'd0;
        left_14_13_write_en = 1'd0;
        left_14_13_clk = 1'd0;
        pe_14_14_top = 32'd0;
        pe_14_14_left = 32'd0;
        pe_14_14_go = 1'd0;
        pe_14_14_clk = 1'd0;
        top_14_14_in = 32'd0;
        top_14_14_write_en = 1'd0;
        top_14_14_clk = 1'd0;
        left_14_14_in = 32'd0;
        left_14_14_write_en = 1'd0;
        left_14_14_clk = 1'd0;
        pe_14_15_top = 32'd0;
        pe_14_15_left = 32'd0;
        pe_14_15_go = 1'd0;
        pe_14_15_clk = 1'd0;
        top_14_15_in = 32'd0;
        top_14_15_write_en = 1'd0;
        top_14_15_clk = 1'd0;
        left_14_15_in = 32'd0;
        left_14_15_write_en = 1'd0;
        left_14_15_clk = 1'd0;
        pe_15_0_top = 32'd0;
        pe_15_0_left = 32'd0;
        pe_15_0_go = 1'd0;
        pe_15_0_clk = 1'd0;
        top_15_0_in = 32'd0;
        top_15_0_write_en = 1'd0;
        top_15_0_clk = 1'd0;
        left_15_0_in = 32'd0;
        left_15_0_write_en = 1'd0;
        left_15_0_clk = 1'd0;
        pe_15_1_top = 32'd0;
        pe_15_1_left = 32'd0;
        pe_15_1_go = 1'd0;
        pe_15_1_clk = 1'd0;
        top_15_1_in = 32'd0;
        top_15_1_write_en = 1'd0;
        top_15_1_clk = 1'd0;
        left_15_1_in = 32'd0;
        left_15_1_write_en = 1'd0;
        left_15_1_clk = 1'd0;
        pe_15_2_top = 32'd0;
        pe_15_2_left = 32'd0;
        pe_15_2_go = 1'd0;
        pe_15_2_clk = 1'd0;
        top_15_2_in = 32'd0;
        top_15_2_write_en = 1'd0;
        top_15_2_clk = 1'd0;
        left_15_2_in = 32'd0;
        left_15_2_write_en = 1'd0;
        left_15_2_clk = 1'd0;
        pe_15_3_top = 32'd0;
        pe_15_3_left = 32'd0;
        pe_15_3_go = 1'd0;
        pe_15_3_clk = 1'd0;
        top_15_3_in = 32'd0;
        top_15_3_write_en = 1'd0;
        top_15_3_clk = 1'd0;
        left_15_3_in = 32'd0;
        left_15_3_write_en = 1'd0;
        left_15_3_clk = 1'd0;
        pe_15_4_top = 32'd0;
        pe_15_4_left = 32'd0;
        pe_15_4_go = 1'd0;
        pe_15_4_clk = 1'd0;
        top_15_4_in = 32'd0;
        top_15_4_write_en = 1'd0;
        top_15_4_clk = 1'd0;
        left_15_4_in = 32'd0;
        left_15_4_write_en = 1'd0;
        left_15_4_clk = 1'd0;
        pe_15_5_top = 32'd0;
        pe_15_5_left = 32'd0;
        pe_15_5_go = 1'd0;
        pe_15_5_clk = 1'd0;
        top_15_5_in = 32'd0;
        top_15_5_write_en = 1'd0;
        top_15_5_clk = 1'd0;
        left_15_5_in = 32'd0;
        left_15_5_write_en = 1'd0;
        left_15_5_clk = 1'd0;
        pe_15_6_top = 32'd0;
        pe_15_6_left = 32'd0;
        pe_15_6_go = 1'd0;
        pe_15_6_clk = 1'd0;
        top_15_6_in = 32'd0;
        top_15_6_write_en = 1'd0;
        top_15_6_clk = 1'd0;
        left_15_6_in = 32'd0;
        left_15_6_write_en = 1'd0;
        left_15_6_clk = 1'd0;
        pe_15_7_top = 32'd0;
        pe_15_7_left = 32'd0;
        pe_15_7_go = 1'd0;
        pe_15_7_clk = 1'd0;
        top_15_7_in = 32'd0;
        top_15_7_write_en = 1'd0;
        top_15_7_clk = 1'd0;
        left_15_7_in = 32'd0;
        left_15_7_write_en = 1'd0;
        left_15_7_clk = 1'd0;
        pe_15_8_top = 32'd0;
        pe_15_8_left = 32'd0;
        pe_15_8_go = 1'd0;
        pe_15_8_clk = 1'd0;
        top_15_8_in = 32'd0;
        top_15_8_write_en = 1'd0;
        top_15_8_clk = 1'd0;
        left_15_8_in = 32'd0;
        left_15_8_write_en = 1'd0;
        left_15_8_clk = 1'd0;
        pe_15_9_top = 32'd0;
        pe_15_9_left = 32'd0;
        pe_15_9_go = 1'd0;
        pe_15_9_clk = 1'd0;
        top_15_9_in = 32'd0;
        top_15_9_write_en = 1'd0;
        top_15_9_clk = 1'd0;
        left_15_9_in = 32'd0;
        left_15_9_write_en = 1'd0;
        left_15_9_clk = 1'd0;
        pe_15_10_top = 32'd0;
        pe_15_10_left = 32'd0;
        pe_15_10_go = 1'd0;
        pe_15_10_clk = 1'd0;
        top_15_10_in = 32'd0;
        top_15_10_write_en = 1'd0;
        top_15_10_clk = 1'd0;
        left_15_10_in = 32'd0;
        left_15_10_write_en = 1'd0;
        left_15_10_clk = 1'd0;
        pe_15_11_top = 32'd0;
        pe_15_11_left = 32'd0;
        pe_15_11_go = 1'd0;
        pe_15_11_clk = 1'd0;
        top_15_11_in = 32'd0;
        top_15_11_write_en = 1'd0;
        top_15_11_clk = 1'd0;
        left_15_11_in = 32'd0;
        left_15_11_write_en = 1'd0;
        left_15_11_clk = 1'd0;
        pe_15_12_top = 32'd0;
        pe_15_12_left = 32'd0;
        pe_15_12_go = 1'd0;
        pe_15_12_clk = 1'd0;
        top_15_12_in = 32'd0;
        top_15_12_write_en = 1'd0;
        top_15_12_clk = 1'd0;
        left_15_12_in = 32'd0;
        left_15_12_write_en = 1'd0;
        left_15_12_clk = 1'd0;
        pe_15_13_top = 32'd0;
        pe_15_13_left = 32'd0;
        pe_15_13_go = 1'd0;
        pe_15_13_clk = 1'd0;
        top_15_13_in = 32'd0;
        top_15_13_write_en = 1'd0;
        top_15_13_clk = 1'd0;
        left_15_13_in = 32'd0;
        left_15_13_write_en = 1'd0;
        left_15_13_clk = 1'd0;
        pe_15_14_top = 32'd0;
        pe_15_14_left = 32'd0;
        pe_15_14_go = 1'd0;
        pe_15_14_clk = 1'd0;
        top_15_14_in = 32'd0;
        top_15_14_write_en = 1'd0;
        top_15_14_clk = 1'd0;
        left_15_14_in = 32'd0;
        left_15_14_write_en = 1'd0;
        left_15_14_clk = 1'd0;
        pe_15_15_top = 32'd0;
        pe_15_15_left = 32'd0;
        pe_15_15_go = 1'd0;
        pe_15_15_clk = 1'd0;
        top_15_15_in = 32'd0;
        top_15_15_write_en = 1'd0;
        top_15_15_clk = 1'd0;
        left_15_15_in = 32'd0;
        left_15_15_write_en = 1'd0;
        left_15_15_clk = 1'd0;
        fsm_in = 1'd0;
        fsm_write_en = 1'd0;
        fsm_clk = 1'd0;
        incr_left = 1'd0;
        incr_right = 1'd0;
        fsm0_in = 1'd0;
        fsm0_write_en = 1'd0;
        fsm0_clk = 1'd0;
        incr0_left = 1'd0;
        incr0_right = 1'd0;
        fsm1_in = 1'd0;
        fsm1_write_en = 1'd0;
        fsm1_clk = 1'd0;
        incr1_left = 1'd0;
        incr1_right = 1'd0;
        fsm2_in = 3'd0;
        fsm2_write_en = 1'd0;
        fsm2_clk = 1'd0;
        incr2_left = 3'd0;
        incr2_right = 3'd0;
        fsm3_in = 1'd0;
        fsm3_write_en = 1'd0;
        fsm3_clk = 1'd0;
        incr3_left = 1'd0;
        incr3_right = 1'd0;
        fsm4_in = 3'd0;
        fsm4_write_en = 1'd0;
        fsm4_clk = 1'd0;
        incr4_left = 3'd0;
        incr4_right = 3'd0;
        fsm5_in = 1'd0;
        fsm5_write_en = 1'd0;
        fsm5_clk = 1'd0;
        incr5_left = 1'd0;
        incr5_right = 1'd0;
        fsm6_in = 3'd0;
        fsm6_write_en = 1'd0;
        fsm6_clk = 1'd0;
        incr6_left = 3'd0;
        incr6_right = 3'd0;
        fsm7_in = 1'd0;
        fsm7_write_en = 1'd0;
        fsm7_clk = 1'd0;
        incr7_left = 1'd0;
        incr7_right = 1'd0;
        fsm8_in = 3'd0;
        fsm8_write_en = 1'd0;
        fsm8_clk = 1'd0;
        incr8_left = 3'd0;
        incr8_right = 3'd0;
        fsm9_in = 1'd0;
        fsm9_write_en = 1'd0;
        fsm9_clk = 1'd0;
        incr9_left = 1'd0;
        incr9_right = 1'd0;
        fsm10_in = 3'd0;
        fsm10_write_en = 1'd0;
        fsm10_clk = 1'd0;
        incr10_left = 3'd0;
        incr10_right = 3'd0;
        fsm11_in = 1'd0;
        fsm11_write_en = 1'd0;
        fsm11_clk = 1'd0;
        incr11_left = 1'd0;
        incr11_right = 1'd0;
        fsm12_in = 3'd0;
        fsm12_write_en = 1'd0;
        fsm12_clk = 1'd0;
        incr12_left = 3'd0;
        incr12_right = 3'd0;
        fsm13_in = 1'd0;
        fsm13_write_en = 1'd0;
        fsm13_clk = 1'd0;
        incr13_left = 1'd0;
        incr13_right = 1'd0;
        fsm14_in = 3'd0;
        fsm14_write_en = 1'd0;
        fsm14_clk = 1'd0;
        incr14_left = 3'd0;
        incr14_right = 3'd0;
        fsm15_in = 1'd0;
        fsm15_write_en = 1'd0;
        fsm15_clk = 1'd0;
        incr15_left = 1'd0;
        incr15_right = 1'd0;
        fsm16_in = 3'd0;
        fsm16_write_en = 1'd0;
        fsm16_clk = 1'd0;
        incr16_left = 3'd0;
        incr16_right = 3'd0;
        fsm17_in = 1'd0;
        fsm17_write_en = 1'd0;
        fsm17_clk = 1'd0;
        incr17_left = 1'd0;
        incr17_right = 1'd0;
        fsm18_in = 3'd0;
        fsm18_write_en = 1'd0;
        fsm18_clk = 1'd0;
        incr18_left = 3'd0;
        incr18_right = 3'd0;
        fsm19_in = 1'd0;
        fsm19_write_en = 1'd0;
        fsm19_clk = 1'd0;
        incr19_left = 1'd0;
        incr19_right = 1'd0;
        fsm20_in = 3'd0;
        fsm20_write_en = 1'd0;
        fsm20_clk = 1'd0;
        incr20_left = 3'd0;
        incr20_right = 3'd0;
        fsm21_in = 1'd0;
        fsm21_write_en = 1'd0;
        fsm21_clk = 1'd0;
        incr21_left = 1'd0;
        incr21_right = 1'd0;
        fsm22_in = 3'd0;
        fsm22_write_en = 1'd0;
        fsm22_clk = 1'd0;
        incr22_left = 3'd0;
        incr22_right = 3'd0;
        fsm23_in = 1'd0;
        fsm23_write_en = 1'd0;
        fsm23_clk = 1'd0;
        incr23_left = 1'd0;
        incr23_right = 1'd0;
        fsm24_in = 3'd0;
        fsm24_write_en = 1'd0;
        fsm24_clk = 1'd0;
        incr24_left = 3'd0;
        incr24_right = 3'd0;
        fsm25_in = 1'd0;
        fsm25_write_en = 1'd0;
        fsm25_clk = 1'd0;
        incr25_left = 1'd0;
        incr25_right = 1'd0;
        fsm26_in = 3'd0;
        fsm26_write_en = 1'd0;
        fsm26_clk = 1'd0;
        incr26_left = 3'd0;
        incr26_right = 3'd0;
        fsm27_in = 1'd0;
        fsm27_write_en = 1'd0;
        fsm27_clk = 1'd0;
        incr27_left = 1'd0;
        incr27_right = 1'd0;
        fsm28_in = 3'd0;
        fsm28_write_en = 1'd0;
        fsm28_clk = 1'd0;
        incr28_left = 3'd0;
        incr28_right = 3'd0;
        fsm29_in = 1'd0;
        fsm29_write_en = 1'd0;
        fsm29_clk = 1'd0;
        incr29_left = 1'd0;
        incr29_right = 1'd0;
        fsm30_in = 3'd0;
        fsm30_write_en = 1'd0;
        fsm30_clk = 1'd0;
        incr30_left = 3'd0;
        incr30_right = 3'd0;
        fsm31_in = 1'd0;
        fsm31_write_en = 1'd0;
        fsm31_clk = 1'd0;
        incr31_left = 1'd0;
        incr31_right = 1'd0;
        fsm32_in = 3'd0;
        fsm32_write_en = 1'd0;
        fsm32_clk = 1'd0;
        incr32_left = 3'd0;
        incr32_right = 3'd0;
        fsm33_in = 1'd0;
        fsm33_write_en = 1'd0;
        fsm33_clk = 1'd0;
        incr33_left = 1'd0;
        incr33_right = 1'd0;
        fsm34_in = 3'd0;
        fsm34_write_en = 1'd0;
        fsm34_clk = 1'd0;
        incr34_left = 3'd0;
        incr34_right = 3'd0;
        fsm35_in = 1'd0;
        fsm35_write_en = 1'd0;
        fsm35_clk = 1'd0;
        incr35_left = 1'd0;
        incr35_right = 1'd0;
        fsm36_in = 3'd0;
        fsm36_write_en = 1'd0;
        fsm36_clk = 1'd0;
        incr36_left = 3'd0;
        incr36_right = 3'd0;
        fsm37_in = 1'd0;
        fsm37_write_en = 1'd0;
        fsm37_clk = 1'd0;
        incr37_left = 1'd0;
        incr37_right = 1'd0;
        fsm38_in = 3'd0;
        fsm38_write_en = 1'd0;
        fsm38_clk = 1'd0;
        incr38_left = 3'd0;
        incr38_right = 3'd0;
        fsm39_in = 1'd0;
        fsm39_write_en = 1'd0;
        fsm39_clk = 1'd0;
        incr39_left = 1'd0;
        incr39_right = 1'd0;
        fsm40_in = 3'd0;
        fsm40_write_en = 1'd0;
        fsm40_clk = 1'd0;
        incr40_left = 3'd0;
        incr40_right = 3'd0;
        fsm41_in = 1'd0;
        fsm41_write_en = 1'd0;
        fsm41_clk = 1'd0;
        incr41_left = 1'd0;
        incr41_right = 1'd0;
        fsm42_in = 3'd0;
        fsm42_write_en = 1'd0;
        fsm42_clk = 1'd0;
        incr42_left = 3'd0;
        incr42_right = 3'd0;
        fsm43_in = 1'd0;
        fsm43_write_en = 1'd0;
        fsm43_clk = 1'd0;
        incr43_left = 1'd0;
        incr43_right = 1'd0;
        fsm44_in = 3'd0;
        fsm44_write_en = 1'd0;
        fsm44_clk = 1'd0;
        incr44_left = 3'd0;
        incr44_right = 3'd0;
        fsm45_in = 1'd0;
        fsm45_write_en = 1'd0;
        fsm45_clk = 1'd0;
        incr45_left = 1'd0;
        incr45_right = 1'd0;
        fsm46_in = 3'd0;
        fsm46_write_en = 1'd0;
        fsm46_clk = 1'd0;
        incr46_left = 3'd0;
        incr46_right = 3'd0;
        fsm47_in = 1'd0;
        fsm47_write_en = 1'd0;
        fsm47_clk = 1'd0;
        incr47_left = 1'd0;
        incr47_right = 1'd0;
        fsm48_in = 3'd0;
        fsm48_write_en = 1'd0;
        fsm48_clk = 1'd0;
        incr48_left = 3'd0;
        incr48_right = 3'd0;
        fsm49_in = 1'd0;
        fsm49_write_en = 1'd0;
        fsm49_clk = 1'd0;
        incr49_left = 1'd0;
        incr49_right = 1'd0;
        fsm50_in = 3'd0;
        fsm50_write_en = 1'd0;
        fsm50_clk = 1'd0;
        incr50_left = 3'd0;
        incr50_right = 3'd0;
        fsm51_in = 1'd0;
        fsm51_write_en = 1'd0;
        fsm51_clk = 1'd0;
        incr51_left = 1'd0;
        incr51_right = 1'd0;
        fsm52_in = 3'd0;
        fsm52_write_en = 1'd0;
        fsm52_clk = 1'd0;
        incr52_left = 3'd0;
        incr52_right = 3'd0;
        fsm53_in = 1'd0;
        fsm53_write_en = 1'd0;
        fsm53_clk = 1'd0;
        incr53_left = 1'd0;
        incr53_right = 1'd0;
        fsm54_in = 3'd0;
        fsm54_write_en = 1'd0;
        fsm54_clk = 1'd0;
        incr54_left = 3'd0;
        incr54_right = 3'd0;
        fsm55_in = 1'd0;
        fsm55_write_en = 1'd0;
        fsm55_clk = 1'd0;
        incr55_left = 1'd0;
        incr55_right = 1'd0;
        fsm56_in = 3'd0;
        fsm56_write_en = 1'd0;
        fsm56_clk = 1'd0;
        incr56_left = 3'd0;
        incr56_right = 3'd0;
        fsm57_in = 1'd0;
        fsm57_write_en = 1'd0;
        fsm57_clk = 1'd0;
        incr57_left = 1'd0;
        incr57_right = 1'd0;
        fsm58_in = 3'd0;
        fsm58_write_en = 1'd0;
        fsm58_clk = 1'd0;
        incr58_left = 3'd0;
        incr58_right = 3'd0;
        fsm59_in = 1'd0;
        fsm59_write_en = 1'd0;
        fsm59_clk = 1'd0;
        incr59_left = 1'd0;
        incr59_right = 1'd0;
        fsm60_in = 3'd0;
        fsm60_write_en = 1'd0;
        fsm60_clk = 1'd0;
        incr60_left = 3'd0;
        incr60_right = 3'd0;
        fsm61_in = 1'd0;
        fsm61_write_en = 1'd0;
        fsm61_clk = 1'd0;
        incr61_left = 1'd0;
        incr61_right = 1'd0;
        fsm62_in = 3'd0;
        fsm62_write_en = 1'd0;
        fsm62_clk = 1'd0;
        incr62_left = 3'd0;
        incr62_right = 3'd0;
        fsm63_in = 1'd0;
        fsm63_write_en = 1'd0;
        fsm63_clk = 1'd0;
        incr63_left = 1'd0;
        incr63_right = 1'd0;
        fsm64_in = 3'd0;
        fsm64_write_en = 1'd0;
        fsm64_clk = 1'd0;
        incr64_left = 3'd0;
        incr64_right = 3'd0;
        fsm65_in = 1'd0;
        fsm65_write_en = 1'd0;
        fsm65_clk = 1'd0;
        incr65_left = 1'd0;
        incr65_right = 1'd0;
        fsm66_in = 3'd0;
        fsm66_write_en = 1'd0;
        fsm66_clk = 1'd0;
        incr66_left = 3'd0;
        incr66_right = 3'd0;
        fsm67_in = 1'd0;
        fsm67_write_en = 1'd0;
        fsm67_clk = 1'd0;
        incr67_left = 1'd0;
        incr67_right = 1'd0;
        fsm68_in = 3'd0;
        fsm68_write_en = 1'd0;
        fsm68_clk = 1'd0;
        incr68_left = 3'd0;
        incr68_right = 3'd0;
        fsm69_in = 1'd0;
        fsm69_write_en = 1'd0;
        fsm69_clk = 1'd0;
        incr69_left = 1'd0;
        incr69_right = 1'd0;
        fsm70_in = 3'd0;
        fsm70_write_en = 1'd0;
        fsm70_clk = 1'd0;
        incr70_left = 3'd0;
        incr70_right = 3'd0;
        fsm71_in = 1'd0;
        fsm71_write_en = 1'd0;
        fsm71_clk = 1'd0;
        incr71_left = 1'd0;
        incr71_right = 1'd0;
        fsm72_in = 3'd0;
        fsm72_write_en = 1'd0;
        fsm72_clk = 1'd0;
        incr72_left = 3'd0;
        incr72_right = 3'd0;
        fsm73_in = 1'd0;
        fsm73_write_en = 1'd0;
        fsm73_clk = 1'd0;
        incr73_left = 1'd0;
        incr73_right = 1'd0;
        fsm74_in = 3'd0;
        fsm74_write_en = 1'd0;
        fsm74_clk = 1'd0;
        incr74_left = 3'd0;
        incr74_right = 3'd0;
        fsm75_in = 1'd0;
        fsm75_write_en = 1'd0;
        fsm75_clk = 1'd0;
        incr75_left = 1'd0;
        incr75_right = 1'd0;
        fsm76_in = 3'd0;
        fsm76_write_en = 1'd0;
        fsm76_clk = 1'd0;
        incr76_left = 3'd0;
        incr76_right = 3'd0;
        fsm77_in = 1'd0;
        fsm77_write_en = 1'd0;
        fsm77_clk = 1'd0;
        incr77_left = 1'd0;
        incr77_right = 1'd0;
        fsm78_in = 3'd0;
        fsm78_write_en = 1'd0;
        fsm78_clk = 1'd0;
        incr78_left = 3'd0;
        incr78_right = 3'd0;
        fsm79_in = 1'd0;
        fsm79_write_en = 1'd0;
        fsm79_clk = 1'd0;
        incr79_left = 1'd0;
        incr79_right = 1'd0;
        fsm80_in = 3'd0;
        fsm80_write_en = 1'd0;
        fsm80_clk = 1'd0;
        incr80_left = 3'd0;
        incr80_right = 3'd0;
        fsm81_in = 1'd0;
        fsm81_write_en = 1'd0;
        fsm81_clk = 1'd0;
        incr81_left = 1'd0;
        incr81_right = 1'd0;
        fsm82_in = 3'd0;
        fsm82_write_en = 1'd0;
        fsm82_clk = 1'd0;
        incr82_left = 3'd0;
        incr82_right = 3'd0;
        fsm83_in = 1'd0;
        fsm83_write_en = 1'd0;
        fsm83_clk = 1'd0;
        incr83_left = 1'd0;
        incr83_right = 1'd0;
        fsm84_in = 3'd0;
        fsm84_write_en = 1'd0;
        fsm84_clk = 1'd0;
        incr84_left = 3'd0;
        incr84_right = 3'd0;
        fsm85_in = 1'd0;
        fsm85_write_en = 1'd0;
        fsm85_clk = 1'd0;
        incr85_left = 1'd0;
        incr85_right = 1'd0;
        fsm86_in = 3'd0;
        fsm86_write_en = 1'd0;
        fsm86_clk = 1'd0;
        incr86_left = 3'd0;
        incr86_right = 3'd0;
        fsm87_in = 1'd0;
        fsm87_write_en = 1'd0;
        fsm87_clk = 1'd0;
        incr87_left = 1'd0;
        incr87_right = 1'd0;
        fsm88_in = 3'd0;
        fsm88_write_en = 1'd0;
        fsm88_clk = 1'd0;
        incr88_left = 3'd0;
        incr88_right = 3'd0;
        fsm89_in = 1'd0;
        fsm89_write_en = 1'd0;
        fsm89_clk = 1'd0;
        incr89_left = 1'd0;
        incr89_right = 1'd0;
        fsm90_in = 3'd0;
        fsm90_write_en = 1'd0;
        fsm90_clk = 1'd0;
        incr90_left = 3'd0;
        incr90_right = 3'd0;
        fsm91_in = 1'd0;
        fsm91_write_en = 1'd0;
        fsm91_clk = 1'd0;
        incr91_left = 1'd0;
        incr91_right = 1'd0;
        fsm92_in = 10'd0;
        fsm92_write_en = 1'd0;
        fsm92_clk = 1'd0;
        incr92_left = 10'd0;
        incr92_right = 10'd0;
    end
    std_reg # (
        .width(5)
    ) t0_idx (
        .clk(t0_idx_clk),
        .done(t0_idx_done),
        .in(t0_idx_in),
        .out(t0_idx_out),
        .write_en(t0_idx_write_en)
    );
    std_add # (
        .width(5)
    ) t0_add (
        .left(t0_add_left),
        .out(t0_add_out),
        .right(t0_add_right)
    );
    std_reg # (
        .width(5)
    ) t1_idx (
        .clk(t1_idx_clk),
        .done(t1_idx_done),
        .in(t1_idx_in),
        .out(t1_idx_out),
        .write_en(t1_idx_write_en)
    );
    std_add # (
        .width(5)
    ) t1_add (
        .left(t1_add_left),
        .out(t1_add_out),
        .right(t1_add_right)
    );
    std_reg # (
        .width(5)
    ) t2_idx (
        .clk(t2_idx_clk),
        .done(t2_idx_done),
        .in(t2_idx_in),
        .out(t2_idx_out),
        .write_en(t2_idx_write_en)
    );
    std_add # (
        .width(5)
    ) t2_add (
        .left(t2_add_left),
        .out(t2_add_out),
        .right(t2_add_right)
    );
    std_reg # (
        .width(5)
    ) t3_idx (
        .clk(t3_idx_clk),
        .done(t3_idx_done),
        .in(t3_idx_in),
        .out(t3_idx_out),
        .write_en(t3_idx_write_en)
    );
    std_add # (
        .width(5)
    ) t3_add (
        .left(t3_add_left),
        .out(t3_add_out),
        .right(t3_add_right)
    );
    std_reg # (
        .width(5)
    ) t4_idx (
        .clk(t4_idx_clk),
        .done(t4_idx_done),
        .in(t4_idx_in),
        .out(t4_idx_out),
        .write_en(t4_idx_write_en)
    );
    std_add # (
        .width(5)
    ) t4_add (
        .left(t4_add_left),
        .out(t4_add_out),
        .right(t4_add_right)
    );
    std_reg # (
        .width(5)
    ) t5_idx (
        .clk(t5_idx_clk),
        .done(t5_idx_done),
        .in(t5_idx_in),
        .out(t5_idx_out),
        .write_en(t5_idx_write_en)
    );
    std_add # (
        .width(5)
    ) t5_add (
        .left(t5_add_left),
        .out(t5_add_out),
        .right(t5_add_right)
    );
    std_reg # (
        .width(5)
    ) t6_idx (
        .clk(t6_idx_clk),
        .done(t6_idx_done),
        .in(t6_idx_in),
        .out(t6_idx_out),
        .write_en(t6_idx_write_en)
    );
    std_add # (
        .width(5)
    ) t6_add (
        .left(t6_add_left),
        .out(t6_add_out),
        .right(t6_add_right)
    );
    std_reg # (
        .width(5)
    ) t7_idx (
        .clk(t7_idx_clk),
        .done(t7_idx_done),
        .in(t7_idx_in),
        .out(t7_idx_out),
        .write_en(t7_idx_write_en)
    );
    std_add # (
        .width(5)
    ) t7_add (
        .left(t7_add_left),
        .out(t7_add_out),
        .right(t7_add_right)
    );
    std_reg # (
        .width(5)
    ) t8_idx (
        .clk(t8_idx_clk),
        .done(t8_idx_done),
        .in(t8_idx_in),
        .out(t8_idx_out),
        .write_en(t8_idx_write_en)
    );
    std_add # (
        .width(5)
    ) t8_add (
        .left(t8_add_left),
        .out(t8_add_out),
        .right(t8_add_right)
    );
    std_reg # (
        .width(5)
    ) t9_idx (
        .clk(t9_idx_clk),
        .done(t9_idx_done),
        .in(t9_idx_in),
        .out(t9_idx_out),
        .write_en(t9_idx_write_en)
    );
    std_add # (
        .width(5)
    ) t9_add (
        .left(t9_add_left),
        .out(t9_add_out),
        .right(t9_add_right)
    );
    std_reg # (
        .width(5)
    ) t10_idx (
        .clk(t10_idx_clk),
        .done(t10_idx_done),
        .in(t10_idx_in),
        .out(t10_idx_out),
        .write_en(t10_idx_write_en)
    );
    std_add # (
        .width(5)
    ) t10_add (
        .left(t10_add_left),
        .out(t10_add_out),
        .right(t10_add_right)
    );
    std_reg # (
        .width(5)
    ) t11_idx (
        .clk(t11_idx_clk),
        .done(t11_idx_done),
        .in(t11_idx_in),
        .out(t11_idx_out),
        .write_en(t11_idx_write_en)
    );
    std_add # (
        .width(5)
    ) t11_add (
        .left(t11_add_left),
        .out(t11_add_out),
        .right(t11_add_right)
    );
    std_reg # (
        .width(5)
    ) t12_idx (
        .clk(t12_idx_clk),
        .done(t12_idx_done),
        .in(t12_idx_in),
        .out(t12_idx_out),
        .write_en(t12_idx_write_en)
    );
    std_add # (
        .width(5)
    ) t12_add (
        .left(t12_add_left),
        .out(t12_add_out),
        .right(t12_add_right)
    );
    std_reg # (
        .width(5)
    ) t13_idx (
        .clk(t13_idx_clk),
        .done(t13_idx_done),
        .in(t13_idx_in),
        .out(t13_idx_out),
        .write_en(t13_idx_write_en)
    );
    std_add # (
        .width(5)
    ) t13_add (
        .left(t13_add_left),
        .out(t13_add_out),
        .right(t13_add_right)
    );
    std_reg # (
        .width(5)
    ) t14_idx (
        .clk(t14_idx_clk),
        .done(t14_idx_done),
        .in(t14_idx_in),
        .out(t14_idx_out),
        .write_en(t14_idx_write_en)
    );
    std_add # (
        .width(5)
    ) t14_add (
        .left(t14_add_left),
        .out(t14_add_out),
        .right(t14_add_right)
    );
    std_reg # (
        .width(5)
    ) t15_idx (
        .clk(t15_idx_clk),
        .done(t15_idx_done),
        .in(t15_idx_in),
        .out(t15_idx_out),
        .write_en(t15_idx_write_en)
    );
    std_add # (
        .width(5)
    ) t15_add (
        .left(t15_add_left),
        .out(t15_add_out),
        .right(t15_add_right)
    );
    std_reg # (
        .width(5)
    ) l0_idx (
        .clk(l0_idx_clk),
        .done(l0_idx_done),
        .in(l0_idx_in),
        .out(l0_idx_out),
        .write_en(l0_idx_write_en)
    );
    std_add # (
        .width(5)
    ) l0_add (
        .left(l0_add_left),
        .out(l0_add_out),
        .right(l0_add_right)
    );
    std_reg # (
        .width(5)
    ) l1_idx (
        .clk(l1_idx_clk),
        .done(l1_idx_done),
        .in(l1_idx_in),
        .out(l1_idx_out),
        .write_en(l1_idx_write_en)
    );
    std_add # (
        .width(5)
    ) l1_add (
        .left(l1_add_left),
        .out(l1_add_out),
        .right(l1_add_right)
    );
    std_reg # (
        .width(5)
    ) l2_idx (
        .clk(l2_idx_clk),
        .done(l2_idx_done),
        .in(l2_idx_in),
        .out(l2_idx_out),
        .write_en(l2_idx_write_en)
    );
    std_add # (
        .width(5)
    ) l2_add (
        .left(l2_add_left),
        .out(l2_add_out),
        .right(l2_add_right)
    );
    std_reg # (
        .width(5)
    ) l3_idx (
        .clk(l3_idx_clk),
        .done(l3_idx_done),
        .in(l3_idx_in),
        .out(l3_idx_out),
        .write_en(l3_idx_write_en)
    );
    std_add # (
        .width(5)
    ) l3_add (
        .left(l3_add_left),
        .out(l3_add_out),
        .right(l3_add_right)
    );
    std_reg # (
        .width(5)
    ) l4_idx (
        .clk(l4_idx_clk),
        .done(l4_idx_done),
        .in(l4_idx_in),
        .out(l4_idx_out),
        .write_en(l4_idx_write_en)
    );
    std_add # (
        .width(5)
    ) l4_add (
        .left(l4_add_left),
        .out(l4_add_out),
        .right(l4_add_right)
    );
    std_reg # (
        .width(5)
    ) l5_idx (
        .clk(l5_idx_clk),
        .done(l5_idx_done),
        .in(l5_idx_in),
        .out(l5_idx_out),
        .write_en(l5_idx_write_en)
    );
    std_add # (
        .width(5)
    ) l5_add (
        .left(l5_add_left),
        .out(l5_add_out),
        .right(l5_add_right)
    );
    std_reg # (
        .width(5)
    ) l6_idx (
        .clk(l6_idx_clk),
        .done(l6_idx_done),
        .in(l6_idx_in),
        .out(l6_idx_out),
        .write_en(l6_idx_write_en)
    );
    std_add # (
        .width(5)
    ) l6_add (
        .left(l6_add_left),
        .out(l6_add_out),
        .right(l6_add_right)
    );
    std_reg # (
        .width(5)
    ) l7_idx (
        .clk(l7_idx_clk),
        .done(l7_idx_done),
        .in(l7_idx_in),
        .out(l7_idx_out),
        .write_en(l7_idx_write_en)
    );
    std_add # (
        .width(5)
    ) l7_add (
        .left(l7_add_left),
        .out(l7_add_out),
        .right(l7_add_right)
    );
    std_reg # (
        .width(5)
    ) l8_idx (
        .clk(l8_idx_clk),
        .done(l8_idx_done),
        .in(l8_idx_in),
        .out(l8_idx_out),
        .write_en(l8_idx_write_en)
    );
    std_add # (
        .width(5)
    ) l8_add (
        .left(l8_add_left),
        .out(l8_add_out),
        .right(l8_add_right)
    );
    std_reg # (
        .width(5)
    ) l9_idx (
        .clk(l9_idx_clk),
        .done(l9_idx_done),
        .in(l9_idx_in),
        .out(l9_idx_out),
        .write_en(l9_idx_write_en)
    );
    std_add # (
        .width(5)
    ) l9_add (
        .left(l9_add_left),
        .out(l9_add_out),
        .right(l9_add_right)
    );
    std_reg # (
        .width(5)
    ) l10_idx (
        .clk(l10_idx_clk),
        .done(l10_idx_done),
        .in(l10_idx_in),
        .out(l10_idx_out),
        .write_en(l10_idx_write_en)
    );
    std_add # (
        .width(5)
    ) l10_add (
        .left(l10_add_left),
        .out(l10_add_out),
        .right(l10_add_right)
    );
    std_reg # (
        .width(5)
    ) l11_idx (
        .clk(l11_idx_clk),
        .done(l11_idx_done),
        .in(l11_idx_in),
        .out(l11_idx_out),
        .write_en(l11_idx_write_en)
    );
    std_add # (
        .width(5)
    ) l11_add (
        .left(l11_add_left),
        .out(l11_add_out),
        .right(l11_add_right)
    );
    std_reg # (
        .width(5)
    ) l12_idx (
        .clk(l12_idx_clk),
        .done(l12_idx_done),
        .in(l12_idx_in),
        .out(l12_idx_out),
        .write_en(l12_idx_write_en)
    );
    std_add # (
        .width(5)
    ) l12_add (
        .left(l12_add_left),
        .out(l12_add_out),
        .right(l12_add_right)
    );
    std_reg # (
        .width(5)
    ) l13_idx (
        .clk(l13_idx_clk),
        .done(l13_idx_done),
        .in(l13_idx_in),
        .out(l13_idx_out),
        .write_en(l13_idx_write_en)
    );
    std_add # (
        .width(5)
    ) l13_add (
        .left(l13_add_left),
        .out(l13_add_out),
        .right(l13_add_right)
    );
    std_reg # (
        .width(5)
    ) l14_idx (
        .clk(l14_idx_clk),
        .done(l14_idx_done),
        .in(l14_idx_in),
        .out(l14_idx_out),
        .write_en(l14_idx_write_en)
    );
    std_add # (
        .width(5)
    ) l14_add (
        .left(l14_add_left),
        .out(l14_add_out),
        .right(l14_add_right)
    );
    std_reg # (
        .width(5)
    ) l15_idx (
        .clk(l15_idx_clk),
        .done(l15_idx_done),
        .in(l15_idx_in),
        .out(l15_idx_out),
        .write_en(l15_idx_write_en)
    );
    std_add # (
        .width(5)
    ) l15_add (
        .left(l15_add_left),
        .out(l15_add_out),
        .right(l15_add_right)
    );
    mac_pe pe_0_0 (
        .clk(pe_0_0_clk),
        .done(pe_0_0_done),
        .go(pe_0_0_go),
        .left(pe_0_0_left),
        .out(pe_0_0_out),
        .top(pe_0_0_top)
    );
    std_reg # (
        .width(32)
    ) top_0_0 (
        .clk(top_0_0_clk),
        .done(top_0_0_done),
        .in(top_0_0_in),
        .out(top_0_0_out),
        .write_en(top_0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_0 (
        .clk(left_0_0_clk),
        .done(left_0_0_done),
        .in(left_0_0_in),
        .out(left_0_0_out),
        .write_en(left_0_0_write_en)
    );
    mac_pe pe_0_1 (
        .clk(pe_0_1_clk),
        .done(pe_0_1_done),
        .go(pe_0_1_go),
        .left(pe_0_1_left),
        .out(pe_0_1_out),
        .top(pe_0_1_top)
    );
    std_reg # (
        .width(32)
    ) top_0_1 (
        .clk(top_0_1_clk),
        .done(top_0_1_done),
        .in(top_0_1_in),
        .out(top_0_1_out),
        .write_en(top_0_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_1 (
        .clk(left_0_1_clk),
        .done(left_0_1_done),
        .in(left_0_1_in),
        .out(left_0_1_out),
        .write_en(left_0_1_write_en)
    );
    mac_pe pe_0_2 (
        .clk(pe_0_2_clk),
        .done(pe_0_2_done),
        .go(pe_0_2_go),
        .left(pe_0_2_left),
        .out(pe_0_2_out),
        .top(pe_0_2_top)
    );
    std_reg # (
        .width(32)
    ) top_0_2 (
        .clk(top_0_2_clk),
        .done(top_0_2_done),
        .in(top_0_2_in),
        .out(top_0_2_out),
        .write_en(top_0_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_2 (
        .clk(left_0_2_clk),
        .done(left_0_2_done),
        .in(left_0_2_in),
        .out(left_0_2_out),
        .write_en(left_0_2_write_en)
    );
    mac_pe pe_0_3 (
        .clk(pe_0_3_clk),
        .done(pe_0_3_done),
        .go(pe_0_3_go),
        .left(pe_0_3_left),
        .out(pe_0_3_out),
        .top(pe_0_3_top)
    );
    std_reg # (
        .width(32)
    ) top_0_3 (
        .clk(top_0_3_clk),
        .done(top_0_3_done),
        .in(top_0_3_in),
        .out(top_0_3_out),
        .write_en(top_0_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_3 (
        .clk(left_0_3_clk),
        .done(left_0_3_done),
        .in(left_0_3_in),
        .out(left_0_3_out),
        .write_en(left_0_3_write_en)
    );
    mac_pe pe_0_4 (
        .clk(pe_0_4_clk),
        .done(pe_0_4_done),
        .go(pe_0_4_go),
        .left(pe_0_4_left),
        .out(pe_0_4_out),
        .top(pe_0_4_top)
    );
    std_reg # (
        .width(32)
    ) top_0_4 (
        .clk(top_0_4_clk),
        .done(top_0_4_done),
        .in(top_0_4_in),
        .out(top_0_4_out),
        .write_en(top_0_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_4 (
        .clk(left_0_4_clk),
        .done(left_0_4_done),
        .in(left_0_4_in),
        .out(left_0_4_out),
        .write_en(left_0_4_write_en)
    );
    mac_pe pe_0_5 (
        .clk(pe_0_5_clk),
        .done(pe_0_5_done),
        .go(pe_0_5_go),
        .left(pe_0_5_left),
        .out(pe_0_5_out),
        .top(pe_0_5_top)
    );
    std_reg # (
        .width(32)
    ) top_0_5 (
        .clk(top_0_5_clk),
        .done(top_0_5_done),
        .in(top_0_5_in),
        .out(top_0_5_out),
        .write_en(top_0_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_5 (
        .clk(left_0_5_clk),
        .done(left_0_5_done),
        .in(left_0_5_in),
        .out(left_0_5_out),
        .write_en(left_0_5_write_en)
    );
    mac_pe pe_0_6 (
        .clk(pe_0_6_clk),
        .done(pe_0_6_done),
        .go(pe_0_6_go),
        .left(pe_0_6_left),
        .out(pe_0_6_out),
        .top(pe_0_6_top)
    );
    std_reg # (
        .width(32)
    ) top_0_6 (
        .clk(top_0_6_clk),
        .done(top_0_6_done),
        .in(top_0_6_in),
        .out(top_0_6_out),
        .write_en(top_0_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_6 (
        .clk(left_0_6_clk),
        .done(left_0_6_done),
        .in(left_0_6_in),
        .out(left_0_6_out),
        .write_en(left_0_6_write_en)
    );
    mac_pe pe_0_7 (
        .clk(pe_0_7_clk),
        .done(pe_0_7_done),
        .go(pe_0_7_go),
        .left(pe_0_7_left),
        .out(pe_0_7_out),
        .top(pe_0_7_top)
    );
    std_reg # (
        .width(32)
    ) top_0_7 (
        .clk(top_0_7_clk),
        .done(top_0_7_done),
        .in(top_0_7_in),
        .out(top_0_7_out),
        .write_en(top_0_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_7 (
        .clk(left_0_7_clk),
        .done(left_0_7_done),
        .in(left_0_7_in),
        .out(left_0_7_out),
        .write_en(left_0_7_write_en)
    );
    mac_pe pe_0_8 (
        .clk(pe_0_8_clk),
        .done(pe_0_8_done),
        .go(pe_0_8_go),
        .left(pe_0_8_left),
        .out(pe_0_8_out),
        .top(pe_0_8_top)
    );
    std_reg # (
        .width(32)
    ) top_0_8 (
        .clk(top_0_8_clk),
        .done(top_0_8_done),
        .in(top_0_8_in),
        .out(top_0_8_out),
        .write_en(top_0_8_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_8 (
        .clk(left_0_8_clk),
        .done(left_0_8_done),
        .in(left_0_8_in),
        .out(left_0_8_out),
        .write_en(left_0_8_write_en)
    );
    mac_pe pe_0_9 (
        .clk(pe_0_9_clk),
        .done(pe_0_9_done),
        .go(pe_0_9_go),
        .left(pe_0_9_left),
        .out(pe_0_9_out),
        .top(pe_0_9_top)
    );
    std_reg # (
        .width(32)
    ) top_0_9 (
        .clk(top_0_9_clk),
        .done(top_0_9_done),
        .in(top_0_9_in),
        .out(top_0_9_out),
        .write_en(top_0_9_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_9 (
        .clk(left_0_9_clk),
        .done(left_0_9_done),
        .in(left_0_9_in),
        .out(left_0_9_out),
        .write_en(left_0_9_write_en)
    );
    mac_pe pe_0_10 (
        .clk(pe_0_10_clk),
        .done(pe_0_10_done),
        .go(pe_0_10_go),
        .left(pe_0_10_left),
        .out(pe_0_10_out),
        .top(pe_0_10_top)
    );
    std_reg # (
        .width(32)
    ) top_0_10 (
        .clk(top_0_10_clk),
        .done(top_0_10_done),
        .in(top_0_10_in),
        .out(top_0_10_out),
        .write_en(top_0_10_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_10 (
        .clk(left_0_10_clk),
        .done(left_0_10_done),
        .in(left_0_10_in),
        .out(left_0_10_out),
        .write_en(left_0_10_write_en)
    );
    mac_pe pe_0_11 (
        .clk(pe_0_11_clk),
        .done(pe_0_11_done),
        .go(pe_0_11_go),
        .left(pe_0_11_left),
        .out(pe_0_11_out),
        .top(pe_0_11_top)
    );
    std_reg # (
        .width(32)
    ) top_0_11 (
        .clk(top_0_11_clk),
        .done(top_0_11_done),
        .in(top_0_11_in),
        .out(top_0_11_out),
        .write_en(top_0_11_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_11 (
        .clk(left_0_11_clk),
        .done(left_0_11_done),
        .in(left_0_11_in),
        .out(left_0_11_out),
        .write_en(left_0_11_write_en)
    );
    mac_pe pe_0_12 (
        .clk(pe_0_12_clk),
        .done(pe_0_12_done),
        .go(pe_0_12_go),
        .left(pe_0_12_left),
        .out(pe_0_12_out),
        .top(pe_0_12_top)
    );
    std_reg # (
        .width(32)
    ) top_0_12 (
        .clk(top_0_12_clk),
        .done(top_0_12_done),
        .in(top_0_12_in),
        .out(top_0_12_out),
        .write_en(top_0_12_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_12 (
        .clk(left_0_12_clk),
        .done(left_0_12_done),
        .in(left_0_12_in),
        .out(left_0_12_out),
        .write_en(left_0_12_write_en)
    );
    mac_pe pe_0_13 (
        .clk(pe_0_13_clk),
        .done(pe_0_13_done),
        .go(pe_0_13_go),
        .left(pe_0_13_left),
        .out(pe_0_13_out),
        .top(pe_0_13_top)
    );
    std_reg # (
        .width(32)
    ) top_0_13 (
        .clk(top_0_13_clk),
        .done(top_0_13_done),
        .in(top_0_13_in),
        .out(top_0_13_out),
        .write_en(top_0_13_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_13 (
        .clk(left_0_13_clk),
        .done(left_0_13_done),
        .in(left_0_13_in),
        .out(left_0_13_out),
        .write_en(left_0_13_write_en)
    );
    mac_pe pe_0_14 (
        .clk(pe_0_14_clk),
        .done(pe_0_14_done),
        .go(pe_0_14_go),
        .left(pe_0_14_left),
        .out(pe_0_14_out),
        .top(pe_0_14_top)
    );
    std_reg # (
        .width(32)
    ) top_0_14 (
        .clk(top_0_14_clk),
        .done(top_0_14_done),
        .in(top_0_14_in),
        .out(top_0_14_out),
        .write_en(top_0_14_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_14 (
        .clk(left_0_14_clk),
        .done(left_0_14_done),
        .in(left_0_14_in),
        .out(left_0_14_out),
        .write_en(left_0_14_write_en)
    );
    mac_pe pe_0_15 (
        .clk(pe_0_15_clk),
        .done(pe_0_15_done),
        .go(pe_0_15_go),
        .left(pe_0_15_left),
        .out(pe_0_15_out),
        .top(pe_0_15_top)
    );
    std_reg # (
        .width(32)
    ) top_0_15 (
        .clk(top_0_15_clk),
        .done(top_0_15_done),
        .in(top_0_15_in),
        .out(top_0_15_out),
        .write_en(top_0_15_write_en)
    );
    std_reg # (
        .width(32)
    ) left_0_15 (
        .clk(left_0_15_clk),
        .done(left_0_15_done),
        .in(left_0_15_in),
        .out(left_0_15_out),
        .write_en(left_0_15_write_en)
    );
    mac_pe pe_1_0 (
        .clk(pe_1_0_clk),
        .done(pe_1_0_done),
        .go(pe_1_0_go),
        .left(pe_1_0_left),
        .out(pe_1_0_out),
        .top(pe_1_0_top)
    );
    std_reg # (
        .width(32)
    ) top_1_0 (
        .clk(top_1_0_clk),
        .done(top_1_0_done),
        .in(top_1_0_in),
        .out(top_1_0_out),
        .write_en(top_1_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_0 (
        .clk(left_1_0_clk),
        .done(left_1_0_done),
        .in(left_1_0_in),
        .out(left_1_0_out),
        .write_en(left_1_0_write_en)
    );
    mac_pe pe_1_1 (
        .clk(pe_1_1_clk),
        .done(pe_1_1_done),
        .go(pe_1_1_go),
        .left(pe_1_1_left),
        .out(pe_1_1_out),
        .top(pe_1_1_top)
    );
    std_reg # (
        .width(32)
    ) top_1_1 (
        .clk(top_1_1_clk),
        .done(top_1_1_done),
        .in(top_1_1_in),
        .out(top_1_1_out),
        .write_en(top_1_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_1 (
        .clk(left_1_1_clk),
        .done(left_1_1_done),
        .in(left_1_1_in),
        .out(left_1_1_out),
        .write_en(left_1_1_write_en)
    );
    mac_pe pe_1_2 (
        .clk(pe_1_2_clk),
        .done(pe_1_2_done),
        .go(pe_1_2_go),
        .left(pe_1_2_left),
        .out(pe_1_2_out),
        .top(pe_1_2_top)
    );
    std_reg # (
        .width(32)
    ) top_1_2 (
        .clk(top_1_2_clk),
        .done(top_1_2_done),
        .in(top_1_2_in),
        .out(top_1_2_out),
        .write_en(top_1_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_2 (
        .clk(left_1_2_clk),
        .done(left_1_2_done),
        .in(left_1_2_in),
        .out(left_1_2_out),
        .write_en(left_1_2_write_en)
    );
    mac_pe pe_1_3 (
        .clk(pe_1_3_clk),
        .done(pe_1_3_done),
        .go(pe_1_3_go),
        .left(pe_1_3_left),
        .out(pe_1_3_out),
        .top(pe_1_3_top)
    );
    std_reg # (
        .width(32)
    ) top_1_3 (
        .clk(top_1_3_clk),
        .done(top_1_3_done),
        .in(top_1_3_in),
        .out(top_1_3_out),
        .write_en(top_1_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_3 (
        .clk(left_1_3_clk),
        .done(left_1_3_done),
        .in(left_1_3_in),
        .out(left_1_3_out),
        .write_en(left_1_3_write_en)
    );
    mac_pe pe_1_4 (
        .clk(pe_1_4_clk),
        .done(pe_1_4_done),
        .go(pe_1_4_go),
        .left(pe_1_4_left),
        .out(pe_1_4_out),
        .top(pe_1_4_top)
    );
    std_reg # (
        .width(32)
    ) top_1_4 (
        .clk(top_1_4_clk),
        .done(top_1_4_done),
        .in(top_1_4_in),
        .out(top_1_4_out),
        .write_en(top_1_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_4 (
        .clk(left_1_4_clk),
        .done(left_1_4_done),
        .in(left_1_4_in),
        .out(left_1_4_out),
        .write_en(left_1_4_write_en)
    );
    mac_pe pe_1_5 (
        .clk(pe_1_5_clk),
        .done(pe_1_5_done),
        .go(pe_1_5_go),
        .left(pe_1_5_left),
        .out(pe_1_5_out),
        .top(pe_1_5_top)
    );
    std_reg # (
        .width(32)
    ) top_1_5 (
        .clk(top_1_5_clk),
        .done(top_1_5_done),
        .in(top_1_5_in),
        .out(top_1_5_out),
        .write_en(top_1_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_5 (
        .clk(left_1_5_clk),
        .done(left_1_5_done),
        .in(left_1_5_in),
        .out(left_1_5_out),
        .write_en(left_1_5_write_en)
    );
    mac_pe pe_1_6 (
        .clk(pe_1_6_clk),
        .done(pe_1_6_done),
        .go(pe_1_6_go),
        .left(pe_1_6_left),
        .out(pe_1_6_out),
        .top(pe_1_6_top)
    );
    std_reg # (
        .width(32)
    ) top_1_6 (
        .clk(top_1_6_clk),
        .done(top_1_6_done),
        .in(top_1_6_in),
        .out(top_1_6_out),
        .write_en(top_1_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_6 (
        .clk(left_1_6_clk),
        .done(left_1_6_done),
        .in(left_1_6_in),
        .out(left_1_6_out),
        .write_en(left_1_6_write_en)
    );
    mac_pe pe_1_7 (
        .clk(pe_1_7_clk),
        .done(pe_1_7_done),
        .go(pe_1_7_go),
        .left(pe_1_7_left),
        .out(pe_1_7_out),
        .top(pe_1_7_top)
    );
    std_reg # (
        .width(32)
    ) top_1_7 (
        .clk(top_1_7_clk),
        .done(top_1_7_done),
        .in(top_1_7_in),
        .out(top_1_7_out),
        .write_en(top_1_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_7 (
        .clk(left_1_7_clk),
        .done(left_1_7_done),
        .in(left_1_7_in),
        .out(left_1_7_out),
        .write_en(left_1_7_write_en)
    );
    mac_pe pe_1_8 (
        .clk(pe_1_8_clk),
        .done(pe_1_8_done),
        .go(pe_1_8_go),
        .left(pe_1_8_left),
        .out(pe_1_8_out),
        .top(pe_1_8_top)
    );
    std_reg # (
        .width(32)
    ) top_1_8 (
        .clk(top_1_8_clk),
        .done(top_1_8_done),
        .in(top_1_8_in),
        .out(top_1_8_out),
        .write_en(top_1_8_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_8 (
        .clk(left_1_8_clk),
        .done(left_1_8_done),
        .in(left_1_8_in),
        .out(left_1_8_out),
        .write_en(left_1_8_write_en)
    );
    mac_pe pe_1_9 (
        .clk(pe_1_9_clk),
        .done(pe_1_9_done),
        .go(pe_1_9_go),
        .left(pe_1_9_left),
        .out(pe_1_9_out),
        .top(pe_1_9_top)
    );
    std_reg # (
        .width(32)
    ) top_1_9 (
        .clk(top_1_9_clk),
        .done(top_1_9_done),
        .in(top_1_9_in),
        .out(top_1_9_out),
        .write_en(top_1_9_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_9 (
        .clk(left_1_9_clk),
        .done(left_1_9_done),
        .in(left_1_9_in),
        .out(left_1_9_out),
        .write_en(left_1_9_write_en)
    );
    mac_pe pe_1_10 (
        .clk(pe_1_10_clk),
        .done(pe_1_10_done),
        .go(pe_1_10_go),
        .left(pe_1_10_left),
        .out(pe_1_10_out),
        .top(pe_1_10_top)
    );
    std_reg # (
        .width(32)
    ) top_1_10 (
        .clk(top_1_10_clk),
        .done(top_1_10_done),
        .in(top_1_10_in),
        .out(top_1_10_out),
        .write_en(top_1_10_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_10 (
        .clk(left_1_10_clk),
        .done(left_1_10_done),
        .in(left_1_10_in),
        .out(left_1_10_out),
        .write_en(left_1_10_write_en)
    );
    mac_pe pe_1_11 (
        .clk(pe_1_11_clk),
        .done(pe_1_11_done),
        .go(pe_1_11_go),
        .left(pe_1_11_left),
        .out(pe_1_11_out),
        .top(pe_1_11_top)
    );
    std_reg # (
        .width(32)
    ) top_1_11 (
        .clk(top_1_11_clk),
        .done(top_1_11_done),
        .in(top_1_11_in),
        .out(top_1_11_out),
        .write_en(top_1_11_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_11 (
        .clk(left_1_11_clk),
        .done(left_1_11_done),
        .in(left_1_11_in),
        .out(left_1_11_out),
        .write_en(left_1_11_write_en)
    );
    mac_pe pe_1_12 (
        .clk(pe_1_12_clk),
        .done(pe_1_12_done),
        .go(pe_1_12_go),
        .left(pe_1_12_left),
        .out(pe_1_12_out),
        .top(pe_1_12_top)
    );
    std_reg # (
        .width(32)
    ) top_1_12 (
        .clk(top_1_12_clk),
        .done(top_1_12_done),
        .in(top_1_12_in),
        .out(top_1_12_out),
        .write_en(top_1_12_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_12 (
        .clk(left_1_12_clk),
        .done(left_1_12_done),
        .in(left_1_12_in),
        .out(left_1_12_out),
        .write_en(left_1_12_write_en)
    );
    mac_pe pe_1_13 (
        .clk(pe_1_13_clk),
        .done(pe_1_13_done),
        .go(pe_1_13_go),
        .left(pe_1_13_left),
        .out(pe_1_13_out),
        .top(pe_1_13_top)
    );
    std_reg # (
        .width(32)
    ) top_1_13 (
        .clk(top_1_13_clk),
        .done(top_1_13_done),
        .in(top_1_13_in),
        .out(top_1_13_out),
        .write_en(top_1_13_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_13 (
        .clk(left_1_13_clk),
        .done(left_1_13_done),
        .in(left_1_13_in),
        .out(left_1_13_out),
        .write_en(left_1_13_write_en)
    );
    mac_pe pe_1_14 (
        .clk(pe_1_14_clk),
        .done(pe_1_14_done),
        .go(pe_1_14_go),
        .left(pe_1_14_left),
        .out(pe_1_14_out),
        .top(pe_1_14_top)
    );
    std_reg # (
        .width(32)
    ) top_1_14 (
        .clk(top_1_14_clk),
        .done(top_1_14_done),
        .in(top_1_14_in),
        .out(top_1_14_out),
        .write_en(top_1_14_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_14 (
        .clk(left_1_14_clk),
        .done(left_1_14_done),
        .in(left_1_14_in),
        .out(left_1_14_out),
        .write_en(left_1_14_write_en)
    );
    mac_pe pe_1_15 (
        .clk(pe_1_15_clk),
        .done(pe_1_15_done),
        .go(pe_1_15_go),
        .left(pe_1_15_left),
        .out(pe_1_15_out),
        .top(pe_1_15_top)
    );
    std_reg # (
        .width(32)
    ) top_1_15 (
        .clk(top_1_15_clk),
        .done(top_1_15_done),
        .in(top_1_15_in),
        .out(top_1_15_out),
        .write_en(top_1_15_write_en)
    );
    std_reg # (
        .width(32)
    ) left_1_15 (
        .clk(left_1_15_clk),
        .done(left_1_15_done),
        .in(left_1_15_in),
        .out(left_1_15_out),
        .write_en(left_1_15_write_en)
    );
    mac_pe pe_2_0 (
        .clk(pe_2_0_clk),
        .done(pe_2_0_done),
        .go(pe_2_0_go),
        .left(pe_2_0_left),
        .out(pe_2_0_out),
        .top(pe_2_0_top)
    );
    std_reg # (
        .width(32)
    ) top_2_0 (
        .clk(top_2_0_clk),
        .done(top_2_0_done),
        .in(top_2_0_in),
        .out(top_2_0_out),
        .write_en(top_2_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_0 (
        .clk(left_2_0_clk),
        .done(left_2_0_done),
        .in(left_2_0_in),
        .out(left_2_0_out),
        .write_en(left_2_0_write_en)
    );
    mac_pe pe_2_1 (
        .clk(pe_2_1_clk),
        .done(pe_2_1_done),
        .go(pe_2_1_go),
        .left(pe_2_1_left),
        .out(pe_2_1_out),
        .top(pe_2_1_top)
    );
    std_reg # (
        .width(32)
    ) top_2_1 (
        .clk(top_2_1_clk),
        .done(top_2_1_done),
        .in(top_2_1_in),
        .out(top_2_1_out),
        .write_en(top_2_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_1 (
        .clk(left_2_1_clk),
        .done(left_2_1_done),
        .in(left_2_1_in),
        .out(left_2_1_out),
        .write_en(left_2_1_write_en)
    );
    mac_pe pe_2_2 (
        .clk(pe_2_2_clk),
        .done(pe_2_2_done),
        .go(pe_2_2_go),
        .left(pe_2_2_left),
        .out(pe_2_2_out),
        .top(pe_2_2_top)
    );
    std_reg # (
        .width(32)
    ) top_2_2 (
        .clk(top_2_2_clk),
        .done(top_2_2_done),
        .in(top_2_2_in),
        .out(top_2_2_out),
        .write_en(top_2_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_2 (
        .clk(left_2_2_clk),
        .done(left_2_2_done),
        .in(left_2_2_in),
        .out(left_2_2_out),
        .write_en(left_2_2_write_en)
    );
    mac_pe pe_2_3 (
        .clk(pe_2_3_clk),
        .done(pe_2_3_done),
        .go(pe_2_3_go),
        .left(pe_2_3_left),
        .out(pe_2_3_out),
        .top(pe_2_3_top)
    );
    std_reg # (
        .width(32)
    ) top_2_3 (
        .clk(top_2_3_clk),
        .done(top_2_3_done),
        .in(top_2_3_in),
        .out(top_2_3_out),
        .write_en(top_2_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_3 (
        .clk(left_2_3_clk),
        .done(left_2_3_done),
        .in(left_2_3_in),
        .out(left_2_3_out),
        .write_en(left_2_3_write_en)
    );
    mac_pe pe_2_4 (
        .clk(pe_2_4_clk),
        .done(pe_2_4_done),
        .go(pe_2_4_go),
        .left(pe_2_4_left),
        .out(pe_2_4_out),
        .top(pe_2_4_top)
    );
    std_reg # (
        .width(32)
    ) top_2_4 (
        .clk(top_2_4_clk),
        .done(top_2_4_done),
        .in(top_2_4_in),
        .out(top_2_4_out),
        .write_en(top_2_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_4 (
        .clk(left_2_4_clk),
        .done(left_2_4_done),
        .in(left_2_4_in),
        .out(left_2_4_out),
        .write_en(left_2_4_write_en)
    );
    mac_pe pe_2_5 (
        .clk(pe_2_5_clk),
        .done(pe_2_5_done),
        .go(pe_2_5_go),
        .left(pe_2_5_left),
        .out(pe_2_5_out),
        .top(pe_2_5_top)
    );
    std_reg # (
        .width(32)
    ) top_2_5 (
        .clk(top_2_5_clk),
        .done(top_2_5_done),
        .in(top_2_5_in),
        .out(top_2_5_out),
        .write_en(top_2_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_5 (
        .clk(left_2_5_clk),
        .done(left_2_5_done),
        .in(left_2_5_in),
        .out(left_2_5_out),
        .write_en(left_2_5_write_en)
    );
    mac_pe pe_2_6 (
        .clk(pe_2_6_clk),
        .done(pe_2_6_done),
        .go(pe_2_6_go),
        .left(pe_2_6_left),
        .out(pe_2_6_out),
        .top(pe_2_6_top)
    );
    std_reg # (
        .width(32)
    ) top_2_6 (
        .clk(top_2_6_clk),
        .done(top_2_6_done),
        .in(top_2_6_in),
        .out(top_2_6_out),
        .write_en(top_2_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_6 (
        .clk(left_2_6_clk),
        .done(left_2_6_done),
        .in(left_2_6_in),
        .out(left_2_6_out),
        .write_en(left_2_6_write_en)
    );
    mac_pe pe_2_7 (
        .clk(pe_2_7_clk),
        .done(pe_2_7_done),
        .go(pe_2_7_go),
        .left(pe_2_7_left),
        .out(pe_2_7_out),
        .top(pe_2_7_top)
    );
    std_reg # (
        .width(32)
    ) top_2_7 (
        .clk(top_2_7_clk),
        .done(top_2_7_done),
        .in(top_2_7_in),
        .out(top_2_7_out),
        .write_en(top_2_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_7 (
        .clk(left_2_7_clk),
        .done(left_2_7_done),
        .in(left_2_7_in),
        .out(left_2_7_out),
        .write_en(left_2_7_write_en)
    );
    mac_pe pe_2_8 (
        .clk(pe_2_8_clk),
        .done(pe_2_8_done),
        .go(pe_2_8_go),
        .left(pe_2_8_left),
        .out(pe_2_8_out),
        .top(pe_2_8_top)
    );
    std_reg # (
        .width(32)
    ) top_2_8 (
        .clk(top_2_8_clk),
        .done(top_2_8_done),
        .in(top_2_8_in),
        .out(top_2_8_out),
        .write_en(top_2_8_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_8 (
        .clk(left_2_8_clk),
        .done(left_2_8_done),
        .in(left_2_8_in),
        .out(left_2_8_out),
        .write_en(left_2_8_write_en)
    );
    mac_pe pe_2_9 (
        .clk(pe_2_9_clk),
        .done(pe_2_9_done),
        .go(pe_2_9_go),
        .left(pe_2_9_left),
        .out(pe_2_9_out),
        .top(pe_2_9_top)
    );
    std_reg # (
        .width(32)
    ) top_2_9 (
        .clk(top_2_9_clk),
        .done(top_2_9_done),
        .in(top_2_9_in),
        .out(top_2_9_out),
        .write_en(top_2_9_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_9 (
        .clk(left_2_9_clk),
        .done(left_2_9_done),
        .in(left_2_9_in),
        .out(left_2_9_out),
        .write_en(left_2_9_write_en)
    );
    mac_pe pe_2_10 (
        .clk(pe_2_10_clk),
        .done(pe_2_10_done),
        .go(pe_2_10_go),
        .left(pe_2_10_left),
        .out(pe_2_10_out),
        .top(pe_2_10_top)
    );
    std_reg # (
        .width(32)
    ) top_2_10 (
        .clk(top_2_10_clk),
        .done(top_2_10_done),
        .in(top_2_10_in),
        .out(top_2_10_out),
        .write_en(top_2_10_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_10 (
        .clk(left_2_10_clk),
        .done(left_2_10_done),
        .in(left_2_10_in),
        .out(left_2_10_out),
        .write_en(left_2_10_write_en)
    );
    mac_pe pe_2_11 (
        .clk(pe_2_11_clk),
        .done(pe_2_11_done),
        .go(pe_2_11_go),
        .left(pe_2_11_left),
        .out(pe_2_11_out),
        .top(pe_2_11_top)
    );
    std_reg # (
        .width(32)
    ) top_2_11 (
        .clk(top_2_11_clk),
        .done(top_2_11_done),
        .in(top_2_11_in),
        .out(top_2_11_out),
        .write_en(top_2_11_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_11 (
        .clk(left_2_11_clk),
        .done(left_2_11_done),
        .in(left_2_11_in),
        .out(left_2_11_out),
        .write_en(left_2_11_write_en)
    );
    mac_pe pe_2_12 (
        .clk(pe_2_12_clk),
        .done(pe_2_12_done),
        .go(pe_2_12_go),
        .left(pe_2_12_left),
        .out(pe_2_12_out),
        .top(pe_2_12_top)
    );
    std_reg # (
        .width(32)
    ) top_2_12 (
        .clk(top_2_12_clk),
        .done(top_2_12_done),
        .in(top_2_12_in),
        .out(top_2_12_out),
        .write_en(top_2_12_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_12 (
        .clk(left_2_12_clk),
        .done(left_2_12_done),
        .in(left_2_12_in),
        .out(left_2_12_out),
        .write_en(left_2_12_write_en)
    );
    mac_pe pe_2_13 (
        .clk(pe_2_13_clk),
        .done(pe_2_13_done),
        .go(pe_2_13_go),
        .left(pe_2_13_left),
        .out(pe_2_13_out),
        .top(pe_2_13_top)
    );
    std_reg # (
        .width(32)
    ) top_2_13 (
        .clk(top_2_13_clk),
        .done(top_2_13_done),
        .in(top_2_13_in),
        .out(top_2_13_out),
        .write_en(top_2_13_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_13 (
        .clk(left_2_13_clk),
        .done(left_2_13_done),
        .in(left_2_13_in),
        .out(left_2_13_out),
        .write_en(left_2_13_write_en)
    );
    mac_pe pe_2_14 (
        .clk(pe_2_14_clk),
        .done(pe_2_14_done),
        .go(pe_2_14_go),
        .left(pe_2_14_left),
        .out(pe_2_14_out),
        .top(pe_2_14_top)
    );
    std_reg # (
        .width(32)
    ) top_2_14 (
        .clk(top_2_14_clk),
        .done(top_2_14_done),
        .in(top_2_14_in),
        .out(top_2_14_out),
        .write_en(top_2_14_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_14 (
        .clk(left_2_14_clk),
        .done(left_2_14_done),
        .in(left_2_14_in),
        .out(left_2_14_out),
        .write_en(left_2_14_write_en)
    );
    mac_pe pe_2_15 (
        .clk(pe_2_15_clk),
        .done(pe_2_15_done),
        .go(pe_2_15_go),
        .left(pe_2_15_left),
        .out(pe_2_15_out),
        .top(pe_2_15_top)
    );
    std_reg # (
        .width(32)
    ) top_2_15 (
        .clk(top_2_15_clk),
        .done(top_2_15_done),
        .in(top_2_15_in),
        .out(top_2_15_out),
        .write_en(top_2_15_write_en)
    );
    std_reg # (
        .width(32)
    ) left_2_15 (
        .clk(left_2_15_clk),
        .done(left_2_15_done),
        .in(left_2_15_in),
        .out(left_2_15_out),
        .write_en(left_2_15_write_en)
    );
    mac_pe pe_3_0 (
        .clk(pe_3_0_clk),
        .done(pe_3_0_done),
        .go(pe_3_0_go),
        .left(pe_3_0_left),
        .out(pe_3_0_out),
        .top(pe_3_0_top)
    );
    std_reg # (
        .width(32)
    ) top_3_0 (
        .clk(top_3_0_clk),
        .done(top_3_0_done),
        .in(top_3_0_in),
        .out(top_3_0_out),
        .write_en(top_3_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_0 (
        .clk(left_3_0_clk),
        .done(left_3_0_done),
        .in(left_3_0_in),
        .out(left_3_0_out),
        .write_en(left_3_0_write_en)
    );
    mac_pe pe_3_1 (
        .clk(pe_3_1_clk),
        .done(pe_3_1_done),
        .go(pe_3_1_go),
        .left(pe_3_1_left),
        .out(pe_3_1_out),
        .top(pe_3_1_top)
    );
    std_reg # (
        .width(32)
    ) top_3_1 (
        .clk(top_3_1_clk),
        .done(top_3_1_done),
        .in(top_3_1_in),
        .out(top_3_1_out),
        .write_en(top_3_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_1 (
        .clk(left_3_1_clk),
        .done(left_3_1_done),
        .in(left_3_1_in),
        .out(left_3_1_out),
        .write_en(left_3_1_write_en)
    );
    mac_pe pe_3_2 (
        .clk(pe_3_2_clk),
        .done(pe_3_2_done),
        .go(pe_3_2_go),
        .left(pe_3_2_left),
        .out(pe_3_2_out),
        .top(pe_3_2_top)
    );
    std_reg # (
        .width(32)
    ) top_3_2 (
        .clk(top_3_2_clk),
        .done(top_3_2_done),
        .in(top_3_2_in),
        .out(top_3_2_out),
        .write_en(top_3_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_2 (
        .clk(left_3_2_clk),
        .done(left_3_2_done),
        .in(left_3_2_in),
        .out(left_3_2_out),
        .write_en(left_3_2_write_en)
    );
    mac_pe pe_3_3 (
        .clk(pe_3_3_clk),
        .done(pe_3_3_done),
        .go(pe_3_3_go),
        .left(pe_3_3_left),
        .out(pe_3_3_out),
        .top(pe_3_3_top)
    );
    std_reg # (
        .width(32)
    ) top_3_3 (
        .clk(top_3_3_clk),
        .done(top_3_3_done),
        .in(top_3_3_in),
        .out(top_3_3_out),
        .write_en(top_3_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_3 (
        .clk(left_3_3_clk),
        .done(left_3_3_done),
        .in(left_3_3_in),
        .out(left_3_3_out),
        .write_en(left_3_3_write_en)
    );
    mac_pe pe_3_4 (
        .clk(pe_3_4_clk),
        .done(pe_3_4_done),
        .go(pe_3_4_go),
        .left(pe_3_4_left),
        .out(pe_3_4_out),
        .top(pe_3_4_top)
    );
    std_reg # (
        .width(32)
    ) top_3_4 (
        .clk(top_3_4_clk),
        .done(top_3_4_done),
        .in(top_3_4_in),
        .out(top_3_4_out),
        .write_en(top_3_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_4 (
        .clk(left_3_4_clk),
        .done(left_3_4_done),
        .in(left_3_4_in),
        .out(left_3_4_out),
        .write_en(left_3_4_write_en)
    );
    mac_pe pe_3_5 (
        .clk(pe_3_5_clk),
        .done(pe_3_5_done),
        .go(pe_3_5_go),
        .left(pe_3_5_left),
        .out(pe_3_5_out),
        .top(pe_3_5_top)
    );
    std_reg # (
        .width(32)
    ) top_3_5 (
        .clk(top_3_5_clk),
        .done(top_3_5_done),
        .in(top_3_5_in),
        .out(top_3_5_out),
        .write_en(top_3_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_5 (
        .clk(left_3_5_clk),
        .done(left_3_5_done),
        .in(left_3_5_in),
        .out(left_3_5_out),
        .write_en(left_3_5_write_en)
    );
    mac_pe pe_3_6 (
        .clk(pe_3_6_clk),
        .done(pe_3_6_done),
        .go(pe_3_6_go),
        .left(pe_3_6_left),
        .out(pe_3_6_out),
        .top(pe_3_6_top)
    );
    std_reg # (
        .width(32)
    ) top_3_6 (
        .clk(top_3_6_clk),
        .done(top_3_6_done),
        .in(top_3_6_in),
        .out(top_3_6_out),
        .write_en(top_3_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_6 (
        .clk(left_3_6_clk),
        .done(left_3_6_done),
        .in(left_3_6_in),
        .out(left_3_6_out),
        .write_en(left_3_6_write_en)
    );
    mac_pe pe_3_7 (
        .clk(pe_3_7_clk),
        .done(pe_3_7_done),
        .go(pe_3_7_go),
        .left(pe_3_7_left),
        .out(pe_3_7_out),
        .top(pe_3_7_top)
    );
    std_reg # (
        .width(32)
    ) top_3_7 (
        .clk(top_3_7_clk),
        .done(top_3_7_done),
        .in(top_3_7_in),
        .out(top_3_7_out),
        .write_en(top_3_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_7 (
        .clk(left_3_7_clk),
        .done(left_3_7_done),
        .in(left_3_7_in),
        .out(left_3_7_out),
        .write_en(left_3_7_write_en)
    );
    mac_pe pe_3_8 (
        .clk(pe_3_8_clk),
        .done(pe_3_8_done),
        .go(pe_3_8_go),
        .left(pe_3_8_left),
        .out(pe_3_8_out),
        .top(pe_3_8_top)
    );
    std_reg # (
        .width(32)
    ) top_3_8 (
        .clk(top_3_8_clk),
        .done(top_3_8_done),
        .in(top_3_8_in),
        .out(top_3_8_out),
        .write_en(top_3_8_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_8 (
        .clk(left_3_8_clk),
        .done(left_3_8_done),
        .in(left_3_8_in),
        .out(left_3_8_out),
        .write_en(left_3_8_write_en)
    );
    mac_pe pe_3_9 (
        .clk(pe_3_9_clk),
        .done(pe_3_9_done),
        .go(pe_3_9_go),
        .left(pe_3_9_left),
        .out(pe_3_9_out),
        .top(pe_3_9_top)
    );
    std_reg # (
        .width(32)
    ) top_3_9 (
        .clk(top_3_9_clk),
        .done(top_3_9_done),
        .in(top_3_9_in),
        .out(top_3_9_out),
        .write_en(top_3_9_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_9 (
        .clk(left_3_9_clk),
        .done(left_3_9_done),
        .in(left_3_9_in),
        .out(left_3_9_out),
        .write_en(left_3_9_write_en)
    );
    mac_pe pe_3_10 (
        .clk(pe_3_10_clk),
        .done(pe_3_10_done),
        .go(pe_3_10_go),
        .left(pe_3_10_left),
        .out(pe_3_10_out),
        .top(pe_3_10_top)
    );
    std_reg # (
        .width(32)
    ) top_3_10 (
        .clk(top_3_10_clk),
        .done(top_3_10_done),
        .in(top_3_10_in),
        .out(top_3_10_out),
        .write_en(top_3_10_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_10 (
        .clk(left_3_10_clk),
        .done(left_3_10_done),
        .in(left_3_10_in),
        .out(left_3_10_out),
        .write_en(left_3_10_write_en)
    );
    mac_pe pe_3_11 (
        .clk(pe_3_11_clk),
        .done(pe_3_11_done),
        .go(pe_3_11_go),
        .left(pe_3_11_left),
        .out(pe_3_11_out),
        .top(pe_3_11_top)
    );
    std_reg # (
        .width(32)
    ) top_3_11 (
        .clk(top_3_11_clk),
        .done(top_3_11_done),
        .in(top_3_11_in),
        .out(top_3_11_out),
        .write_en(top_3_11_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_11 (
        .clk(left_3_11_clk),
        .done(left_3_11_done),
        .in(left_3_11_in),
        .out(left_3_11_out),
        .write_en(left_3_11_write_en)
    );
    mac_pe pe_3_12 (
        .clk(pe_3_12_clk),
        .done(pe_3_12_done),
        .go(pe_3_12_go),
        .left(pe_3_12_left),
        .out(pe_3_12_out),
        .top(pe_3_12_top)
    );
    std_reg # (
        .width(32)
    ) top_3_12 (
        .clk(top_3_12_clk),
        .done(top_3_12_done),
        .in(top_3_12_in),
        .out(top_3_12_out),
        .write_en(top_3_12_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_12 (
        .clk(left_3_12_clk),
        .done(left_3_12_done),
        .in(left_3_12_in),
        .out(left_3_12_out),
        .write_en(left_3_12_write_en)
    );
    mac_pe pe_3_13 (
        .clk(pe_3_13_clk),
        .done(pe_3_13_done),
        .go(pe_3_13_go),
        .left(pe_3_13_left),
        .out(pe_3_13_out),
        .top(pe_3_13_top)
    );
    std_reg # (
        .width(32)
    ) top_3_13 (
        .clk(top_3_13_clk),
        .done(top_3_13_done),
        .in(top_3_13_in),
        .out(top_3_13_out),
        .write_en(top_3_13_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_13 (
        .clk(left_3_13_clk),
        .done(left_3_13_done),
        .in(left_3_13_in),
        .out(left_3_13_out),
        .write_en(left_3_13_write_en)
    );
    mac_pe pe_3_14 (
        .clk(pe_3_14_clk),
        .done(pe_3_14_done),
        .go(pe_3_14_go),
        .left(pe_3_14_left),
        .out(pe_3_14_out),
        .top(pe_3_14_top)
    );
    std_reg # (
        .width(32)
    ) top_3_14 (
        .clk(top_3_14_clk),
        .done(top_3_14_done),
        .in(top_3_14_in),
        .out(top_3_14_out),
        .write_en(top_3_14_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_14 (
        .clk(left_3_14_clk),
        .done(left_3_14_done),
        .in(left_3_14_in),
        .out(left_3_14_out),
        .write_en(left_3_14_write_en)
    );
    mac_pe pe_3_15 (
        .clk(pe_3_15_clk),
        .done(pe_3_15_done),
        .go(pe_3_15_go),
        .left(pe_3_15_left),
        .out(pe_3_15_out),
        .top(pe_3_15_top)
    );
    std_reg # (
        .width(32)
    ) top_3_15 (
        .clk(top_3_15_clk),
        .done(top_3_15_done),
        .in(top_3_15_in),
        .out(top_3_15_out),
        .write_en(top_3_15_write_en)
    );
    std_reg # (
        .width(32)
    ) left_3_15 (
        .clk(left_3_15_clk),
        .done(left_3_15_done),
        .in(left_3_15_in),
        .out(left_3_15_out),
        .write_en(left_3_15_write_en)
    );
    mac_pe pe_4_0 (
        .clk(pe_4_0_clk),
        .done(pe_4_0_done),
        .go(pe_4_0_go),
        .left(pe_4_0_left),
        .out(pe_4_0_out),
        .top(pe_4_0_top)
    );
    std_reg # (
        .width(32)
    ) top_4_0 (
        .clk(top_4_0_clk),
        .done(top_4_0_done),
        .in(top_4_0_in),
        .out(top_4_0_out),
        .write_en(top_4_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_0 (
        .clk(left_4_0_clk),
        .done(left_4_0_done),
        .in(left_4_0_in),
        .out(left_4_0_out),
        .write_en(left_4_0_write_en)
    );
    mac_pe pe_4_1 (
        .clk(pe_4_1_clk),
        .done(pe_4_1_done),
        .go(pe_4_1_go),
        .left(pe_4_1_left),
        .out(pe_4_1_out),
        .top(pe_4_1_top)
    );
    std_reg # (
        .width(32)
    ) top_4_1 (
        .clk(top_4_1_clk),
        .done(top_4_1_done),
        .in(top_4_1_in),
        .out(top_4_1_out),
        .write_en(top_4_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_1 (
        .clk(left_4_1_clk),
        .done(left_4_1_done),
        .in(left_4_1_in),
        .out(left_4_1_out),
        .write_en(left_4_1_write_en)
    );
    mac_pe pe_4_2 (
        .clk(pe_4_2_clk),
        .done(pe_4_2_done),
        .go(pe_4_2_go),
        .left(pe_4_2_left),
        .out(pe_4_2_out),
        .top(pe_4_2_top)
    );
    std_reg # (
        .width(32)
    ) top_4_2 (
        .clk(top_4_2_clk),
        .done(top_4_2_done),
        .in(top_4_2_in),
        .out(top_4_2_out),
        .write_en(top_4_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_2 (
        .clk(left_4_2_clk),
        .done(left_4_2_done),
        .in(left_4_2_in),
        .out(left_4_2_out),
        .write_en(left_4_2_write_en)
    );
    mac_pe pe_4_3 (
        .clk(pe_4_3_clk),
        .done(pe_4_3_done),
        .go(pe_4_3_go),
        .left(pe_4_3_left),
        .out(pe_4_3_out),
        .top(pe_4_3_top)
    );
    std_reg # (
        .width(32)
    ) top_4_3 (
        .clk(top_4_3_clk),
        .done(top_4_3_done),
        .in(top_4_3_in),
        .out(top_4_3_out),
        .write_en(top_4_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_3 (
        .clk(left_4_3_clk),
        .done(left_4_3_done),
        .in(left_4_3_in),
        .out(left_4_3_out),
        .write_en(left_4_3_write_en)
    );
    mac_pe pe_4_4 (
        .clk(pe_4_4_clk),
        .done(pe_4_4_done),
        .go(pe_4_4_go),
        .left(pe_4_4_left),
        .out(pe_4_4_out),
        .top(pe_4_4_top)
    );
    std_reg # (
        .width(32)
    ) top_4_4 (
        .clk(top_4_4_clk),
        .done(top_4_4_done),
        .in(top_4_4_in),
        .out(top_4_4_out),
        .write_en(top_4_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_4 (
        .clk(left_4_4_clk),
        .done(left_4_4_done),
        .in(left_4_4_in),
        .out(left_4_4_out),
        .write_en(left_4_4_write_en)
    );
    mac_pe pe_4_5 (
        .clk(pe_4_5_clk),
        .done(pe_4_5_done),
        .go(pe_4_5_go),
        .left(pe_4_5_left),
        .out(pe_4_5_out),
        .top(pe_4_5_top)
    );
    std_reg # (
        .width(32)
    ) top_4_5 (
        .clk(top_4_5_clk),
        .done(top_4_5_done),
        .in(top_4_5_in),
        .out(top_4_5_out),
        .write_en(top_4_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_5 (
        .clk(left_4_5_clk),
        .done(left_4_5_done),
        .in(left_4_5_in),
        .out(left_4_5_out),
        .write_en(left_4_5_write_en)
    );
    mac_pe pe_4_6 (
        .clk(pe_4_6_clk),
        .done(pe_4_6_done),
        .go(pe_4_6_go),
        .left(pe_4_6_left),
        .out(pe_4_6_out),
        .top(pe_4_6_top)
    );
    std_reg # (
        .width(32)
    ) top_4_6 (
        .clk(top_4_6_clk),
        .done(top_4_6_done),
        .in(top_4_6_in),
        .out(top_4_6_out),
        .write_en(top_4_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_6 (
        .clk(left_4_6_clk),
        .done(left_4_6_done),
        .in(left_4_6_in),
        .out(left_4_6_out),
        .write_en(left_4_6_write_en)
    );
    mac_pe pe_4_7 (
        .clk(pe_4_7_clk),
        .done(pe_4_7_done),
        .go(pe_4_7_go),
        .left(pe_4_7_left),
        .out(pe_4_7_out),
        .top(pe_4_7_top)
    );
    std_reg # (
        .width(32)
    ) top_4_7 (
        .clk(top_4_7_clk),
        .done(top_4_7_done),
        .in(top_4_7_in),
        .out(top_4_7_out),
        .write_en(top_4_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_7 (
        .clk(left_4_7_clk),
        .done(left_4_7_done),
        .in(left_4_7_in),
        .out(left_4_7_out),
        .write_en(left_4_7_write_en)
    );
    mac_pe pe_4_8 (
        .clk(pe_4_8_clk),
        .done(pe_4_8_done),
        .go(pe_4_8_go),
        .left(pe_4_8_left),
        .out(pe_4_8_out),
        .top(pe_4_8_top)
    );
    std_reg # (
        .width(32)
    ) top_4_8 (
        .clk(top_4_8_clk),
        .done(top_4_8_done),
        .in(top_4_8_in),
        .out(top_4_8_out),
        .write_en(top_4_8_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_8 (
        .clk(left_4_8_clk),
        .done(left_4_8_done),
        .in(left_4_8_in),
        .out(left_4_8_out),
        .write_en(left_4_8_write_en)
    );
    mac_pe pe_4_9 (
        .clk(pe_4_9_clk),
        .done(pe_4_9_done),
        .go(pe_4_9_go),
        .left(pe_4_9_left),
        .out(pe_4_9_out),
        .top(pe_4_9_top)
    );
    std_reg # (
        .width(32)
    ) top_4_9 (
        .clk(top_4_9_clk),
        .done(top_4_9_done),
        .in(top_4_9_in),
        .out(top_4_9_out),
        .write_en(top_4_9_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_9 (
        .clk(left_4_9_clk),
        .done(left_4_9_done),
        .in(left_4_9_in),
        .out(left_4_9_out),
        .write_en(left_4_9_write_en)
    );
    mac_pe pe_4_10 (
        .clk(pe_4_10_clk),
        .done(pe_4_10_done),
        .go(pe_4_10_go),
        .left(pe_4_10_left),
        .out(pe_4_10_out),
        .top(pe_4_10_top)
    );
    std_reg # (
        .width(32)
    ) top_4_10 (
        .clk(top_4_10_clk),
        .done(top_4_10_done),
        .in(top_4_10_in),
        .out(top_4_10_out),
        .write_en(top_4_10_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_10 (
        .clk(left_4_10_clk),
        .done(left_4_10_done),
        .in(left_4_10_in),
        .out(left_4_10_out),
        .write_en(left_4_10_write_en)
    );
    mac_pe pe_4_11 (
        .clk(pe_4_11_clk),
        .done(pe_4_11_done),
        .go(pe_4_11_go),
        .left(pe_4_11_left),
        .out(pe_4_11_out),
        .top(pe_4_11_top)
    );
    std_reg # (
        .width(32)
    ) top_4_11 (
        .clk(top_4_11_clk),
        .done(top_4_11_done),
        .in(top_4_11_in),
        .out(top_4_11_out),
        .write_en(top_4_11_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_11 (
        .clk(left_4_11_clk),
        .done(left_4_11_done),
        .in(left_4_11_in),
        .out(left_4_11_out),
        .write_en(left_4_11_write_en)
    );
    mac_pe pe_4_12 (
        .clk(pe_4_12_clk),
        .done(pe_4_12_done),
        .go(pe_4_12_go),
        .left(pe_4_12_left),
        .out(pe_4_12_out),
        .top(pe_4_12_top)
    );
    std_reg # (
        .width(32)
    ) top_4_12 (
        .clk(top_4_12_clk),
        .done(top_4_12_done),
        .in(top_4_12_in),
        .out(top_4_12_out),
        .write_en(top_4_12_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_12 (
        .clk(left_4_12_clk),
        .done(left_4_12_done),
        .in(left_4_12_in),
        .out(left_4_12_out),
        .write_en(left_4_12_write_en)
    );
    mac_pe pe_4_13 (
        .clk(pe_4_13_clk),
        .done(pe_4_13_done),
        .go(pe_4_13_go),
        .left(pe_4_13_left),
        .out(pe_4_13_out),
        .top(pe_4_13_top)
    );
    std_reg # (
        .width(32)
    ) top_4_13 (
        .clk(top_4_13_clk),
        .done(top_4_13_done),
        .in(top_4_13_in),
        .out(top_4_13_out),
        .write_en(top_4_13_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_13 (
        .clk(left_4_13_clk),
        .done(left_4_13_done),
        .in(left_4_13_in),
        .out(left_4_13_out),
        .write_en(left_4_13_write_en)
    );
    mac_pe pe_4_14 (
        .clk(pe_4_14_clk),
        .done(pe_4_14_done),
        .go(pe_4_14_go),
        .left(pe_4_14_left),
        .out(pe_4_14_out),
        .top(pe_4_14_top)
    );
    std_reg # (
        .width(32)
    ) top_4_14 (
        .clk(top_4_14_clk),
        .done(top_4_14_done),
        .in(top_4_14_in),
        .out(top_4_14_out),
        .write_en(top_4_14_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_14 (
        .clk(left_4_14_clk),
        .done(left_4_14_done),
        .in(left_4_14_in),
        .out(left_4_14_out),
        .write_en(left_4_14_write_en)
    );
    mac_pe pe_4_15 (
        .clk(pe_4_15_clk),
        .done(pe_4_15_done),
        .go(pe_4_15_go),
        .left(pe_4_15_left),
        .out(pe_4_15_out),
        .top(pe_4_15_top)
    );
    std_reg # (
        .width(32)
    ) top_4_15 (
        .clk(top_4_15_clk),
        .done(top_4_15_done),
        .in(top_4_15_in),
        .out(top_4_15_out),
        .write_en(top_4_15_write_en)
    );
    std_reg # (
        .width(32)
    ) left_4_15 (
        .clk(left_4_15_clk),
        .done(left_4_15_done),
        .in(left_4_15_in),
        .out(left_4_15_out),
        .write_en(left_4_15_write_en)
    );
    mac_pe pe_5_0 (
        .clk(pe_5_0_clk),
        .done(pe_5_0_done),
        .go(pe_5_0_go),
        .left(pe_5_0_left),
        .out(pe_5_0_out),
        .top(pe_5_0_top)
    );
    std_reg # (
        .width(32)
    ) top_5_0 (
        .clk(top_5_0_clk),
        .done(top_5_0_done),
        .in(top_5_0_in),
        .out(top_5_0_out),
        .write_en(top_5_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_0 (
        .clk(left_5_0_clk),
        .done(left_5_0_done),
        .in(left_5_0_in),
        .out(left_5_0_out),
        .write_en(left_5_0_write_en)
    );
    mac_pe pe_5_1 (
        .clk(pe_5_1_clk),
        .done(pe_5_1_done),
        .go(pe_5_1_go),
        .left(pe_5_1_left),
        .out(pe_5_1_out),
        .top(pe_5_1_top)
    );
    std_reg # (
        .width(32)
    ) top_5_1 (
        .clk(top_5_1_clk),
        .done(top_5_1_done),
        .in(top_5_1_in),
        .out(top_5_1_out),
        .write_en(top_5_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_1 (
        .clk(left_5_1_clk),
        .done(left_5_1_done),
        .in(left_5_1_in),
        .out(left_5_1_out),
        .write_en(left_5_1_write_en)
    );
    mac_pe pe_5_2 (
        .clk(pe_5_2_clk),
        .done(pe_5_2_done),
        .go(pe_5_2_go),
        .left(pe_5_2_left),
        .out(pe_5_2_out),
        .top(pe_5_2_top)
    );
    std_reg # (
        .width(32)
    ) top_5_2 (
        .clk(top_5_2_clk),
        .done(top_5_2_done),
        .in(top_5_2_in),
        .out(top_5_2_out),
        .write_en(top_5_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_2 (
        .clk(left_5_2_clk),
        .done(left_5_2_done),
        .in(left_5_2_in),
        .out(left_5_2_out),
        .write_en(left_5_2_write_en)
    );
    mac_pe pe_5_3 (
        .clk(pe_5_3_clk),
        .done(pe_5_3_done),
        .go(pe_5_3_go),
        .left(pe_5_3_left),
        .out(pe_5_3_out),
        .top(pe_5_3_top)
    );
    std_reg # (
        .width(32)
    ) top_5_3 (
        .clk(top_5_3_clk),
        .done(top_5_3_done),
        .in(top_5_3_in),
        .out(top_5_3_out),
        .write_en(top_5_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_3 (
        .clk(left_5_3_clk),
        .done(left_5_3_done),
        .in(left_5_3_in),
        .out(left_5_3_out),
        .write_en(left_5_3_write_en)
    );
    mac_pe pe_5_4 (
        .clk(pe_5_4_clk),
        .done(pe_5_4_done),
        .go(pe_5_4_go),
        .left(pe_5_4_left),
        .out(pe_5_4_out),
        .top(pe_5_4_top)
    );
    std_reg # (
        .width(32)
    ) top_5_4 (
        .clk(top_5_4_clk),
        .done(top_5_4_done),
        .in(top_5_4_in),
        .out(top_5_4_out),
        .write_en(top_5_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_4 (
        .clk(left_5_4_clk),
        .done(left_5_4_done),
        .in(left_5_4_in),
        .out(left_5_4_out),
        .write_en(left_5_4_write_en)
    );
    mac_pe pe_5_5 (
        .clk(pe_5_5_clk),
        .done(pe_5_5_done),
        .go(pe_5_5_go),
        .left(pe_5_5_left),
        .out(pe_5_5_out),
        .top(pe_5_5_top)
    );
    std_reg # (
        .width(32)
    ) top_5_5 (
        .clk(top_5_5_clk),
        .done(top_5_5_done),
        .in(top_5_5_in),
        .out(top_5_5_out),
        .write_en(top_5_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_5 (
        .clk(left_5_5_clk),
        .done(left_5_5_done),
        .in(left_5_5_in),
        .out(left_5_5_out),
        .write_en(left_5_5_write_en)
    );
    mac_pe pe_5_6 (
        .clk(pe_5_6_clk),
        .done(pe_5_6_done),
        .go(pe_5_6_go),
        .left(pe_5_6_left),
        .out(pe_5_6_out),
        .top(pe_5_6_top)
    );
    std_reg # (
        .width(32)
    ) top_5_6 (
        .clk(top_5_6_clk),
        .done(top_5_6_done),
        .in(top_5_6_in),
        .out(top_5_6_out),
        .write_en(top_5_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_6 (
        .clk(left_5_6_clk),
        .done(left_5_6_done),
        .in(left_5_6_in),
        .out(left_5_6_out),
        .write_en(left_5_6_write_en)
    );
    mac_pe pe_5_7 (
        .clk(pe_5_7_clk),
        .done(pe_5_7_done),
        .go(pe_5_7_go),
        .left(pe_5_7_left),
        .out(pe_5_7_out),
        .top(pe_5_7_top)
    );
    std_reg # (
        .width(32)
    ) top_5_7 (
        .clk(top_5_7_clk),
        .done(top_5_7_done),
        .in(top_5_7_in),
        .out(top_5_7_out),
        .write_en(top_5_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_7 (
        .clk(left_5_7_clk),
        .done(left_5_7_done),
        .in(left_5_7_in),
        .out(left_5_7_out),
        .write_en(left_5_7_write_en)
    );
    mac_pe pe_5_8 (
        .clk(pe_5_8_clk),
        .done(pe_5_8_done),
        .go(pe_5_8_go),
        .left(pe_5_8_left),
        .out(pe_5_8_out),
        .top(pe_5_8_top)
    );
    std_reg # (
        .width(32)
    ) top_5_8 (
        .clk(top_5_8_clk),
        .done(top_5_8_done),
        .in(top_5_8_in),
        .out(top_5_8_out),
        .write_en(top_5_8_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_8 (
        .clk(left_5_8_clk),
        .done(left_5_8_done),
        .in(left_5_8_in),
        .out(left_5_8_out),
        .write_en(left_5_8_write_en)
    );
    mac_pe pe_5_9 (
        .clk(pe_5_9_clk),
        .done(pe_5_9_done),
        .go(pe_5_9_go),
        .left(pe_5_9_left),
        .out(pe_5_9_out),
        .top(pe_5_9_top)
    );
    std_reg # (
        .width(32)
    ) top_5_9 (
        .clk(top_5_9_clk),
        .done(top_5_9_done),
        .in(top_5_9_in),
        .out(top_5_9_out),
        .write_en(top_5_9_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_9 (
        .clk(left_5_9_clk),
        .done(left_5_9_done),
        .in(left_5_9_in),
        .out(left_5_9_out),
        .write_en(left_5_9_write_en)
    );
    mac_pe pe_5_10 (
        .clk(pe_5_10_clk),
        .done(pe_5_10_done),
        .go(pe_5_10_go),
        .left(pe_5_10_left),
        .out(pe_5_10_out),
        .top(pe_5_10_top)
    );
    std_reg # (
        .width(32)
    ) top_5_10 (
        .clk(top_5_10_clk),
        .done(top_5_10_done),
        .in(top_5_10_in),
        .out(top_5_10_out),
        .write_en(top_5_10_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_10 (
        .clk(left_5_10_clk),
        .done(left_5_10_done),
        .in(left_5_10_in),
        .out(left_5_10_out),
        .write_en(left_5_10_write_en)
    );
    mac_pe pe_5_11 (
        .clk(pe_5_11_clk),
        .done(pe_5_11_done),
        .go(pe_5_11_go),
        .left(pe_5_11_left),
        .out(pe_5_11_out),
        .top(pe_5_11_top)
    );
    std_reg # (
        .width(32)
    ) top_5_11 (
        .clk(top_5_11_clk),
        .done(top_5_11_done),
        .in(top_5_11_in),
        .out(top_5_11_out),
        .write_en(top_5_11_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_11 (
        .clk(left_5_11_clk),
        .done(left_5_11_done),
        .in(left_5_11_in),
        .out(left_5_11_out),
        .write_en(left_5_11_write_en)
    );
    mac_pe pe_5_12 (
        .clk(pe_5_12_clk),
        .done(pe_5_12_done),
        .go(pe_5_12_go),
        .left(pe_5_12_left),
        .out(pe_5_12_out),
        .top(pe_5_12_top)
    );
    std_reg # (
        .width(32)
    ) top_5_12 (
        .clk(top_5_12_clk),
        .done(top_5_12_done),
        .in(top_5_12_in),
        .out(top_5_12_out),
        .write_en(top_5_12_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_12 (
        .clk(left_5_12_clk),
        .done(left_5_12_done),
        .in(left_5_12_in),
        .out(left_5_12_out),
        .write_en(left_5_12_write_en)
    );
    mac_pe pe_5_13 (
        .clk(pe_5_13_clk),
        .done(pe_5_13_done),
        .go(pe_5_13_go),
        .left(pe_5_13_left),
        .out(pe_5_13_out),
        .top(pe_5_13_top)
    );
    std_reg # (
        .width(32)
    ) top_5_13 (
        .clk(top_5_13_clk),
        .done(top_5_13_done),
        .in(top_5_13_in),
        .out(top_5_13_out),
        .write_en(top_5_13_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_13 (
        .clk(left_5_13_clk),
        .done(left_5_13_done),
        .in(left_5_13_in),
        .out(left_5_13_out),
        .write_en(left_5_13_write_en)
    );
    mac_pe pe_5_14 (
        .clk(pe_5_14_clk),
        .done(pe_5_14_done),
        .go(pe_5_14_go),
        .left(pe_5_14_left),
        .out(pe_5_14_out),
        .top(pe_5_14_top)
    );
    std_reg # (
        .width(32)
    ) top_5_14 (
        .clk(top_5_14_clk),
        .done(top_5_14_done),
        .in(top_5_14_in),
        .out(top_5_14_out),
        .write_en(top_5_14_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_14 (
        .clk(left_5_14_clk),
        .done(left_5_14_done),
        .in(left_5_14_in),
        .out(left_5_14_out),
        .write_en(left_5_14_write_en)
    );
    mac_pe pe_5_15 (
        .clk(pe_5_15_clk),
        .done(pe_5_15_done),
        .go(pe_5_15_go),
        .left(pe_5_15_left),
        .out(pe_5_15_out),
        .top(pe_5_15_top)
    );
    std_reg # (
        .width(32)
    ) top_5_15 (
        .clk(top_5_15_clk),
        .done(top_5_15_done),
        .in(top_5_15_in),
        .out(top_5_15_out),
        .write_en(top_5_15_write_en)
    );
    std_reg # (
        .width(32)
    ) left_5_15 (
        .clk(left_5_15_clk),
        .done(left_5_15_done),
        .in(left_5_15_in),
        .out(left_5_15_out),
        .write_en(left_5_15_write_en)
    );
    mac_pe pe_6_0 (
        .clk(pe_6_0_clk),
        .done(pe_6_0_done),
        .go(pe_6_0_go),
        .left(pe_6_0_left),
        .out(pe_6_0_out),
        .top(pe_6_0_top)
    );
    std_reg # (
        .width(32)
    ) top_6_0 (
        .clk(top_6_0_clk),
        .done(top_6_0_done),
        .in(top_6_0_in),
        .out(top_6_0_out),
        .write_en(top_6_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_0 (
        .clk(left_6_0_clk),
        .done(left_6_0_done),
        .in(left_6_0_in),
        .out(left_6_0_out),
        .write_en(left_6_0_write_en)
    );
    mac_pe pe_6_1 (
        .clk(pe_6_1_clk),
        .done(pe_6_1_done),
        .go(pe_6_1_go),
        .left(pe_6_1_left),
        .out(pe_6_1_out),
        .top(pe_6_1_top)
    );
    std_reg # (
        .width(32)
    ) top_6_1 (
        .clk(top_6_1_clk),
        .done(top_6_1_done),
        .in(top_6_1_in),
        .out(top_6_1_out),
        .write_en(top_6_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_1 (
        .clk(left_6_1_clk),
        .done(left_6_1_done),
        .in(left_6_1_in),
        .out(left_6_1_out),
        .write_en(left_6_1_write_en)
    );
    mac_pe pe_6_2 (
        .clk(pe_6_2_clk),
        .done(pe_6_2_done),
        .go(pe_6_2_go),
        .left(pe_6_2_left),
        .out(pe_6_2_out),
        .top(pe_6_2_top)
    );
    std_reg # (
        .width(32)
    ) top_6_2 (
        .clk(top_6_2_clk),
        .done(top_6_2_done),
        .in(top_6_2_in),
        .out(top_6_2_out),
        .write_en(top_6_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_2 (
        .clk(left_6_2_clk),
        .done(left_6_2_done),
        .in(left_6_2_in),
        .out(left_6_2_out),
        .write_en(left_6_2_write_en)
    );
    mac_pe pe_6_3 (
        .clk(pe_6_3_clk),
        .done(pe_6_3_done),
        .go(pe_6_3_go),
        .left(pe_6_3_left),
        .out(pe_6_3_out),
        .top(pe_6_3_top)
    );
    std_reg # (
        .width(32)
    ) top_6_3 (
        .clk(top_6_3_clk),
        .done(top_6_3_done),
        .in(top_6_3_in),
        .out(top_6_3_out),
        .write_en(top_6_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_3 (
        .clk(left_6_3_clk),
        .done(left_6_3_done),
        .in(left_6_3_in),
        .out(left_6_3_out),
        .write_en(left_6_3_write_en)
    );
    mac_pe pe_6_4 (
        .clk(pe_6_4_clk),
        .done(pe_6_4_done),
        .go(pe_6_4_go),
        .left(pe_6_4_left),
        .out(pe_6_4_out),
        .top(pe_6_4_top)
    );
    std_reg # (
        .width(32)
    ) top_6_4 (
        .clk(top_6_4_clk),
        .done(top_6_4_done),
        .in(top_6_4_in),
        .out(top_6_4_out),
        .write_en(top_6_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_4 (
        .clk(left_6_4_clk),
        .done(left_6_4_done),
        .in(left_6_4_in),
        .out(left_6_4_out),
        .write_en(left_6_4_write_en)
    );
    mac_pe pe_6_5 (
        .clk(pe_6_5_clk),
        .done(pe_6_5_done),
        .go(pe_6_5_go),
        .left(pe_6_5_left),
        .out(pe_6_5_out),
        .top(pe_6_5_top)
    );
    std_reg # (
        .width(32)
    ) top_6_5 (
        .clk(top_6_5_clk),
        .done(top_6_5_done),
        .in(top_6_5_in),
        .out(top_6_5_out),
        .write_en(top_6_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_5 (
        .clk(left_6_5_clk),
        .done(left_6_5_done),
        .in(left_6_5_in),
        .out(left_6_5_out),
        .write_en(left_6_5_write_en)
    );
    mac_pe pe_6_6 (
        .clk(pe_6_6_clk),
        .done(pe_6_6_done),
        .go(pe_6_6_go),
        .left(pe_6_6_left),
        .out(pe_6_6_out),
        .top(pe_6_6_top)
    );
    std_reg # (
        .width(32)
    ) top_6_6 (
        .clk(top_6_6_clk),
        .done(top_6_6_done),
        .in(top_6_6_in),
        .out(top_6_6_out),
        .write_en(top_6_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_6 (
        .clk(left_6_6_clk),
        .done(left_6_6_done),
        .in(left_6_6_in),
        .out(left_6_6_out),
        .write_en(left_6_6_write_en)
    );
    mac_pe pe_6_7 (
        .clk(pe_6_7_clk),
        .done(pe_6_7_done),
        .go(pe_6_7_go),
        .left(pe_6_7_left),
        .out(pe_6_7_out),
        .top(pe_6_7_top)
    );
    std_reg # (
        .width(32)
    ) top_6_7 (
        .clk(top_6_7_clk),
        .done(top_6_7_done),
        .in(top_6_7_in),
        .out(top_6_7_out),
        .write_en(top_6_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_7 (
        .clk(left_6_7_clk),
        .done(left_6_7_done),
        .in(left_6_7_in),
        .out(left_6_7_out),
        .write_en(left_6_7_write_en)
    );
    mac_pe pe_6_8 (
        .clk(pe_6_8_clk),
        .done(pe_6_8_done),
        .go(pe_6_8_go),
        .left(pe_6_8_left),
        .out(pe_6_8_out),
        .top(pe_6_8_top)
    );
    std_reg # (
        .width(32)
    ) top_6_8 (
        .clk(top_6_8_clk),
        .done(top_6_8_done),
        .in(top_6_8_in),
        .out(top_6_8_out),
        .write_en(top_6_8_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_8 (
        .clk(left_6_8_clk),
        .done(left_6_8_done),
        .in(left_6_8_in),
        .out(left_6_8_out),
        .write_en(left_6_8_write_en)
    );
    mac_pe pe_6_9 (
        .clk(pe_6_9_clk),
        .done(pe_6_9_done),
        .go(pe_6_9_go),
        .left(pe_6_9_left),
        .out(pe_6_9_out),
        .top(pe_6_9_top)
    );
    std_reg # (
        .width(32)
    ) top_6_9 (
        .clk(top_6_9_clk),
        .done(top_6_9_done),
        .in(top_6_9_in),
        .out(top_6_9_out),
        .write_en(top_6_9_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_9 (
        .clk(left_6_9_clk),
        .done(left_6_9_done),
        .in(left_6_9_in),
        .out(left_6_9_out),
        .write_en(left_6_9_write_en)
    );
    mac_pe pe_6_10 (
        .clk(pe_6_10_clk),
        .done(pe_6_10_done),
        .go(pe_6_10_go),
        .left(pe_6_10_left),
        .out(pe_6_10_out),
        .top(pe_6_10_top)
    );
    std_reg # (
        .width(32)
    ) top_6_10 (
        .clk(top_6_10_clk),
        .done(top_6_10_done),
        .in(top_6_10_in),
        .out(top_6_10_out),
        .write_en(top_6_10_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_10 (
        .clk(left_6_10_clk),
        .done(left_6_10_done),
        .in(left_6_10_in),
        .out(left_6_10_out),
        .write_en(left_6_10_write_en)
    );
    mac_pe pe_6_11 (
        .clk(pe_6_11_clk),
        .done(pe_6_11_done),
        .go(pe_6_11_go),
        .left(pe_6_11_left),
        .out(pe_6_11_out),
        .top(pe_6_11_top)
    );
    std_reg # (
        .width(32)
    ) top_6_11 (
        .clk(top_6_11_clk),
        .done(top_6_11_done),
        .in(top_6_11_in),
        .out(top_6_11_out),
        .write_en(top_6_11_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_11 (
        .clk(left_6_11_clk),
        .done(left_6_11_done),
        .in(left_6_11_in),
        .out(left_6_11_out),
        .write_en(left_6_11_write_en)
    );
    mac_pe pe_6_12 (
        .clk(pe_6_12_clk),
        .done(pe_6_12_done),
        .go(pe_6_12_go),
        .left(pe_6_12_left),
        .out(pe_6_12_out),
        .top(pe_6_12_top)
    );
    std_reg # (
        .width(32)
    ) top_6_12 (
        .clk(top_6_12_clk),
        .done(top_6_12_done),
        .in(top_6_12_in),
        .out(top_6_12_out),
        .write_en(top_6_12_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_12 (
        .clk(left_6_12_clk),
        .done(left_6_12_done),
        .in(left_6_12_in),
        .out(left_6_12_out),
        .write_en(left_6_12_write_en)
    );
    mac_pe pe_6_13 (
        .clk(pe_6_13_clk),
        .done(pe_6_13_done),
        .go(pe_6_13_go),
        .left(pe_6_13_left),
        .out(pe_6_13_out),
        .top(pe_6_13_top)
    );
    std_reg # (
        .width(32)
    ) top_6_13 (
        .clk(top_6_13_clk),
        .done(top_6_13_done),
        .in(top_6_13_in),
        .out(top_6_13_out),
        .write_en(top_6_13_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_13 (
        .clk(left_6_13_clk),
        .done(left_6_13_done),
        .in(left_6_13_in),
        .out(left_6_13_out),
        .write_en(left_6_13_write_en)
    );
    mac_pe pe_6_14 (
        .clk(pe_6_14_clk),
        .done(pe_6_14_done),
        .go(pe_6_14_go),
        .left(pe_6_14_left),
        .out(pe_6_14_out),
        .top(pe_6_14_top)
    );
    std_reg # (
        .width(32)
    ) top_6_14 (
        .clk(top_6_14_clk),
        .done(top_6_14_done),
        .in(top_6_14_in),
        .out(top_6_14_out),
        .write_en(top_6_14_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_14 (
        .clk(left_6_14_clk),
        .done(left_6_14_done),
        .in(left_6_14_in),
        .out(left_6_14_out),
        .write_en(left_6_14_write_en)
    );
    mac_pe pe_6_15 (
        .clk(pe_6_15_clk),
        .done(pe_6_15_done),
        .go(pe_6_15_go),
        .left(pe_6_15_left),
        .out(pe_6_15_out),
        .top(pe_6_15_top)
    );
    std_reg # (
        .width(32)
    ) top_6_15 (
        .clk(top_6_15_clk),
        .done(top_6_15_done),
        .in(top_6_15_in),
        .out(top_6_15_out),
        .write_en(top_6_15_write_en)
    );
    std_reg # (
        .width(32)
    ) left_6_15 (
        .clk(left_6_15_clk),
        .done(left_6_15_done),
        .in(left_6_15_in),
        .out(left_6_15_out),
        .write_en(left_6_15_write_en)
    );
    mac_pe pe_7_0 (
        .clk(pe_7_0_clk),
        .done(pe_7_0_done),
        .go(pe_7_0_go),
        .left(pe_7_0_left),
        .out(pe_7_0_out),
        .top(pe_7_0_top)
    );
    std_reg # (
        .width(32)
    ) top_7_0 (
        .clk(top_7_0_clk),
        .done(top_7_0_done),
        .in(top_7_0_in),
        .out(top_7_0_out),
        .write_en(top_7_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_0 (
        .clk(left_7_0_clk),
        .done(left_7_0_done),
        .in(left_7_0_in),
        .out(left_7_0_out),
        .write_en(left_7_0_write_en)
    );
    mac_pe pe_7_1 (
        .clk(pe_7_1_clk),
        .done(pe_7_1_done),
        .go(pe_7_1_go),
        .left(pe_7_1_left),
        .out(pe_7_1_out),
        .top(pe_7_1_top)
    );
    std_reg # (
        .width(32)
    ) top_7_1 (
        .clk(top_7_1_clk),
        .done(top_7_1_done),
        .in(top_7_1_in),
        .out(top_7_1_out),
        .write_en(top_7_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_1 (
        .clk(left_7_1_clk),
        .done(left_7_1_done),
        .in(left_7_1_in),
        .out(left_7_1_out),
        .write_en(left_7_1_write_en)
    );
    mac_pe pe_7_2 (
        .clk(pe_7_2_clk),
        .done(pe_7_2_done),
        .go(pe_7_2_go),
        .left(pe_7_2_left),
        .out(pe_7_2_out),
        .top(pe_7_2_top)
    );
    std_reg # (
        .width(32)
    ) top_7_2 (
        .clk(top_7_2_clk),
        .done(top_7_2_done),
        .in(top_7_2_in),
        .out(top_7_2_out),
        .write_en(top_7_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_2 (
        .clk(left_7_2_clk),
        .done(left_7_2_done),
        .in(left_7_2_in),
        .out(left_7_2_out),
        .write_en(left_7_2_write_en)
    );
    mac_pe pe_7_3 (
        .clk(pe_7_3_clk),
        .done(pe_7_3_done),
        .go(pe_7_3_go),
        .left(pe_7_3_left),
        .out(pe_7_3_out),
        .top(pe_7_3_top)
    );
    std_reg # (
        .width(32)
    ) top_7_3 (
        .clk(top_7_3_clk),
        .done(top_7_3_done),
        .in(top_7_3_in),
        .out(top_7_3_out),
        .write_en(top_7_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_3 (
        .clk(left_7_3_clk),
        .done(left_7_3_done),
        .in(left_7_3_in),
        .out(left_7_3_out),
        .write_en(left_7_3_write_en)
    );
    mac_pe pe_7_4 (
        .clk(pe_7_4_clk),
        .done(pe_7_4_done),
        .go(pe_7_4_go),
        .left(pe_7_4_left),
        .out(pe_7_4_out),
        .top(pe_7_4_top)
    );
    std_reg # (
        .width(32)
    ) top_7_4 (
        .clk(top_7_4_clk),
        .done(top_7_4_done),
        .in(top_7_4_in),
        .out(top_7_4_out),
        .write_en(top_7_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_4 (
        .clk(left_7_4_clk),
        .done(left_7_4_done),
        .in(left_7_4_in),
        .out(left_7_4_out),
        .write_en(left_7_4_write_en)
    );
    mac_pe pe_7_5 (
        .clk(pe_7_5_clk),
        .done(pe_7_5_done),
        .go(pe_7_5_go),
        .left(pe_7_5_left),
        .out(pe_7_5_out),
        .top(pe_7_5_top)
    );
    std_reg # (
        .width(32)
    ) top_7_5 (
        .clk(top_7_5_clk),
        .done(top_7_5_done),
        .in(top_7_5_in),
        .out(top_7_5_out),
        .write_en(top_7_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_5 (
        .clk(left_7_5_clk),
        .done(left_7_5_done),
        .in(left_7_5_in),
        .out(left_7_5_out),
        .write_en(left_7_5_write_en)
    );
    mac_pe pe_7_6 (
        .clk(pe_7_6_clk),
        .done(pe_7_6_done),
        .go(pe_7_6_go),
        .left(pe_7_6_left),
        .out(pe_7_6_out),
        .top(pe_7_6_top)
    );
    std_reg # (
        .width(32)
    ) top_7_6 (
        .clk(top_7_6_clk),
        .done(top_7_6_done),
        .in(top_7_6_in),
        .out(top_7_6_out),
        .write_en(top_7_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_6 (
        .clk(left_7_6_clk),
        .done(left_7_6_done),
        .in(left_7_6_in),
        .out(left_7_6_out),
        .write_en(left_7_6_write_en)
    );
    mac_pe pe_7_7 (
        .clk(pe_7_7_clk),
        .done(pe_7_7_done),
        .go(pe_7_7_go),
        .left(pe_7_7_left),
        .out(pe_7_7_out),
        .top(pe_7_7_top)
    );
    std_reg # (
        .width(32)
    ) top_7_7 (
        .clk(top_7_7_clk),
        .done(top_7_7_done),
        .in(top_7_7_in),
        .out(top_7_7_out),
        .write_en(top_7_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_7 (
        .clk(left_7_7_clk),
        .done(left_7_7_done),
        .in(left_7_7_in),
        .out(left_7_7_out),
        .write_en(left_7_7_write_en)
    );
    mac_pe pe_7_8 (
        .clk(pe_7_8_clk),
        .done(pe_7_8_done),
        .go(pe_7_8_go),
        .left(pe_7_8_left),
        .out(pe_7_8_out),
        .top(pe_7_8_top)
    );
    std_reg # (
        .width(32)
    ) top_7_8 (
        .clk(top_7_8_clk),
        .done(top_7_8_done),
        .in(top_7_8_in),
        .out(top_7_8_out),
        .write_en(top_7_8_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_8 (
        .clk(left_7_8_clk),
        .done(left_7_8_done),
        .in(left_7_8_in),
        .out(left_7_8_out),
        .write_en(left_7_8_write_en)
    );
    mac_pe pe_7_9 (
        .clk(pe_7_9_clk),
        .done(pe_7_9_done),
        .go(pe_7_9_go),
        .left(pe_7_9_left),
        .out(pe_7_9_out),
        .top(pe_7_9_top)
    );
    std_reg # (
        .width(32)
    ) top_7_9 (
        .clk(top_7_9_clk),
        .done(top_7_9_done),
        .in(top_7_9_in),
        .out(top_7_9_out),
        .write_en(top_7_9_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_9 (
        .clk(left_7_9_clk),
        .done(left_7_9_done),
        .in(left_7_9_in),
        .out(left_7_9_out),
        .write_en(left_7_9_write_en)
    );
    mac_pe pe_7_10 (
        .clk(pe_7_10_clk),
        .done(pe_7_10_done),
        .go(pe_7_10_go),
        .left(pe_7_10_left),
        .out(pe_7_10_out),
        .top(pe_7_10_top)
    );
    std_reg # (
        .width(32)
    ) top_7_10 (
        .clk(top_7_10_clk),
        .done(top_7_10_done),
        .in(top_7_10_in),
        .out(top_7_10_out),
        .write_en(top_7_10_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_10 (
        .clk(left_7_10_clk),
        .done(left_7_10_done),
        .in(left_7_10_in),
        .out(left_7_10_out),
        .write_en(left_7_10_write_en)
    );
    mac_pe pe_7_11 (
        .clk(pe_7_11_clk),
        .done(pe_7_11_done),
        .go(pe_7_11_go),
        .left(pe_7_11_left),
        .out(pe_7_11_out),
        .top(pe_7_11_top)
    );
    std_reg # (
        .width(32)
    ) top_7_11 (
        .clk(top_7_11_clk),
        .done(top_7_11_done),
        .in(top_7_11_in),
        .out(top_7_11_out),
        .write_en(top_7_11_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_11 (
        .clk(left_7_11_clk),
        .done(left_7_11_done),
        .in(left_7_11_in),
        .out(left_7_11_out),
        .write_en(left_7_11_write_en)
    );
    mac_pe pe_7_12 (
        .clk(pe_7_12_clk),
        .done(pe_7_12_done),
        .go(pe_7_12_go),
        .left(pe_7_12_left),
        .out(pe_7_12_out),
        .top(pe_7_12_top)
    );
    std_reg # (
        .width(32)
    ) top_7_12 (
        .clk(top_7_12_clk),
        .done(top_7_12_done),
        .in(top_7_12_in),
        .out(top_7_12_out),
        .write_en(top_7_12_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_12 (
        .clk(left_7_12_clk),
        .done(left_7_12_done),
        .in(left_7_12_in),
        .out(left_7_12_out),
        .write_en(left_7_12_write_en)
    );
    mac_pe pe_7_13 (
        .clk(pe_7_13_clk),
        .done(pe_7_13_done),
        .go(pe_7_13_go),
        .left(pe_7_13_left),
        .out(pe_7_13_out),
        .top(pe_7_13_top)
    );
    std_reg # (
        .width(32)
    ) top_7_13 (
        .clk(top_7_13_clk),
        .done(top_7_13_done),
        .in(top_7_13_in),
        .out(top_7_13_out),
        .write_en(top_7_13_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_13 (
        .clk(left_7_13_clk),
        .done(left_7_13_done),
        .in(left_7_13_in),
        .out(left_7_13_out),
        .write_en(left_7_13_write_en)
    );
    mac_pe pe_7_14 (
        .clk(pe_7_14_clk),
        .done(pe_7_14_done),
        .go(pe_7_14_go),
        .left(pe_7_14_left),
        .out(pe_7_14_out),
        .top(pe_7_14_top)
    );
    std_reg # (
        .width(32)
    ) top_7_14 (
        .clk(top_7_14_clk),
        .done(top_7_14_done),
        .in(top_7_14_in),
        .out(top_7_14_out),
        .write_en(top_7_14_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_14 (
        .clk(left_7_14_clk),
        .done(left_7_14_done),
        .in(left_7_14_in),
        .out(left_7_14_out),
        .write_en(left_7_14_write_en)
    );
    mac_pe pe_7_15 (
        .clk(pe_7_15_clk),
        .done(pe_7_15_done),
        .go(pe_7_15_go),
        .left(pe_7_15_left),
        .out(pe_7_15_out),
        .top(pe_7_15_top)
    );
    std_reg # (
        .width(32)
    ) top_7_15 (
        .clk(top_7_15_clk),
        .done(top_7_15_done),
        .in(top_7_15_in),
        .out(top_7_15_out),
        .write_en(top_7_15_write_en)
    );
    std_reg # (
        .width(32)
    ) left_7_15 (
        .clk(left_7_15_clk),
        .done(left_7_15_done),
        .in(left_7_15_in),
        .out(left_7_15_out),
        .write_en(left_7_15_write_en)
    );
    mac_pe pe_8_0 (
        .clk(pe_8_0_clk),
        .done(pe_8_0_done),
        .go(pe_8_0_go),
        .left(pe_8_0_left),
        .out(pe_8_0_out),
        .top(pe_8_0_top)
    );
    std_reg # (
        .width(32)
    ) top_8_0 (
        .clk(top_8_0_clk),
        .done(top_8_0_done),
        .in(top_8_0_in),
        .out(top_8_0_out),
        .write_en(top_8_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_8_0 (
        .clk(left_8_0_clk),
        .done(left_8_0_done),
        .in(left_8_0_in),
        .out(left_8_0_out),
        .write_en(left_8_0_write_en)
    );
    mac_pe pe_8_1 (
        .clk(pe_8_1_clk),
        .done(pe_8_1_done),
        .go(pe_8_1_go),
        .left(pe_8_1_left),
        .out(pe_8_1_out),
        .top(pe_8_1_top)
    );
    std_reg # (
        .width(32)
    ) top_8_1 (
        .clk(top_8_1_clk),
        .done(top_8_1_done),
        .in(top_8_1_in),
        .out(top_8_1_out),
        .write_en(top_8_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_8_1 (
        .clk(left_8_1_clk),
        .done(left_8_1_done),
        .in(left_8_1_in),
        .out(left_8_1_out),
        .write_en(left_8_1_write_en)
    );
    mac_pe pe_8_2 (
        .clk(pe_8_2_clk),
        .done(pe_8_2_done),
        .go(pe_8_2_go),
        .left(pe_8_2_left),
        .out(pe_8_2_out),
        .top(pe_8_2_top)
    );
    std_reg # (
        .width(32)
    ) top_8_2 (
        .clk(top_8_2_clk),
        .done(top_8_2_done),
        .in(top_8_2_in),
        .out(top_8_2_out),
        .write_en(top_8_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_8_2 (
        .clk(left_8_2_clk),
        .done(left_8_2_done),
        .in(left_8_2_in),
        .out(left_8_2_out),
        .write_en(left_8_2_write_en)
    );
    mac_pe pe_8_3 (
        .clk(pe_8_3_clk),
        .done(pe_8_3_done),
        .go(pe_8_3_go),
        .left(pe_8_3_left),
        .out(pe_8_3_out),
        .top(pe_8_3_top)
    );
    std_reg # (
        .width(32)
    ) top_8_3 (
        .clk(top_8_3_clk),
        .done(top_8_3_done),
        .in(top_8_3_in),
        .out(top_8_3_out),
        .write_en(top_8_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_8_3 (
        .clk(left_8_3_clk),
        .done(left_8_3_done),
        .in(left_8_3_in),
        .out(left_8_3_out),
        .write_en(left_8_3_write_en)
    );
    mac_pe pe_8_4 (
        .clk(pe_8_4_clk),
        .done(pe_8_4_done),
        .go(pe_8_4_go),
        .left(pe_8_4_left),
        .out(pe_8_4_out),
        .top(pe_8_4_top)
    );
    std_reg # (
        .width(32)
    ) top_8_4 (
        .clk(top_8_4_clk),
        .done(top_8_4_done),
        .in(top_8_4_in),
        .out(top_8_4_out),
        .write_en(top_8_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_8_4 (
        .clk(left_8_4_clk),
        .done(left_8_4_done),
        .in(left_8_4_in),
        .out(left_8_4_out),
        .write_en(left_8_4_write_en)
    );
    mac_pe pe_8_5 (
        .clk(pe_8_5_clk),
        .done(pe_8_5_done),
        .go(pe_8_5_go),
        .left(pe_8_5_left),
        .out(pe_8_5_out),
        .top(pe_8_5_top)
    );
    std_reg # (
        .width(32)
    ) top_8_5 (
        .clk(top_8_5_clk),
        .done(top_8_5_done),
        .in(top_8_5_in),
        .out(top_8_5_out),
        .write_en(top_8_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_8_5 (
        .clk(left_8_5_clk),
        .done(left_8_5_done),
        .in(left_8_5_in),
        .out(left_8_5_out),
        .write_en(left_8_5_write_en)
    );
    mac_pe pe_8_6 (
        .clk(pe_8_6_clk),
        .done(pe_8_6_done),
        .go(pe_8_6_go),
        .left(pe_8_6_left),
        .out(pe_8_6_out),
        .top(pe_8_6_top)
    );
    std_reg # (
        .width(32)
    ) top_8_6 (
        .clk(top_8_6_clk),
        .done(top_8_6_done),
        .in(top_8_6_in),
        .out(top_8_6_out),
        .write_en(top_8_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_8_6 (
        .clk(left_8_6_clk),
        .done(left_8_6_done),
        .in(left_8_6_in),
        .out(left_8_6_out),
        .write_en(left_8_6_write_en)
    );
    mac_pe pe_8_7 (
        .clk(pe_8_7_clk),
        .done(pe_8_7_done),
        .go(pe_8_7_go),
        .left(pe_8_7_left),
        .out(pe_8_7_out),
        .top(pe_8_7_top)
    );
    std_reg # (
        .width(32)
    ) top_8_7 (
        .clk(top_8_7_clk),
        .done(top_8_7_done),
        .in(top_8_7_in),
        .out(top_8_7_out),
        .write_en(top_8_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_8_7 (
        .clk(left_8_7_clk),
        .done(left_8_7_done),
        .in(left_8_7_in),
        .out(left_8_7_out),
        .write_en(left_8_7_write_en)
    );
    mac_pe pe_8_8 (
        .clk(pe_8_8_clk),
        .done(pe_8_8_done),
        .go(pe_8_8_go),
        .left(pe_8_8_left),
        .out(pe_8_8_out),
        .top(pe_8_8_top)
    );
    std_reg # (
        .width(32)
    ) top_8_8 (
        .clk(top_8_8_clk),
        .done(top_8_8_done),
        .in(top_8_8_in),
        .out(top_8_8_out),
        .write_en(top_8_8_write_en)
    );
    std_reg # (
        .width(32)
    ) left_8_8 (
        .clk(left_8_8_clk),
        .done(left_8_8_done),
        .in(left_8_8_in),
        .out(left_8_8_out),
        .write_en(left_8_8_write_en)
    );
    mac_pe pe_8_9 (
        .clk(pe_8_9_clk),
        .done(pe_8_9_done),
        .go(pe_8_9_go),
        .left(pe_8_9_left),
        .out(pe_8_9_out),
        .top(pe_8_9_top)
    );
    std_reg # (
        .width(32)
    ) top_8_9 (
        .clk(top_8_9_clk),
        .done(top_8_9_done),
        .in(top_8_9_in),
        .out(top_8_9_out),
        .write_en(top_8_9_write_en)
    );
    std_reg # (
        .width(32)
    ) left_8_9 (
        .clk(left_8_9_clk),
        .done(left_8_9_done),
        .in(left_8_9_in),
        .out(left_8_9_out),
        .write_en(left_8_9_write_en)
    );
    mac_pe pe_8_10 (
        .clk(pe_8_10_clk),
        .done(pe_8_10_done),
        .go(pe_8_10_go),
        .left(pe_8_10_left),
        .out(pe_8_10_out),
        .top(pe_8_10_top)
    );
    std_reg # (
        .width(32)
    ) top_8_10 (
        .clk(top_8_10_clk),
        .done(top_8_10_done),
        .in(top_8_10_in),
        .out(top_8_10_out),
        .write_en(top_8_10_write_en)
    );
    std_reg # (
        .width(32)
    ) left_8_10 (
        .clk(left_8_10_clk),
        .done(left_8_10_done),
        .in(left_8_10_in),
        .out(left_8_10_out),
        .write_en(left_8_10_write_en)
    );
    mac_pe pe_8_11 (
        .clk(pe_8_11_clk),
        .done(pe_8_11_done),
        .go(pe_8_11_go),
        .left(pe_8_11_left),
        .out(pe_8_11_out),
        .top(pe_8_11_top)
    );
    std_reg # (
        .width(32)
    ) top_8_11 (
        .clk(top_8_11_clk),
        .done(top_8_11_done),
        .in(top_8_11_in),
        .out(top_8_11_out),
        .write_en(top_8_11_write_en)
    );
    std_reg # (
        .width(32)
    ) left_8_11 (
        .clk(left_8_11_clk),
        .done(left_8_11_done),
        .in(left_8_11_in),
        .out(left_8_11_out),
        .write_en(left_8_11_write_en)
    );
    mac_pe pe_8_12 (
        .clk(pe_8_12_clk),
        .done(pe_8_12_done),
        .go(pe_8_12_go),
        .left(pe_8_12_left),
        .out(pe_8_12_out),
        .top(pe_8_12_top)
    );
    std_reg # (
        .width(32)
    ) top_8_12 (
        .clk(top_8_12_clk),
        .done(top_8_12_done),
        .in(top_8_12_in),
        .out(top_8_12_out),
        .write_en(top_8_12_write_en)
    );
    std_reg # (
        .width(32)
    ) left_8_12 (
        .clk(left_8_12_clk),
        .done(left_8_12_done),
        .in(left_8_12_in),
        .out(left_8_12_out),
        .write_en(left_8_12_write_en)
    );
    mac_pe pe_8_13 (
        .clk(pe_8_13_clk),
        .done(pe_8_13_done),
        .go(pe_8_13_go),
        .left(pe_8_13_left),
        .out(pe_8_13_out),
        .top(pe_8_13_top)
    );
    std_reg # (
        .width(32)
    ) top_8_13 (
        .clk(top_8_13_clk),
        .done(top_8_13_done),
        .in(top_8_13_in),
        .out(top_8_13_out),
        .write_en(top_8_13_write_en)
    );
    std_reg # (
        .width(32)
    ) left_8_13 (
        .clk(left_8_13_clk),
        .done(left_8_13_done),
        .in(left_8_13_in),
        .out(left_8_13_out),
        .write_en(left_8_13_write_en)
    );
    mac_pe pe_8_14 (
        .clk(pe_8_14_clk),
        .done(pe_8_14_done),
        .go(pe_8_14_go),
        .left(pe_8_14_left),
        .out(pe_8_14_out),
        .top(pe_8_14_top)
    );
    std_reg # (
        .width(32)
    ) top_8_14 (
        .clk(top_8_14_clk),
        .done(top_8_14_done),
        .in(top_8_14_in),
        .out(top_8_14_out),
        .write_en(top_8_14_write_en)
    );
    std_reg # (
        .width(32)
    ) left_8_14 (
        .clk(left_8_14_clk),
        .done(left_8_14_done),
        .in(left_8_14_in),
        .out(left_8_14_out),
        .write_en(left_8_14_write_en)
    );
    mac_pe pe_8_15 (
        .clk(pe_8_15_clk),
        .done(pe_8_15_done),
        .go(pe_8_15_go),
        .left(pe_8_15_left),
        .out(pe_8_15_out),
        .top(pe_8_15_top)
    );
    std_reg # (
        .width(32)
    ) top_8_15 (
        .clk(top_8_15_clk),
        .done(top_8_15_done),
        .in(top_8_15_in),
        .out(top_8_15_out),
        .write_en(top_8_15_write_en)
    );
    std_reg # (
        .width(32)
    ) left_8_15 (
        .clk(left_8_15_clk),
        .done(left_8_15_done),
        .in(left_8_15_in),
        .out(left_8_15_out),
        .write_en(left_8_15_write_en)
    );
    mac_pe pe_9_0 (
        .clk(pe_9_0_clk),
        .done(pe_9_0_done),
        .go(pe_9_0_go),
        .left(pe_9_0_left),
        .out(pe_9_0_out),
        .top(pe_9_0_top)
    );
    std_reg # (
        .width(32)
    ) top_9_0 (
        .clk(top_9_0_clk),
        .done(top_9_0_done),
        .in(top_9_0_in),
        .out(top_9_0_out),
        .write_en(top_9_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_9_0 (
        .clk(left_9_0_clk),
        .done(left_9_0_done),
        .in(left_9_0_in),
        .out(left_9_0_out),
        .write_en(left_9_0_write_en)
    );
    mac_pe pe_9_1 (
        .clk(pe_9_1_clk),
        .done(pe_9_1_done),
        .go(pe_9_1_go),
        .left(pe_9_1_left),
        .out(pe_9_1_out),
        .top(pe_9_1_top)
    );
    std_reg # (
        .width(32)
    ) top_9_1 (
        .clk(top_9_1_clk),
        .done(top_9_1_done),
        .in(top_9_1_in),
        .out(top_9_1_out),
        .write_en(top_9_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_9_1 (
        .clk(left_9_1_clk),
        .done(left_9_1_done),
        .in(left_9_1_in),
        .out(left_9_1_out),
        .write_en(left_9_1_write_en)
    );
    mac_pe pe_9_2 (
        .clk(pe_9_2_clk),
        .done(pe_9_2_done),
        .go(pe_9_2_go),
        .left(pe_9_2_left),
        .out(pe_9_2_out),
        .top(pe_9_2_top)
    );
    std_reg # (
        .width(32)
    ) top_9_2 (
        .clk(top_9_2_clk),
        .done(top_9_2_done),
        .in(top_9_2_in),
        .out(top_9_2_out),
        .write_en(top_9_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_9_2 (
        .clk(left_9_2_clk),
        .done(left_9_2_done),
        .in(left_9_2_in),
        .out(left_9_2_out),
        .write_en(left_9_2_write_en)
    );
    mac_pe pe_9_3 (
        .clk(pe_9_3_clk),
        .done(pe_9_3_done),
        .go(pe_9_3_go),
        .left(pe_9_3_left),
        .out(pe_9_3_out),
        .top(pe_9_3_top)
    );
    std_reg # (
        .width(32)
    ) top_9_3 (
        .clk(top_9_3_clk),
        .done(top_9_3_done),
        .in(top_9_3_in),
        .out(top_9_3_out),
        .write_en(top_9_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_9_3 (
        .clk(left_9_3_clk),
        .done(left_9_3_done),
        .in(left_9_3_in),
        .out(left_9_3_out),
        .write_en(left_9_3_write_en)
    );
    mac_pe pe_9_4 (
        .clk(pe_9_4_clk),
        .done(pe_9_4_done),
        .go(pe_9_4_go),
        .left(pe_9_4_left),
        .out(pe_9_4_out),
        .top(pe_9_4_top)
    );
    std_reg # (
        .width(32)
    ) top_9_4 (
        .clk(top_9_4_clk),
        .done(top_9_4_done),
        .in(top_9_4_in),
        .out(top_9_4_out),
        .write_en(top_9_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_9_4 (
        .clk(left_9_4_clk),
        .done(left_9_4_done),
        .in(left_9_4_in),
        .out(left_9_4_out),
        .write_en(left_9_4_write_en)
    );
    mac_pe pe_9_5 (
        .clk(pe_9_5_clk),
        .done(pe_9_5_done),
        .go(pe_9_5_go),
        .left(pe_9_5_left),
        .out(pe_9_5_out),
        .top(pe_9_5_top)
    );
    std_reg # (
        .width(32)
    ) top_9_5 (
        .clk(top_9_5_clk),
        .done(top_9_5_done),
        .in(top_9_5_in),
        .out(top_9_5_out),
        .write_en(top_9_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_9_5 (
        .clk(left_9_5_clk),
        .done(left_9_5_done),
        .in(left_9_5_in),
        .out(left_9_5_out),
        .write_en(left_9_5_write_en)
    );
    mac_pe pe_9_6 (
        .clk(pe_9_6_clk),
        .done(pe_9_6_done),
        .go(pe_9_6_go),
        .left(pe_9_6_left),
        .out(pe_9_6_out),
        .top(pe_9_6_top)
    );
    std_reg # (
        .width(32)
    ) top_9_6 (
        .clk(top_9_6_clk),
        .done(top_9_6_done),
        .in(top_9_6_in),
        .out(top_9_6_out),
        .write_en(top_9_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_9_6 (
        .clk(left_9_6_clk),
        .done(left_9_6_done),
        .in(left_9_6_in),
        .out(left_9_6_out),
        .write_en(left_9_6_write_en)
    );
    mac_pe pe_9_7 (
        .clk(pe_9_7_clk),
        .done(pe_9_7_done),
        .go(pe_9_7_go),
        .left(pe_9_7_left),
        .out(pe_9_7_out),
        .top(pe_9_7_top)
    );
    std_reg # (
        .width(32)
    ) top_9_7 (
        .clk(top_9_7_clk),
        .done(top_9_7_done),
        .in(top_9_7_in),
        .out(top_9_7_out),
        .write_en(top_9_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_9_7 (
        .clk(left_9_7_clk),
        .done(left_9_7_done),
        .in(left_9_7_in),
        .out(left_9_7_out),
        .write_en(left_9_7_write_en)
    );
    mac_pe pe_9_8 (
        .clk(pe_9_8_clk),
        .done(pe_9_8_done),
        .go(pe_9_8_go),
        .left(pe_9_8_left),
        .out(pe_9_8_out),
        .top(pe_9_8_top)
    );
    std_reg # (
        .width(32)
    ) top_9_8 (
        .clk(top_9_8_clk),
        .done(top_9_8_done),
        .in(top_9_8_in),
        .out(top_9_8_out),
        .write_en(top_9_8_write_en)
    );
    std_reg # (
        .width(32)
    ) left_9_8 (
        .clk(left_9_8_clk),
        .done(left_9_8_done),
        .in(left_9_8_in),
        .out(left_9_8_out),
        .write_en(left_9_8_write_en)
    );
    mac_pe pe_9_9 (
        .clk(pe_9_9_clk),
        .done(pe_9_9_done),
        .go(pe_9_9_go),
        .left(pe_9_9_left),
        .out(pe_9_9_out),
        .top(pe_9_9_top)
    );
    std_reg # (
        .width(32)
    ) top_9_9 (
        .clk(top_9_9_clk),
        .done(top_9_9_done),
        .in(top_9_9_in),
        .out(top_9_9_out),
        .write_en(top_9_9_write_en)
    );
    std_reg # (
        .width(32)
    ) left_9_9 (
        .clk(left_9_9_clk),
        .done(left_9_9_done),
        .in(left_9_9_in),
        .out(left_9_9_out),
        .write_en(left_9_9_write_en)
    );
    mac_pe pe_9_10 (
        .clk(pe_9_10_clk),
        .done(pe_9_10_done),
        .go(pe_9_10_go),
        .left(pe_9_10_left),
        .out(pe_9_10_out),
        .top(pe_9_10_top)
    );
    std_reg # (
        .width(32)
    ) top_9_10 (
        .clk(top_9_10_clk),
        .done(top_9_10_done),
        .in(top_9_10_in),
        .out(top_9_10_out),
        .write_en(top_9_10_write_en)
    );
    std_reg # (
        .width(32)
    ) left_9_10 (
        .clk(left_9_10_clk),
        .done(left_9_10_done),
        .in(left_9_10_in),
        .out(left_9_10_out),
        .write_en(left_9_10_write_en)
    );
    mac_pe pe_9_11 (
        .clk(pe_9_11_clk),
        .done(pe_9_11_done),
        .go(pe_9_11_go),
        .left(pe_9_11_left),
        .out(pe_9_11_out),
        .top(pe_9_11_top)
    );
    std_reg # (
        .width(32)
    ) top_9_11 (
        .clk(top_9_11_clk),
        .done(top_9_11_done),
        .in(top_9_11_in),
        .out(top_9_11_out),
        .write_en(top_9_11_write_en)
    );
    std_reg # (
        .width(32)
    ) left_9_11 (
        .clk(left_9_11_clk),
        .done(left_9_11_done),
        .in(left_9_11_in),
        .out(left_9_11_out),
        .write_en(left_9_11_write_en)
    );
    mac_pe pe_9_12 (
        .clk(pe_9_12_clk),
        .done(pe_9_12_done),
        .go(pe_9_12_go),
        .left(pe_9_12_left),
        .out(pe_9_12_out),
        .top(pe_9_12_top)
    );
    std_reg # (
        .width(32)
    ) top_9_12 (
        .clk(top_9_12_clk),
        .done(top_9_12_done),
        .in(top_9_12_in),
        .out(top_9_12_out),
        .write_en(top_9_12_write_en)
    );
    std_reg # (
        .width(32)
    ) left_9_12 (
        .clk(left_9_12_clk),
        .done(left_9_12_done),
        .in(left_9_12_in),
        .out(left_9_12_out),
        .write_en(left_9_12_write_en)
    );
    mac_pe pe_9_13 (
        .clk(pe_9_13_clk),
        .done(pe_9_13_done),
        .go(pe_9_13_go),
        .left(pe_9_13_left),
        .out(pe_9_13_out),
        .top(pe_9_13_top)
    );
    std_reg # (
        .width(32)
    ) top_9_13 (
        .clk(top_9_13_clk),
        .done(top_9_13_done),
        .in(top_9_13_in),
        .out(top_9_13_out),
        .write_en(top_9_13_write_en)
    );
    std_reg # (
        .width(32)
    ) left_9_13 (
        .clk(left_9_13_clk),
        .done(left_9_13_done),
        .in(left_9_13_in),
        .out(left_9_13_out),
        .write_en(left_9_13_write_en)
    );
    mac_pe pe_9_14 (
        .clk(pe_9_14_clk),
        .done(pe_9_14_done),
        .go(pe_9_14_go),
        .left(pe_9_14_left),
        .out(pe_9_14_out),
        .top(pe_9_14_top)
    );
    std_reg # (
        .width(32)
    ) top_9_14 (
        .clk(top_9_14_clk),
        .done(top_9_14_done),
        .in(top_9_14_in),
        .out(top_9_14_out),
        .write_en(top_9_14_write_en)
    );
    std_reg # (
        .width(32)
    ) left_9_14 (
        .clk(left_9_14_clk),
        .done(left_9_14_done),
        .in(left_9_14_in),
        .out(left_9_14_out),
        .write_en(left_9_14_write_en)
    );
    mac_pe pe_9_15 (
        .clk(pe_9_15_clk),
        .done(pe_9_15_done),
        .go(pe_9_15_go),
        .left(pe_9_15_left),
        .out(pe_9_15_out),
        .top(pe_9_15_top)
    );
    std_reg # (
        .width(32)
    ) top_9_15 (
        .clk(top_9_15_clk),
        .done(top_9_15_done),
        .in(top_9_15_in),
        .out(top_9_15_out),
        .write_en(top_9_15_write_en)
    );
    std_reg # (
        .width(32)
    ) left_9_15 (
        .clk(left_9_15_clk),
        .done(left_9_15_done),
        .in(left_9_15_in),
        .out(left_9_15_out),
        .write_en(left_9_15_write_en)
    );
    mac_pe pe_10_0 (
        .clk(pe_10_0_clk),
        .done(pe_10_0_done),
        .go(pe_10_0_go),
        .left(pe_10_0_left),
        .out(pe_10_0_out),
        .top(pe_10_0_top)
    );
    std_reg # (
        .width(32)
    ) top_10_0 (
        .clk(top_10_0_clk),
        .done(top_10_0_done),
        .in(top_10_0_in),
        .out(top_10_0_out),
        .write_en(top_10_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_10_0 (
        .clk(left_10_0_clk),
        .done(left_10_0_done),
        .in(left_10_0_in),
        .out(left_10_0_out),
        .write_en(left_10_0_write_en)
    );
    mac_pe pe_10_1 (
        .clk(pe_10_1_clk),
        .done(pe_10_1_done),
        .go(pe_10_1_go),
        .left(pe_10_1_left),
        .out(pe_10_1_out),
        .top(pe_10_1_top)
    );
    std_reg # (
        .width(32)
    ) top_10_1 (
        .clk(top_10_1_clk),
        .done(top_10_1_done),
        .in(top_10_1_in),
        .out(top_10_1_out),
        .write_en(top_10_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_10_1 (
        .clk(left_10_1_clk),
        .done(left_10_1_done),
        .in(left_10_1_in),
        .out(left_10_1_out),
        .write_en(left_10_1_write_en)
    );
    mac_pe pe_10_2 (
        .clk(pe_10_2_clk),
        .done(pe_10_2_done),
        .go(pe_10_2_go),
        .left(pe_10_2_left),
        .out(pe_10_2_out),
        .top(pe_10_2_top)
    );
    std_reg # (
        .width(32)
    ) top_10_2 (
        .clk(top_10_2_clk),
        .done(top_10_2_done),
        .in(top_10_2_in),
        .out(top_10_2_out),
        .write_en(top_10_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_10_2 (
        .clk(left_10_2_clk),
        .done(left_10_2_done),
        .in(left_10_2_in),
        .out(left_10_2_out),
        .write_en(left_10_2_write_en)
    );
    mac_pe pe_10_3 (
        .clk(pe_10_3_clk),
        .done(pe_10_3_done),
        .go(pe_10_3_go),
        .left(pe_10_3_left),
        .out(pe_10_3_out),
        .top(pe_10_3_top)
    );
    std_reg # (
        .width(32)
    ) top_10_3 (
        .clk(top_10_3_clk),
        .done(top_10_3_done),
        .in(top_10_3_in),
        .out(top_10_3_out),
        .write_en(top_10_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_10_3 (
        .clk(left_10_3_clk),
        .done(left_10_3_done),
        .in(left_10_3_in),
        .out(left_10_3_out),
        .write_en(left_10_3_write_en)
    );
    mac_pe pe_10_4 (
        .clk(pe_10_4_clk),
        .done(pe_10_4_done),
        .go(pe_10_4_go),
        .left(pe_10_4_left),
        .out(pe_10_4_out),
        .top(pe_10_4_top)
    );
    std_reg # (
        .width(32)
    ) top_10_4 (
        .clk(top_10_4_clk),
        .done(top_10_4_done),
        .in(top_10_4_in),
        .out(top_10_4_out),
        .write_en(top_10_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_10_4 (
        .clk(left_10_4_clk),
        .done(left_10_4_done),
        .in(left_10_4_in),
        .out(left_10_4_out),
        .write_en(left_10_4_write_en)
    );
    mac_pe pe_10_5 (
        .clk(pe_10_5_clk),
        .done(pe_10_5_done),
        .go(pe_10_5_go),
        .left(pe_10_5_left),
        .out(pe_10_5_out),
        .top(pe_10_5_top)
    );
    std_reg # (
        .width(32)
    ) top_10_5 (
        .clk(top_10_5_clk),
        .done(top_10_5_done),
        .in(top_10_5_in),
        .out(top_10_5_out),
        .write_en(top_10_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_10_5 (
        .clk(left_10_5_clk),
        .done(left_10_5_done),
        .in(left_10_5_in),
        .out(left_10_5_out),
        .write_en(left_10_5_write_en)
    );
    mac_pe pe_10_6 (
        .clk(pe_10_6_clk),
        .done(pe_10_6_done),
        .go(pe_10_6_go),
        .left(pe_10_6_left),
        .out(pe_10_6_out),
        .top(pe_10_6_top)
    );
    std_reg # (
        .width(32)
    ) top_10_6 (
        .clk(top_10_6_clk),
        .done(top_10_6_done),
        .in(top_10_6_in),
        .out(top_10_6_out),
        .write_en(top_10_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_10_6 (
        .clk(left_10_6_clk),
        .done(left_10_6_done),
        .in(left_10_6_in),
        .out(left_10_6_out),
        .write_en(left_10_6_write_en)
    );
    mac_pe pe_10_7 (
        .clk(pe_10_7_clk),
        .done(pe_10_7_done),
        .go(pe_10_7_go),
        .left(pe_10_7_left),
        .out(pe_10_7_out),
        .top(pe_10_7_top)
    );
    std_reg # (
        .width(32)
    ) top_10_7 (
        .clk(top_10_7_clk),
        .done(top_10_7_done),
        .in(top_10_7_in),
        .out(top_10_7_out),
        .write_en(top_10_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_10_7 (
        .clk(left_10_7_clk),
        .done(left_10_7_done),
        .in(left_10_7_in),
        .out(left_10_7_out),
        .write_en(left_10_7_write_en)
    );
    mac_pe pe_10_8 (
        .clk(pe_10_8_clk),
        .done(pe_10_8_done),
        .go(pe_10_8_go),
        .left(pe_10_8_left),
        .out(pe_10_8_out),
        .top(pe_10_8_top)
    );
    std_reg # (
        .width(32)
    ) top_10_8 (
        .clk(top_10_8_clk),
        .done(top_10_8_done),
        .in(top_10_8_in),
        .out(top_10_8_out),
        .write_en(top_10_8_write_en)
    );
    std_reg # (
        .width(32)
    ) left_10_8 (
        .clk(left_10_8_clk),
        .done(left_10_8_done),
        .in(left_10_8_in),
        .out(left_10_8_out),
        .write_en(left_10_8_write_en)
    );
    mac_pe pe_10_9 (
        .clk(pe_10_9_clk),
        .done(pe_10_9_done),
        .go(pe_10_9_go),
        .left(pe_10_9_left),
        .out(pe_10_9_out),
        .top(pe_10_9_top)
    );
    std_reg # (
        .width(32)
    ) top_10_9 (
        .clk(top_10_9_clk),
        .done(top_10_9_done),
        .in(top_10_9_in),
        .out(top_10_9_out),
        .write_en(top_10_9_write_en)
    );
    std_reg # (
        .width(32)
    ) left_10_9 (
        .clk(left_10_9_clk),
        .done(left_10_9_done),
        .in(left_10_9_in),
        .out(left_10_9_out),
        .write_en(left_10_9_write_en)
    );
    mac_pe pe_10_10 (
        .clk(pe_10_10_clk),
        .done(pe_10_10_done),
        .go(pe_10_10_go),
        .left(pe_10_10_left),
        .out(pe_10_10_out),
        .top(pe_10_10_top)
    );
    std_reg # (
        .width(32)
    ) top_10_10 (
        .clk(top_10_10_clk),
        .done(top_10_10_done),
        .in(top_10_10_in),
        .out(top_10_10_out),
        .write_en(top_10_10_write_en)
    );
    std_reg # (
        .width(32)
    ) left_10_10 (
        .clk(left_10_10_clk),
        .done(left_10_10_done),
        .in(left_10_10_in),
        .out(left_10_10_out),
        .write_en(left_10_10_write_en)
    );
    mac_pe pe_10_11 (
        .clk(pe_10_11_clk),
        .done(pe_10_11_done),
        .go(pe_10_11_go),
        .left(pe_10_11_left),
        .out(pe_10_11_out),
        .top(pe_10_11_top)
    );
    std_reg # (
        .width(32)
    ) top_10_11 (
        .clk(top_10_11_clk),
        .done(top_10_11_done),
        .in(top_10_11_in),
        .out(top_10_11_out),
        .write_en(top_10_11_write_en)
    );
    std_reg # (
        .width(32)
    ) left_10_11 (
        .clk(left_10_11_clk),
        .done(left_10_11_done),
        .in(left_10_11_in),
        .out(left_10_11_out),
        .write_en(left_10_11_write_en)
    );
    mac_pe pe_10_12 (
        .clk(pe_10_12_clk),
        .done(pe_10_12_done),
        .go(pe_10_12_go),
        .left(pe_10_12_left),
        .out(pe_10_12_out),
        .top(pe_10_12_top)
    );
    std_reg # (
        .width(32)
    ) top_10_12 (
        .clk(top_10_12_clk),
        .done(top_10_12_done),
        .in(top_10_12_in),
        .out(top_10_12_out),
        .write_en(top_10_12_write_en)
    );
    std_reg # (
        .width(32)
    ) left_10_12 (
        .clk(left_10_12_clk),
        .done(left_10_12_done),
        .in(left_10_12_in),
        .out(left_10_12_out),
        .write_en(left_10_12_write_en)
    );
    mac_pe pe_10_13 (
        .clk(pe_10_13_clk),
        .done(pe_10_13_done),
        .go(pe_10_13_go),
        .left(pe_10_13_left),
        .out(pe_10_13_out),
        .top(pe_10_13_top)
    );
    std_reg # (
        .width(32)
    ) top_10_13 (
        .clk(top_10_13_clk),
        .done(top_10_13_done),
        .in(top_10_13_in),
        .out(top_10_13_out),
        .write_en(top_10_13_write_en)
    );
    std_reg # (
        .width(32)
    ) left_10_13 (
        .clk(left_10_13_clk),
        .done(left_10_13_done),
        .in(left_10_13_in),
        .out(left_10_13_out),
        .write_en(left_10_13_write_en)
    );
    mac_pe pe_10_14 (
        .clk(pe_10_14_clk),
        .done(pe_10_14_done),
        .go(pe_10_14_go),
        .left(pe_10_14_left),
        .out(pe_10_14_out),
        .top(pe_10_14_top)
    );
    std_reg # (
        .width(32)
    ) top_10_14 (
        .clk(top_10_14_clk),
        .done(top_10_14_done),
        .in(top_10_14_in),
        .out(top_10_14_out),
        .write_en(top_10_14_write_en)
    );
    std_reg # (
        .width(32)
    ) left_10_14 (
        .clk(left_10_14_clk),
        .done(left_10_14_done),
        .in(left_10_14_in),
        .out(left_10_14_out),
        .write_en(left_10_14_write_en)
    );
    mac_pe pe_10_15 (
        .clk(pe_10_15_clk),
        .done(pe_10_15_done),
        .go(pe_10_15_go),
        .left(pe_10_15_left),
        .out(pe_10_15_out),
        .top(pe_10_15_top)
    );
    std_reg # (
        .width(32)
    ) top_10_15 (
        .clk(top_10_15_clk),
        .done(top_10_15_done),
        .in(top_10_15_in),
        .out(top_10_15_out),
        .write_en(top_10_15_write_en)
    );
    std_reg # (
        .width(32)
    ) left_10_15 (
        .clk(left_10_15_clk),
        .done(left_10_15_done),
        .in(left_10_15_in),
        .out(left_10_15_out),
        .write_en(left_10_15_write_en)
    );
    mac_pe pe_11_0 (
        .clk(pe_11_0_clk),
        .done(pe_11_0_done),
        .go(pe_11_0_go),
        .left(pe_11_0_left),
        .out(pe_11_0_out),
        .top(pe_11_0_top)
    );
    std_reg # (
        .width(32)
    ) top_11_0 (
        .clk(top_11_0_clk),
        .done(top_11_0_done),
        .in(top_11_0_in),
        .out(top_11_0_out),
        .write_en(top_11_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_11_0 (
        .clk(left_11_0_clk),
        .done(left_11_0_done),
        .in(left_11_0_in),
        .out(left_11_0_out),
        .write_en(left_11_0_write_en)
    );
    mac_pe pe_11_1 (
        .clk(pe_11_1_clk),
        .done(pe_11_1_done),
        .go(pe_11_1_go),
        .left(pe_11_1_left),
        .out(pe_11_1_out),
        .top(pe_11_1_top)
    );
    std_reg # (
        .width(32)
    ) top_11_1 (
        .clk(top_11_1_clk),
        .done(top_11_1_done),
        .in(top_11_1_in),
        .out(top_11_1_out),
        .write_en(top_11_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_11_1 (
        .clk(left_11_1_clk),
        .done(left_11_1_done),
        .in(left_11_1_in),
        .out(left_11_1_out),
        .write_en(left_11_1_write_en)
    );
    mac_pe pe_11_2 (
        .clk(pe_11_2_clk),
        .done(pe_11_2_done),
        .go(pe_11_2_go),
        .left(pe_11_2_left),
        .out(pe_11_2_out),
        .top(pe_11_2_top)
    );
    std_reg # (
        .width(32)
    ) top_11_2 (
        .clk(top_11_2_clk),
        .done(top_11_2_done),
        .in(top_11_2_in),
        .out(top_11_2_out),
        .write_en(top_11_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_11_2 (
        .clk(left_11_2_clk),
        .done(left_11_2_done),
        .in(left_11_2_in),
        .out(left_11_2_out),
        .write_en(left_11_2_write_en)
    );
    mac_pe pe_11_3 (
        .clk(pe_11_3_clk),
        .done(pe_11_3_done),
        .go(pe_11_3_go),
        .left(pe_11_3_left),
        .out(pe_11_3_out),
        .top(pe_11_3_top)
    );
    std_reg # (
        .width(32)
    ) top_11_3 (
        .clk(top_11_3_clk),
        .done(top_11_3_done),
        .in(top_11_3_in),
        .out(top_11_3_out),
        .write_en(top_11_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_11_3 (
        .clk(left_11_3_clk),
        .done(left_11_3_done),
        .in(left_11_3_in),
        .out(left_11_3_out),
        .write_en(left_11_3_write_en)
    );
    mac_pe pe_11_4 (
        .clk(pe_11_4_clk),
        .done(pe_11_4_done),
        .go(pe_11_4_go),
        .left(pe_11_4_left),
        .out(pe_11_4_out),
        .top(pe_11_4_top)
    );
    std_reg # (
        .width(32)
    ) top_11_4 (
        .clk(top_11_4_clk),
        .done(top_11_4_done),
        .in(top_11_4_in),
        .out(top_11_4_out),
        .write_en(top_11_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_11_4 (
        .clk(left_11_4_clk),
        .done(left_11_4_done),
        .in(left_11_4_in),
        .out(left_11_4_out),
        .write_en(left_11_4_write_en)
    );
    mac_pe pe_11_5 (
        .clk(pe_11_5_clk),
        .done(pe_11_5_done),
        .go(pe_11_5_go),
        .left(pe_11_5_left),
        .out(pe_11_5_out),
        .top(pe_11_5_top)
    );
    std_reg # (
        .width(32)
    ) top_11_5 (
        .clk(top_11_5_clk),
        .done(top_11_5_done),
        .in(top_11_5_in),
        .out(top_11_5_out),
        .write_en(top_11_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_11_5 (
        .clk(left_11_5_clk),
        .done(left_11_5_done),
        .in(left_11_5_in),
        .out(left_11_5_out),
        .write_en(left_11_5_write_en)
    );
    mac_pe pe_11_6 (
        .clk(pe_11_6_clk),
        .done(pe_11_6_done),
        .go(pe_11_6_go),
        .left(pe_11_6_left),
        .out(pe_11_6_out),
        .top(pe_11_6_top)
    );
    std_reg # (
        .width(32)
    ) top_11_6 (
        .clk(top_11_6_clk),
        .done(top_11_6_done),
        .in(top_11_6_in),
        .out(top_11_6_out),
        .write_en(top_11_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_11_6 (
        .clk(left_11_6_clk),
        .done(left_11_6_done),
        .in(left_11_6_in),
        .out(left_11_6_out),
        .write_en(left_11_6_write_en)
    );
    mac_pe pe_11_7 (
        .clk(pe_11_7_clk),
        .done(pe_11_7_done),
        .go(pe_11_7_go),
        .left(pe_11_7_left),
        .out(pe_11_7_out),
        .top(pe_11_7_top)
    );
    std_reg # (
        .width(32)
    ) top_11_7 (
        .clk(top_11_7_clk),
        .done(top_11_7_done),
        .in(top_11_7_in),
        .out(top_11_7_out),
        .write_en(top_11_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_11_7 (
        .clk(left_11_7_clk),
        .done(left_11_7_done),
        .in(left_11_7_in),
        .out(left_11_7_out),
        .write_en(left_11_7_write_en)
    );
    mac_pe pe_11_8 (
        .clk(pe_11_8_clk),
        .done(pe_11_8_done),
        .go(pe_11_8_go),
        .left(pe_11_8_left),
        .out(pe_11_8_out),
        .top(pe_11_8_top)
    );
    std_reg # (
        .width(32)
    ) top_11_8 (
        .clk(top_11_8_clk),
        .done(top_11_8_done),
        .in(top_11_8_in),
        .out(top_11_8_out),
        .write_en(top_11_8_write_en)
    );
    std_reg # (
        .width(32)
    ) left_11_8 (
        .clk(left_11_8_clk),
        .done(left_11_8_done),
        .in(left_11_8_in),
        .out(left_11_8_out),
        .write_en(left_11_8_write_en)
    );
    mac_pe pe_11_9 (
        .clk(pe_11_9_clk),
        .done(pe_11_9_done),
        .go(pe_11_9_go),
        .left(pe_11_9_left),
        .out(pe_11_9_out),
        .top(pe_11_9_top)
    );
    std_reg # (
        .width(32)
    ) top_11_9 (
        .clk(top_11_9_clk),
        .done(top_11_9_done),
        .in(top_11_9_in),
        .out(top_11_9_out),
        .write_en(top_11_9_write_en)
    );
    std_reg # (
        .width(32)
    ) left_11_9 (
        .clk(left_11_9_clk),
        .done(left_11_9_done),
        .in(left_11_9_in),
        .out(left_11_9_out),
        .write_en(left_11_9_write_en)
    );
    mac_pe pe_11_10 (
        .clk(pe_11_10_clk),
        .done(pe_11_10_done),
        .go(pe_11_10_go),
        .left(pe_11_10_left),
        .out(pe_11_10_out),
        .top(pe_11_10_top)
    );
    std_reg # (
        .width(32)
    ) top_11_10 (
        .clk(top_11_10_clk),
        .done(top_11_10_done),
        .in(top_11_10_in),
        .out(top_11_10_out),
        .write_en(top_11_10_write_en)
    );
    std_reg # (
        .width(32)
    ) left_11_10 (
        .clk(left_11_10_clk),
        .done(left_11_10_done),
        .in(left_11_10_in),
        .out(left_11_10_out),
        .write_en(left_11_10_write_en)
    );
    mac_pe pe_11_11 (
        .clk(pe_11_11_clk),
        .done(pe_11_11_done),
        .go(pe_11_11_go),
        .left(pe_11_11_left),
        .out(pe_11_11_out),
        .top(pe_11_11_top)
    );
    std_reg # (
        .width(32)
    ) top_11_11 (
        .clk(top_11_11_clk),
        .done(top_11_11_done),
        .in(top_11_11_in),
        .out(top_11_11_out),
        .write_en(top_11_11_write_en)
    );
    std_reg # (
        .width(32)
    ) left_11_11 (
        .clk(left_11_11_clk),
        .done(left_11_11_done),
        .in(left_11_11_in),
        .out(left_11_11_out),
        .write_en(left_11_11_write_en)
    );
    mac_pe pe_11_12 (
        .clk(pe_11_12_clk),
        .done(pe_11_12_done),
        .go(pe_11_12_go),
        .left(pe_11_12_left),
        .out(pe_11_12_out),
        .top(pe_11_12_top)
    );
    std_reg # (
        .width(32)
    ) top_11_12 (
        .clk(top_11_12_clk),
        .done(top_11_12_done),
        .in(top_11_12_in),
        .out(top_11_12_out),
        .write_en(top_11_12_write_en)
    );
    std_reg # (
        .width(32)
    ) left_11_12 (
        .clk(left_11_12_clk),
        .done(left_11_12_done),
        .in(left_11_12_in),
        .out(left_11_12_out),
        .write_en(left_11_12_write_en)
    );
    mac_pe pe_11_13 (
        .clk(pe_11_13_clk),
        .done(pe_11_13_done),
        .go(pe_11_13_go),
        .left(pe_11_13_left),
        .out(pe_11_13_out),
        .top(pe_11_13_top)
    );
    std_reg # (
        .width(32)
    ) top_11_13 (
        .clk(top_11_13_clk),
        .done(top_11_13_done),
        .in(top_11_13_in),
        .out(top_11_13_out),
        .write_en(top_11_13_write_en)
    );
    std_reg # (
        .width(32)
    ) left_11_13 (
        .clk(left_11_13_clk),
        .done(left_11_13_done),
        .in(left_11_13_in),
        .out(left_11_13_out),
        .write_en(left_11_13_write_en)
    );
    mac_pe pe_11_14 (
        .clk(pe_11_14_clk),
        .done(pe_11_14_done),
        .go(pe_11_14_go),
        .left(pe_11_14_left),
        .out(pe_11_14_out),
        .top(pe_11_14_top)
    );
    std_reg # (
        .width(32)
    ) top_11_14 (
        .clk(top_11_14_clk),
        .done(top_11_14_done),
        .in(top_11_14_in),
        .out(top_11_14_out),
        .write_en(top_11_14_write_en)
    );
    std_reg # (
        .width(32)
    ) left_11_14 (
        .clk(left_11_14_clk),
        .done(left_11_14_done),
        .in(left_11_14_in),
        .out(left_11_14_out),
        .write_en(left_11_14_write_en)
    );
    mac_pe pe_11_15 (
        .clk(pe_11_15_clk),
        .done(pe_11_15_done),
        .go(pe_11_15_go),
        .left(pe_11_15_left),
        .out(pe_11_15_out),
        .top(pe_11_15_top)
    );
    std_reg # (
        .width(32)
    ) top_11_15 (
        .clk(top_11_15_clk),
        .done(top_11_15_done),
        .in(top_11_15_in),
        .out(top_11_15_out),
        .write_en(top_11_15_write_en)
    );
    std_reg # (
        .width(32)
    ) left_11_15 (
        .clk(left_11_15_clk),
        .done(left_11_15_done),
        .in(left_11_15_in),
        .out(left_11_15_out),
        .write_en(left_11_15_write_en)
    );
    mac_pe pe_12_0 (
        .clk(pe_12_0_clk),
        .done(pe_12_0_done),
        .go(pe_12_0_go),
        .left(pe_12_0_left),
        .out(pe_12_0_out),
        .top(pe_12_0_top)
    );
    std_reg # (
        .width(32)
    ) top_12_0 (
        .clk(top_12_0_clk),
        .done(top_12_0_done),
        .in(top_12_0_in),
        .out(top_12_0_out),
        .write_en(top_12_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_12_0 (
        .clk(left_12_0_clk),
        .done(left_12_0_done),
        .in(left_12_0_in),
        .out(left_12_0_out),
        .write_en(left_12_0_write_en)
    );
    mac_pe pe_12_1 (
        .clk(pe_12_1_clk),
        .done(pe_12_1_done),
        .go(pe_12_1_go),
        .left(pe_12_1_left),
        .out(pe_12_1_out),
        .top(pe_12_1_top)
    );
    std_reg # (
        .width(32)
    ) top_12_1 (
        .clk(top_12_1_clk),
        .done(top_12_1_done),
        .in(top_12_1_in),
        .out(top_12_1_out),
        .write_en(top_12_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_12_1 (
        .clk(left_12_1_clk),
        .done(left_12_1_done),
        .in(left_12_1_in),
        .out(left_12_1_out),
        .write_en(left_12_1_write_en)
    );
    mac_pe pe_12_2 (
        .clk(pe_12_2_clk),
        .done(pe_12_2_done),
        .go(pe_12_2_go),
        .left(pe_12_2_left),
        .out(pe_12_2_out),
        .top(pe_12_2_top)
    );
    std_reg # (
        .width(32)
    ) top_12_2 (
        .clk(top_12_2_clk),
        .done(top_12_2_done),
        .in(top_12_2_in),
        .out(top_12_2_out),
        .write_en(top_12_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_12_2 (
        .clk(left_12_2_clk),
        .done(left_12_2_done),
        .in(left_12_2_in),
        .out(left_12_2_out),
        .write_en(left_12_2_write_en)
    );
    mac_pe pe_12_3 (
        .clk(pe_12_3_clk),
        .done(pe_12_3_done),
        .go(pe_12_3_go),
        .left(pe_12_3_left),
        .out(pe_12_3_out),
        .top(pe_12_3_top)
    );
    std_reg # (
        .width(32)
    ) top_12_3 (
        .clk(top_12_3_clk),
        .done(top_12_3_done),
        .in(top_12_3_in),
        .out(top_12_3_out),
        .write_en(top_12_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_12_3 (
        .clk(left_12_3_clk),
        .done(left_12_3_done),
        .in(left_12_3_in),
        .out(left_12_3_out),
        .write_en(left_12_3_write_en)
    );
    mac_pe pe_12_4 (
        .clk(pe_12_4_clk),
        .done(pe_12_4_done),
        .go(pe_12_4_go),
        .left(pe_12_4_left),
        .out(pe_12_4_out),
        .top(pe_12_4_top)
    );
    std_reg # (
        .width(32)
    ) top_12_4 (
        .clk(top_12_4_clk),
        .done(top_12_4_done),
        .in(top_12_4_in),
        .out(top_12_4_out),
        .write_en(top_12_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_12_4 (
        .clk(left_12_4_clk),
        .done(left_12_4_done),
        .in(left_12_4_in),
        .out(left_12_4_out),
        .write_en(left_12_4_write_en)
    );
    mac_pe pe_12_5 (
        .clk(pe_12_5_clk),
        .done(pe_12_5_done),
        .go(pe_12_5_go),
        .left(pe_12_5_left),
        .out(pe_12_5_out),
        .top(pe_12_5_top)
    );
    std_reg # (
        .width(32)
    ) top_12_5 (
        .clk(top_12_5_clk),
        .done(top_12_5_done),
        .in(top_12_5_in),
        .out(top_12_5_out),
        .write_en(top_12_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_12_5 (
        .clk(left_12_5_clk),
        .done(left_12_5_done),
        .in(left_12_5_in),
        .out(left_12_5_out),
        .write_en(left_12_5_write_en)
    );
    mac_pe pe_12_6 (
        .clk(pe_12_6_clk),
        .done(pe_12_6_done),
        .go(pe_12_6_go),
        .left(pe_12_6_left),
        .out(pe_12_6_out),
        .top(pe_12_6_top)
    );
    std_reg # (
        .width(32)
    ) top_12_6 (
        .clk(top_12_6_clk),
        .done(top_12_6_done),
        .in(top_12_6_in),
        .out(top_12_6_out),
        .write_en(top_12_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_12_6 (
        .clk(left_12_6_clk),
        .done(left_12_6_done),
        .in(left_12_6_in),
        .out(left_12_6_out),
        .write_en(left_12_6_write_en)
    );
    mac_pe pe_12_7 (
        .clk(pe_12_7_clk),
        .done(pe_12_7_done),
        .go(pe_12_7_go),
        .left(pe_12_7_left),
        .out(pe_12_7_out),
        .top(pe_12_7_top)
    );
    std_reg # (
        .width(32)
    ) top_12_7 (
        .clk(top_12_7_clk),
        .done(top_12_7_done),
        .in(top_12_7_in),
        .out(top_12_7_out),
        .write_en(top_12_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_12_7 (
        .clk(left_12_7_clk),
        .done(left_12_7_done),
        .in(left_12_7_in),
        .out(left_12_7_out),
        .write_en(left_12_7_write_en)
    );
    mac_pe pe_12_8 (
        .clk(pe_12_8_clk),
        .done(pe_12_8_done),
        .go(pe_12_8_go),
        .left(pe_12_8_left),
        .out(pe_12_8_out),
        .top(pe_12_8_top)
    );
    std_reg # (
        .width(32)
    ) top_12_8 (
        .clk(top_12_8_clk),
        .done(top_12_8_done),
        .in(top_12_8_in),
        .out(top_12_8_out),
        .write_en(top_12_8_write_en)
    );
    std_reg # (
        .width(32)
    ) left_12_8 (
        .clk(left_12_8_clk),
        .done(left_12_8_done),
        .in(left_12_8_in),
        .out(left_12_8_out),
        .write_en(left_12_8_write_en)
    );
    mac_pe pe_12_9 (
        .clk(pe_12_9_clk),
        .done(pe_12_9_done),
        .go(pe_12_9_go),
        .left(pe_12_9_left),
        .out(pe_12_9_out),
        .top(pe_12_9_top)
    );
    std_reg # (
        .width(32)
    ) top_12_9 (
        .clk(top_12_9_clk),
        .done(top_12_9_done),
        .in(top_12_9_in),
        .out(top_12_9_out),
        .write_en(top_12_9_write_en)
    );
    std_reg # (
        .width(32)
    ) left_12_9 (
        .clk(left_12_9_clk),
        .done(left_12_9_done),
        .in(left_12_9_in),
        .out(left_12_9_out),
        .write_en(left_12_9_write_en)
    );
    mac_pe pe_12_10 (
        .clk(pe_12_10_clk),
        .done(pe_12_10_done),
        .go(pe_12_10_go),
        .left(pe_12_10_left),
        .out(pe_12_10_out),
        .top(pe_12_10_top)
    );
    std_reg # (
        .width(32)
    ) top_12_10 (
        .clk(top_12_10_clk),
        .done(top_12_10_done),
        .in(top_12_10_in),
        .out(top_12_10_out),
        .write_en(top_12_10_write_en)
    );
    std_reg # (
        .width(32)
    ) left_12_10 (
        .clk(left_12_10_clk),
        .done(left_12_10_done),
        .in(left_12_10_in),
        .out(left_12_10_out),
        .write_en(left_12_10_write_en)
    );
    mac_pe pe_12_11 (
        .clk(pe_12_11_clk),
        .done(pe_12_11_done),
        .go(pe_12_11_go),
        .left(pe_12_11_left),
        .out(pe_12_11_out),
        .top(pe_12_11_top)
    );
    std_reg # (
        .width(32)
    ) top_12_11 (
        .clk(top_12_11_clk),
        .done(top_12_11_done),
        .in(top_12_11_in),
        .out(top_12_11_out),
        .write_en(top_12_11_write_en)
    );
    std_reg # (
        .width(32)
    ) left_12_11 (
        .clk(left_12_11_clk),
        .done(left_12_11_done),
        .in(left_12_11_in),
        .out(left_12_11_out),
        .write_en(left_12_11_write_en)
    );
    mac_pe pe_12_12 (
        .clk(pe_12_12_clk),
        .done(pe_12_12_done),
        .go(pe_12_12_go),
        .left(pe_12_12_left),
        .out(pe_12_12_out),
        .top(pe_12_12_top)
    );
    std_reg # (
        .width(32)
    ) top_12_12 (
        .clk(top_12_12_clk),
        .done(top_12_12_done),
        .in(top_12_12_in),
        .out(top_12_12_out),
        .write_en(top_12_12_write_en)
    );
    std_reg # (
        .width(32)
    ) left_12_12 (
        .clk(left_12_12_clk),
        .done(left_12_12_done),
        .in(left_12_12_in),
        .out(left_12_12_out),
        .write_en(left_12_12_write_en)
    );
    mac_pe pe_12_13 (
        .clk(pe_12_13_clk),
        .done(pe_12_13_done),
        .go(pe_12_13_go),
        .left(pe_12_13_left),
        .out(pe_12_13_out),
        .top(pe_12_13_top)
    );
    std_reg # (
        .width(32)
    ) top_12_13 (
        .clk(top_12_13_clk),
        .done(top_12_13_done),
        .in(top_12_13_in),
        .out(top_12_13_out),
        .write_en(top_12_13_write_en)
    );
    std_reg # (
        .width(32)
    ) left_12_13 (
        .clk(left_12_13_clk),
        .done(left_12_13_done),
        .in(left_12_13_in),
        .out(left_12_13_out),
        .write_en(left_12_13_write_en)
    );
    mac_pe pe_12_14 (
        .clk(pe_12_14_clk),
        .done(pe_12_14_done),
        .go(pe_12_14_go),
        .left(pe_12_14_left),
        .out(pe_12_14_out),
        .top(pe_12_14_top)
    );
    std_reg # (
        .width(32)
    ) top_12_14 (
        .clk(top_12_14_clk),
        .done(top_12_14_done),
        .in(top_12_14_in),
        .out(top_12_14_out),
        .write_en(top_12_14_write_en)
    );
    std_reg # (
        .width(32)
    ) left_12_14 (
        .clk(left_12_14_clk),
        .done(left_12_14_done),
        .in(left_12_14_in),
        .out(left_12_14_out),
        .write_en(left_12_14_write_en)
    );
    mac_pe pe_12_15 (
        .clk(pe_12_15_clk),
        .done(pe_12_15_done),
        .go(pe_12_15_go),
        .left(pe_12_15_left),
        .out(pe_12_15_out),
        .top(pe_12_15_top)
    );
    std_reg # (
        .width(32)
    ) top_12_15 (
        .clk(top_12_15_clk),
        .done(top_12_15_done),
        .in(top_12_15_in),
        .out(top_12_15_out),
        .write_en(top_12_15_write_en)
    );
    std_reg # (
        .width(32)
    ) left_12_15 (
        .clk(left_12_15_clk),
        .done(left_12_15_done),
        .in(left_12_15_in),
        .out(left_12_15_out),
        .write_en(left_12_15_write_en)
    );
    mac_pe pe_13_0 (
        .clk(pe_13_0_clk),
        .done(pe_13_0_done),
        .go(pe_13_0_go),
        .left(pe_13_0_left),
        .out(pe_13_0_out),
        .top(pe_13_0_top)
    );
    std_reg # (
        .width(32)
    ) top_13_0 (
        .clk(top_13_0_clk),
        .done(top_13_0_done),
        .in(top_13_0_in),
        .out(top_13_0_out),
        .write_en(top_13_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_13_0 (
        .clk(left_13_0_clk),
        .done(left_13_0_done),
        .in(left_13_0_in),
        .out(left_13_0_out),
        .write_en(left_13_0_write_en)
    );
    mac_pe pe_13_1 (
        .clk(pe_13_1_clk),
        .done(pe_13_1_done),
        .go(pe_13_1_go),
        .left(pe_13_1_left),
        .out(pe_13_1_out),
        .top(pe_13_1_top)
    );
    std_reg # (
        .width(32)
    ) top_13_1 (
        .clk(top_13_1_clk),
        .done(top_13_1_done),
        .in(top_13_1_in),
        .out(top_13_1_out),
        .write_en(top_13_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_13_1 (
        .clk(left_13_1_clk),
        .done(left_13_1_done),
        .in(left_13_1_in),
        .out(left_13_1_out),
        .write_en(left_13_1_write_en)
    );
    mac_pe pe_13_2 (
        .clk(pe_13_2_clk),
        .done(pe_13_2_done),
        .go(pe_13_2_go),
        .left(pe_13_2_left),
        .out(pe_13_2_out),
        .top(pe_13_2_top)
    );
    std_reg # (
        .width(32)
    ) top_13_2 (
        .clk(top_13_2_clk),
        .done(top_13_2_done),
        .in(top_13_2_in),
        .out(top_13_2_out),
        .write_en(top_13_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_13_2 (
        .clk(left_13_2_clk),
        .done(left_13_2_done),
        .in(left_13_2_in),
        .out(left_13_2_out),
        .write_en(left_13_2_write_en)
    );
    mac_pe pe_13_3 (
        .clk(pe_13_3_clk),
        .done(pe_13_3_done),
        .go(pe_13_3_go),
        .left(pe_13_3_left),
        .out(pe_13_3_out),
        .top(pe_13_3_top)
    );
    std_reg # (
        .width(32)
    ) top_13_3 (
        .clk(top_13_3_clk),
        .done(top_13_3_done),
        .in(top_13_3_in),
        .out(top_13_3_out),
        .write_en(top_13_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_13_3 (
        .clk(left_13_3_clk),
        .done(left_13_3_done),
        .in(left_13_3_in),
        .out(left_13_3_out),
        .write_en(left_13_3_write_en)
    );
    mac_pe pe_13_4 (
        .clk(pe_13_4_clk),
        .done(pe_13_4_done),
        .go(pe_13_4_go),
        .left(pe_13_4_left),
        .out(pe_13_4_out),
        .top(pe_13_4_top)
    );
    std_reg # (
        .width(32)
    ) top_13_4 (
        .clk(top_13_4_clk),
        .done(top_13_4_done),
        .in(top_13_4_in),
        .out(top_13_4_out),
        .write_en(top_13_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_13_4 (
        .clk(left_13_4_clk),
        .done(left_13_4_done),
        .in(left_13_4_in),
        .out(left_13_4_out),
        .write_en(left_13_4_write_en)
    );
    mac_pe pe_13_5 (
        .clk(pe_13_5_clk),
        .done(pe_13_5_done),
        .go(pe_13_5_go),
        .left(pe_13_5_left),
        .out(pe_13_5_out),
        .top(pe_13_5_top)
    );
    std_reg # (
        .width(32)
    ) top_13_5 (
        .clk(top_13_5_clk),
        .done(top_13_5_done),
        .in(top_13_5_in),
        .out(top_13_5_out),
        .write_en(top_13_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_13_5 (
        .clk(left_13_5_clk),
        .done(left_13_5_done),
        .in(left_13_5_in),
        .out(left_13_5_out),
        .write_en(left_13_5_write_en)
    );
    mac_pe pe_13_6 (
        .clk(pe_13_6_clk),
        .done(pe_13_6_done),
        .go(pe_13_6_go),
        .left(pe_13_6_left),
        .out(pe_13_6_out),
        .top(pe_13_6_top)
    );
    std_reg # (
        .width(32)
    ) top_13_6 (
        .clk(top_13_6_clk),
        .done(top_13_6_done),
        .in(top_13_6_in),
        .out(top_13_6_out),
        .write_en(top_13_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_13_6 (
        .clk(left_13_6_clk),
        .done(left_13_6_done),
        .in(left_13_6_in),
        .out(left_13_6_out),
        .write_en(left_13_6_write_en)
    );
    mac_pe pe_13_7 (
        .clk(pe_13_7_clk),
        .done(pe_13_7_done),
        .go(pe_13_7_go),
        .left(pe_13_7_left),
        .out(pe_13_7_out),
        .top(pe_13_7_top)
    );
    std_reg # (
        .width(32)
    ) top_13_7 (
        .clk(top_13_7_clk),
        .done(top_13_7_done),
        .in(top_13_7_in),
        .out(top_13_7_out),
        .write_en(top_13_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_13_7 (
        .clk(left_13_7_clk),
        .done(left_13_7_done),
        .in(left_13_7_in),
        .out(left_13_7_out),
        .write_en(left_13_7_write_en)
    );
    mac_pe pe_13_8 (
        .clk(pe_13_8_clk),
        .done(pe_13_8_done),
        .go(pe_13_8_go),
        .left(pe_13_8_left),
        .out(pe_13_8_out),
        .top(pe_13_8_top)
    );
    std_reg # (
        .width(32)
    ) top_13_8 (
        .clk(top_13_8_clk),
        .done(top_13_8_done),
        .in(top_13_8_in),
        .out(top_13_8_out),
        .write_en(top_13_8_write_en)
    );
    std_reg # (
        .width(32)
    ) left_13_8 (
        .clk(left_13_8_clk),
        .done(left_13_8_done),
        .in(left_13_8_in),
        .out(left_13_8_out),
        .write_en(left_13_8_write_en)
    );
    mac_pe pe_13_9 (
        .clk(pe_13_9_clk),
        .done(pe_13_9_done),
        .go(pe_13_9_go),
        .left(pe_13_9_left),
        .out(pe_13_9_out),
        .top(pe_13_9_top)
    );
    std_reg # (
        .width(32)
    ) top_13_9 (
        .clk(top_13_9_clk),
        .done(top_13_9_done),
        .in(top_13_9_in),
        .out(top_13_9_out),
        .write_en(top_13_9_write_en)
    );
    std_reg # (
        .width(32)
    ) left_13_9 (
        .clk(left_13_9_clk),
        .done(left_13_9_done),
        .in(left_13_9_in),
        .out(left_13_9_out),
        .write_en(left_13_9_write_en)
    );
    mac_pe pe_13_10 (
        .clk(pe_13_10_clk),
        .done(pe_13_10_done),
        .go(pe_13_10_go),
        .left(pe_13_10_left),
        .out(pe_13_10_out),
        .top(pe_13_10_top)
    );
    std_reg # (
        .width(32)
    ) top_13_10 (
        .clk(top_13_10_clk),
        .done(top_13_10_done),
        .in(top_13_10_in),
        .out(top_13_10_out),
        .write_en(top_13_10_write_en)
    );
    std_reg # (
        .width(32)
    ) left_13_10 (
        .clk(left_13_10_clk),
        .done(left_13_10_done),
        .in(left_13_10_in),
        .out(left_13_10_out),
        .write_en(left_13_10_write_en)
    );
    mac_pe pe_13_11 (
        .clk(pe_13_11_clk),
        .done(pe_13_11_done),
        .go(pe_13_11_go),
        .left(pe_13_11_left),
        .out(pe_13_11_out),
        .top(pe_13_11_top)
    );
    std_reg # (
        .width(32)
    ) top_13_11 (
        .clk(top_13_11_clk),
        .done(top_13_11_done),
        .in(top_13_11_in),
        .out(top_13_11_out),
        .write_en(top_13_11_write_en)
    );
    std_reg # (
        .width(32)
    ) left_13_11 (
        .clk(left_13_11_clk),
        .done(left_13_11_done),
        .in(left_13_11_in),
        .out(left_13_11_out),
        .write_en(left_13_11_write_en)
    );
    mac_pe pe_13_12 (
        .clk(pe_13_12_clk),
        .done(pe_13_12_done),
        .go(pe_13_12_go),
        .left(pe_13_12_left),
        .out(pe_13_12_out),
        .top(pe_13_12_top)
    );
    std_reg # (
        .width(32)
    ) top_13_12 (
        .clk(top_13_12_clk),
        .done(top_13_12_done),
        .in(top_13_12_in),
        .out(top_13_12_out),
        .write_en(top_13_12_write_en)
    );
    std_reg # (
        .width(32)
    ) left_13_12 (
        .clk(left_13_12_clk),
        .done(left_13_12_done),
        .in(left_13_12_in),
        .out(left_13_12_out),
        .write_en(left_13_12_write_en)
    );
    mac_pe pe_13_13 (
        .clk(pe_13_13_clk),
        .done(pe_13_13_done),
        .go(pe_13_13_go),
        .left(pe_13_13_left),
        .out(pe_13_13_out),
        .top(pe_13_13_top)
    );
    std_reg # (
        .width(32)
    ) top_13_13 (
        .clk(top_13_13_clk),
        .done(top_13_13_done),
        .in(top_13_13_in),
        .out(top_13_13_out),
        .write_en(top_13_13_write_en)
    );
    std_reg # (
        .width(32)
    ) left_13_13 (
        .clk(left_13_13_clk),
        .done(left_13_13_done),
        .in(left_13_13_in),
        .out(left_13_13_out),
        .write_en(left_13_13_write_en)
    );
    mac_pe pe_13_14 (
        .clk(pe_13_14_clk),
        .done(pe_13_14_done),
        .go(pe_13_14_go),
        .left(pe_13_14_left),
        .out(pe_13_14_out),
        .top(pe_13_14_top)
    );
    std_reg # (
        .width(32)
    ) top_13_14 (
        .clk(top_13_14_clk),
        .done(top_13_14_done),
        .in(top_13_14_in),
        .out(top_13_14_out),
        .write_en(top_13_14_write_en)
    );
    std_reg # (
        .width(32)
    ) left_13_14 (
        .clk(left_13_14_clk),
        .done(left_13_14_done),
        .in(left_13_14_in),
        .out(left_13_14_out),
        .write_en(left_13_14_write_en)
    );
    mac_pe pe_13_15 (
        .clk(pe_13_15_clk),
        .done(pe_13_15_done),
        .go(pe_13_15_go),
        .left(pe_13_15_left),
        .out(pe_13_15_out),
        .top(pe_13_15_top)
    );
    std_reg # (
        .width(32)
    ) top_13_15 (
        .clk(top_13_15_clk),
        .done(top_13_15_done),
        .in(top_13_15_in),
        .out(top_13_15_out),
        .write_en(top_13_15_write_en)
    );
    std_reg # (
        .width(32)
    ) left_13_15 (
        .clk(left_13_15_clk),
        .done(left_13_15_done),
        .in(left_13_15_in),
        .out(left_13_15_out),
        .write_en(left_13_15_write_en)
    );
    mac_pe pe_14_0 (
        .clk(pe_14_0_clk),
        .done(pe_14_0_done),
        .go(pe_14_0_go),
        .left(pe_14_0_left),
        .out(pe_14_0_out),
        .top(pe_14_0_top)
    );
    std_reg # (
        .width(32)
    ) top_14_0 (
        .clk(top_14_0_clk),
        .done(top_14_0_done),
        .in(top_14_0_in),
        .out(top_14_0_out),
        .write_en(top_14_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_14_0 (
        .clk(left_14_0_clk),
        .done(left_14_0_done),
        .in(left_14_0_in),
        .out(left_14_0_out),
        .write_en(left_14_0_write_en)
    );
    mac_pe pe_14_1 (
        .clk(pe_14_1_clk),
        .done(pe_14_1_done),
        .go(pe_14_1_go),
        .left(pe_14_1_left),
        .out(pe_14_1_out),
        .top(pe_14_1_top)
    );
    std_reg # (
        .width(32)
    ) top_14_1 (
        .clk(top_14_1_clk),
        .done(top_14_1_done),
        .in(top_14_1_in),
        .out(top_14_1_out),
        .write_en(top_14_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_14_1 (
        .clk(left_14_1_clk),
        .done(left_14_1_done),
        .in(left_14_1_in),
        .out(left_14_1_out),
        .write_en(left_14_1_write_en)
    );
    mac_pe pe_14_2 (
        .clk(pe_14_2_clk),
        .done(pe_14_2_done),
        .go(pe_14_2_go),
        .left(pe_14_2_left),
        .out(pe_14_2_out),
        .top(pe_14_2_top)
    );
    std_reg # (
        .width(32)
    ) top_14_2 (
        .clk(top_14_2_clk),
        .done(top_14_2_done),
        .in(top_14_2_in),
        .out(top_14_2_out),
        .write_en(top_14_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_14_2 (
        .clk(left_14_2_clk),
        .done(left_14_2_done),
        .in(left_14_2_in),
        .out(left_14_2_out),
        .write_en(left_14_2_write_en)
    );
    mac_pe pe_14_3 (
        .clk(pe_14_3_clk),
        .done(pe_14_3_done),
        .go(pe_14_3_go),
        .left(pe_14_3_left),
        .out(pe_14_3_out),
        .top(pe_14_3_top)
    );
    std_reg # (
        .width(32)
    ) top_14_3 (
        .clk(top_14_3_clk),
        .done(top_14_3_done),
        .in(top_14_3_in),
        .out(top_14_3_out),
        .write_en(top_14_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_14_3 (
        .clk(left_14_3_clk),
        .done(left_14_3_done),
        .in(left_14_3_in),
        .out(left_14_3_out),
        .write_en(left_14_3_write_en)
    );
    mac_pe pe_14_4 (
        .clk(pe_14_4_clk),
        .done(pe_14_4_done),
        .go(pe_14_4_go),
        .left(pe_14_4_left),
        .out(pe_14_4_out),
        .top(pe_14_4_top)
    );
    std_reg # (
        .width(32)
    ) top_14_4 (
        .clk(top_14_4_clk),
        .done(top_14_4_done),
        .in(top_14_4_in),
        .out(top_14_4_out),
        .write_en(top_14_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_14_4 (
        .clk(left_14_4_clk),
        .done(left_14_4_done),
        .in(left_14_4_in),
        .out(left_14_4_out),
        .write_en(left_14_4_write_en)
    );
    mac_pe pe_14_5 (
        .clk(pe_14_5_clk),
        .done(pe_14_5_done),
        .go(pe_14_5_go),
        .left(pe_14_5_left),
        .out(pe_14_5_out),
        .top(pe_14_5_top)
    );
    std_reg # (
        .width(32)
    ) top_14_5 (
        .clk(top_14_5_clk),
        .done(top_14_5_done),
        .in(top_14_5_in),
        .out(top_14_5_out),
        .write_en(top_14_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_14_5 (
        .clk(left_14_5_clk),
        .done(left_14_5_done),
        .in(left_14_5_in),
        .out(left_14_5_out),
        .write_en(left_14_5_write_en)
    );
    mac_pe pe_14_6 (
        .clk(pe_14_6_clk),
        .done(pe_14_6_done),
        .go(pe_14_6_go),
        .left(pe_14_6_left),
        .out(pe_14_6_out),
        .top(pe_14_6_top)
    );
    std_reg # (
        .width(32)
    ) top_14_6 (
        .clk(top_14_6_clk),
        .done(top_14_6_done),
        .in(top_14_6_in),
        .out(top_14_6_out),
        .write_en(top_14_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_14_6 (
        .clk(left_14_6_clk),
        .done(left_14_6_done),
        .in(left_14_6_in),
        .out(left_14_6_out),
        .write_en(left_14_6_write_en)
    );
    mac_pe pe_14_7 (
        .clk(pe_14_7_clk),
        .done(pe_14_7_done),
        .go(pe_14_7_go),
        .left(pe_14_7_left),
        .out(pe_14_7_out),
        .top(pe_14_7_top)
    );
    std_reg # (
        .width(32)
    ) top_14_7 (
        .clk(top_14_7_clk),
        .done(top_14_7_done),
        .in(top_14_7_in),
        .out(top_14_7_out),
        .write_en(top_14_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_14_7 (
        .clk(left_14_7_clk),
        .done(left_14_7_done),
        .in(left_14_7_in),
        .out(left_14_7_out),
        .write_en(left_14_7_write_en)
    );
    mac_pe pe_14_8 (
        .clk(pe_14_8_clk),
        .done(pe_14_8_done),
        .go(pe_14_8_go),
        .left(pe_14_8_left),
        .out(pe_14_8_out),
        .top(pe_14_8_top)
    );
    std_reg # (
        .width(32)
    ) top_14_8 (
        .clk(top_14_8_clk),
        .done(top_14_8_done),
        .in(top_14_8_in),
        .out(top_14_8_out),
        .write_en(top_14_8_write_en)
    );
    std_reg # (
        .width(32)
    ) left_14_8 (
        .clk(left_14_8_clk),
        .done(left_14_8_done),
        .in(left_14_8_in),
        .out(left_14_8_out),
        .write_en(left_14_8_write_en)
    );
    mac_pe pe_14_9 (
        .clk(pe_14_9_clk),
        .done(pe_14_9_done),
        .go(pe_14_9_go),
        .left(pe_14_9_left),
        .out(pe_14_9_out),
        .top(pe_14_9_top)
    );
    std_reg # (
        .width(32)
    ) top_14_9 (
        .clk(top_14_9_clk),
        .done(top_14_9_done),
        .in(top_14_9_in),
        .out(top_14_9_out),
        .write_en(top_14_9_write_en)
    );
    std_reg # (
        .width(32)
    ) left_14_9 (
        .clk(left_14_9_clk),
        .done(left_14_9_done),
        .in(left_14_9_in),
        .out(left_14_9_out),
        .write_en(left_14_9_write_en)
    );
    mac_pe pe_14_10 (
        .clk(pe_14_10_clk),
        .done(pe_14_10_done),
        .go(pe_14_10_go),
        .left(pe_14_10_left),
        .out(pe_14_10_out),
        .top(pe_14_10_top)
    );
    std_reg # (
        .width(32)
    ) top_14_10 (
        .clk(top_14_10_clk),
        .done(top_14_10_done),
        .in(top_14_10_in),
        .out(top_14_10_out),
        .write_en(top_14_10_write_en)
    );
    std_reg # (
        .width(32)
    ) left_14_10 (
        .clk(left_14_10_clk),
        .done(left_14_10_done),
        .in(left_14_10_in),
        .out(left_14_10_out),
        .write_en(left_14_10_write_en)
    );
    mac_pe pe_14_11 (
        .clk(pe_14_11_clk),
        .done(pe_14_11_done),
        .go(pe_14_11_go),
        .left(pe_14_11_left),
        .out(pe_14_11_out),
        .top(pe_14_11_top)
    );
    std_reg # (
        .width(32)
    ) top_14_11 (
        .clk(top_14_11_clk),
        .done(top_14_11_done),
        .in(top_14_11_in),
        .out(top_14_11_out),
        .write_en(top_14_11_write_en)
    );
    std_reg # (
        .width(32)
    ) left_14_11 (
        .clk(left_14_11_clk),
        .done(left_14_11_done),
        .in(left_14_11_in),
        .out(left_14_11_out),
        .write_en(left_14_11_write_en)
    );
    mac_pe pe_14_12 (
        .clk(pe_14_12_clk),
        .done(pe_14_12_done),
        .go(pe_14_12_go),
        .left(pe_14_12_left),
        .out(pe_14_12_out),
        .top(pe_14_12_top)
    );
    std_reg # (
        .width(32)
    ) top_14_12 (
        .clk(top_14_12_clk),
        .done(top_14_12_done),
        .in(top_14_12_in),
        .out(top_14_12_out),
        .write_en(top_14_12_write_en)
    );
    std_reg # (
        .width(32)
    ) left_14_12 (
        .clk(left_14_12_clk),
        .done(left_14_12_done),
        .in(left_14_12_in),
        .out(left_14_12_out),
        .write_en(left_14_12_write_en)
    );
    mac_pe pe_14_13 (
        .clk(pe_14_13_clk),
        .done(pe_14_13_done),
        .go(pe_14_13_go),
        .left(pe_14_13_left),
        .out(pe_14_13_out),
        .top(pe_14_13_top)
    );
    std_reg # (
        .width(32)
    ) top_14_13 (
        .clk(top_14_13_clk),
        .done(top_14_13_done),
        .in(top_14_13_in),
        .out(top_14_13_out),
        .write_en(top_14_13_write_en)
    );
    std_reg # (
        .width(32)
    ) left_14_13 (
        .clk(left_14_13_clk),
        .done(left_14_13_done),
        .in(left_14_13_in),
        .out(left_14_13_out),
        .write_en(left_14_13_write_en)
    );
    mac_pe pe_14_14 (
        .clk(pe_14_14_clk),
        .done(pe_14_14_done),
        .go(pe_14_14_go),
        .left(pe_14_14_left),
        .out(pe_14_14_out),
        .top(pe_14_14_top)
    );
    std_reg # (
        .width(32)
    ) top_14_14 (
        .clk(top_14_14_clk),
        .done(top_14_14_done),
        .in(top_14_14_in),
        .out(top_14_14_out),
        .write_en(top_14_14_write_en)
    );
    std_reg # (
        .width(32)
    ) left_14_14 (
        .clk(left_14_14_clk),
        .done(left_14_14_done),
        .in(left_14_14_in),
        .out(left_14_14_out),
        .write_en(left_14_14_write_en)
    );
    mac_pe pe_14_15 (
        .clk(pe_14_15_clk),
        .done(pe_14_15_done),
        .go(pe_14_15_go),
        .left(pe_14_15_left),
        .out(pe_14_15_out),
        .top(pe_14_15_top)
    );
    std_reg # (
        .width(32)
    ) top_14_15 (
        .clk(top_14_15_clk),
        .done(top_14_15_done),
        .in(top_14_15_in),
        .out(top_14_15_out),
        .write_en(top_14_15_write_en)
    );
    std_reg # (
        .width(32)
    ) left_14_15 (
        .clk(left_14_15_clk),
        .done(left_14_15_done),
        .in(left_14_15_in),
        .out(left_14_15_out),
        .write_en(left_14_15_write_en)
    );
    mac_pe pe_15_0 (
        .clk(pe_15_0_clk),
        .done(pe_15_0_done),
        .go(pe_15_0_go),
        .left(pe_15_0_left),
        .out(pe_15_0_out),
        .top(pe_15_0_top)
    );
    std_reg # (
        .width(32)
    ) top_15_0 (
        .clk(top_15_0_clk),
        .done(top_15_0_done),
        .in(top_15_0_in),
        .out(top_15_0_out),
        .write_en(top_15_0_write_en)
    );
    std_reg # (
        .width(32)
    ) left_15_0 (
        .clk(left_15_0_clk),
        .done(left_15_0_done),
        .in(left_15_0_in),
        .out(left_15_0_out),
        .write_en(left_15_0_write_en)
    );
    mac_pe pe_15_1 (
        .clk(pe_15_1_clk),
        .done(pe_15_1_done),
        .go(pe_15_1_go),
        .left(pe_15_1_left),
        .out(pe_15_1_out),
        .top(pe_15_1_top)
    );
    std_reg # (
        .width(32)
    ) top_15_1 (
        .clk(top_15_1_clk),
        .done(top_15_1_done),
        .in(top_15_1_in),
        .out(top_15_1_out),
        .write_en(top_15_1_write_en)
    );
    std_reg # (
        .width(32)
    ) left_15_1 (
        .clk(left_15_1_clk),
        .done(left_15_1_done),
        .in(left_15_1_in),
        .out(left_15_1_out),
        .write_en(left_15_1_write_en)
    );
    mac_pe pe_15_2 (
        .clk(pe_15_2_clk),
        .done(pe_15_2_done),
        .go(pe_15_2_go),
        .left(pe_15_2_left),
        .out(pe_15_2_out),
        .top(pe_15_2_top)
    );
    std_reg # (
        .width(32)
    ) top_15_2 (
        .clk(top_15_2_clk),
        .done(top_15_2_done),
        .in(top_15_2_in),
        .out(top_15_2_out),
        .write_en(top_15_2_write_en)
    );
    std_reg # (
        .width(32)
    ) left_15_2 (
        .clk(left_15_2_clk),
        .done(left_15_2_done),
        .in(left_15_2_in),
        .out(left_15_2_out),
        .write_en(left_15_2_write_en)
    );
    mac_pe pe_15_3 (
        .clk(pe_15_3_clk),
        .done(pe_15_3_done),
        .go(pe_15_3_go),
        .left(pe_15_3_left),
        .out(pe_15_3_out),
        .top(pe_15_3_top)
    );
    std_reg # (
        .width(32)
    ) top_15_3 (
        .clk(top_15_3_clk),
        .done(top_15_3_done),
        .in(top_15_3_in),
        .out(top_15_3_out),
        .write_en(top_15_3_write_en)
    );
    std_reg # (
        .width(32)
    ) left_15_3 (
        .clk(left_15_3_clk),
        .done(left_15_3_done),
        .in(left_15_3_in),
        .out(left_15_3_out),
        .write_en(left_15_3_write_en)
    );
    mac_pe pe_15_4 (
        .clk(pe_15_4_clk),
        .done(pe_15_4_done),
        .go(pe_15_4_go),
        .left(pe_15_4_left),
        .out(pe_15_4_out),
        .top(pe_15_4_top)
    );
    std_reg # (
        .width(32)
    ) top_15_4 (
        .clk(top_15_4_clk),
        .done(top_15_4_done),
        .in(top_15_4_in),
        .out(top_15_4_out),
        .write_en(top_15_4_write_en)
    );
    std_reg # (
        .width(32)
    ) left_15_4 (
        .clk(left_15_4_clk),
        .done(left_15_4_done),
        .in(left_15_4_in),
        .out(left_15_4_out),
        .write_en(left_15_4_write_en)
    );
    mac_pe pe_15_5 (
        .clk(pe_15_5_clk),
        .done(pe_15_5_done),
        .go(pe_15_5_go),
        .left(pe_15_5_left),
        .out(pe_15_5_out),
        .top(pe_15_5_top)
    );
    std_reg # (
        .width(32)
    ) top_15_5 (
        .clk(top_15_5_clk),
        .done(top_15_5_done),
        .in(top_15_5_in),
        .out(top_15_5_out),
        .write_en(top_15_5_write_en)
    );
    std_reg # (
        .width(32)
    ) left_15_5 (
        .clk(left_15_5_clk),
        .done(left_15_5_done),
        .in(left_15_5_in),
        .out(left_15_5_out),
        .write_en(left_15_5_write_en)
    );
    mac_pe pe_15_6 (
        .clk(pe_15_6_clk),
        .done(pe_15_6_done),
        .go(pe_15_6_go),
        .left(pe_15_6_left),
        .out(pe_15_6_out),
        .top(pe_15_6_top)
    );
    std_reg # (
        .width(32)
    ) top_15_6 (
        .clk(top_15_6_clk),
        .done(top_15_6_done),
        .in(top_15_6_in),
        .out(top_15_6_out),
        .write_en(top_15_6_write_en)
    );
    std_reg # (
        .width(32)
    ) left_15_6 (
        .clk(left_15_6_clk),
        .done(left_15_6_done),
        .in(left_15_6_in),
        .out(left_15_6_out),
        .write_en(left_15_6_write_en)
    );
    mac_pe pe_15_7 (
        .clk(pe_15_7_clk),
        .done(pe_15_7_done),
        .go(pe_15_7_go),
        .left(pe_15_7_left),
        .out(pe_15_7_out),
        .top(pe_15_7_top)
    );
    std_reg # (
        .width(32)
    ) top_15_7 (
        .clk(top_15_7_clk),
        .done(top_15_7_done),
        .in(top_15_7_in),
        .out(top_15_7_out),
        .write_en(top_15_7_write_en)
    );
    std_reg # (
        .width(32)
    ) left_15_7 (
        .clk(left_15_7_clk),
        .done(left_15_7_done),
        .in(left_15_7_in),
        .out(left_15_7_out),
        .write_en(left_15_7_write_en)
    );
    mac_pe pe_15_8 (
        .clk(pe_15_8_clk),
        .done(pe_15_8_done),
        .go(pe_15_8_go),
        .left(pe_15_8_left),
        .out(pe_15_8_out),
        .top(pe_15_8_top)
    );
    std_reg # (
        .width(32)
    ) top_15_8 (
        .clk(top_15_8_clk),
        .done(top_15_8_done),
        .in(top_15_8_in),
        .out(top_15_8_out),
        .write_en(top_15_8_write_en)
    );
    std_reg # (
        .width(32)
    ) left_15_8 (
        .clk(left_15_8_clk),
        .done(left_15_8_done),
        .in(left_15_8_in),
        .out(left_15_8_out),
        .write_en(left_15_8_write_en)
    );
    mac_pe pe_15_9 (
        .clk(pe_15_9_clk),
        .done(pe_15_9_done),
        .go(pe_15_9_go),
        .left(pe_15_9_left),
        .out(pe_15_9_out),
        .top(pe_15_9_top)
    );
    std_reg # (
        .width(32)
    ) top_15_9 (
        .clk(top_15_9_clk),
        .done(top_15_9_done),
        .in(top_15_9_in),
        .out(top_15_9_out),
        .write_en(top_15_9_write_en)
    );
    std_reg # (
        .width(32)
    ) left_15_9 (
        .clk(left_15_9_clk),
        .done(left_15_9_done),
        .in(left_15_9_in),
        .out(left_15_9_out),
        .write_en(left_15_9_write_en)
    );
    mac_pe pe_15_10 (
        .clk(pe_15_10_clk),
        .done(pe_15_10_done),
        .go(pe_15_10_go),
        .left(pe_15_10_left),
        .out(pe_15_10_out),
        .top(pe_15_10_top)
    );
    std_reg # (
        .width(32)
    ) top_15_10 (
        .clk(top_15_10_clk),
        .done(top_15_10_done),
        .in(top_15_10_in),
        .out(top_15_10_out),
        .write_en(top_15_10_write_en)
    );
    std_reg # (
        .width(32)
    ) left_15_10 (
        .clk(left_15_10_clk),
        .done(left_15_10_done),
        .in(left_15_10_in),
        .out(left_15_10_out),
        .write_en(left_15_10_write_en)
    );
    mac_pe pe_15_11 (
        .clk(pe_15_11_clk),
        .done(pe_15_11_done),
        .go(pe_15_11_go),
        .left(pe_15_11_left),
        .out(pe_15_11_out),
        .top(pe_15_11_top)
    );
    std_reg # (
        .width(32)
    ) top_15_11 (
        .clk(top_15_11_clk),
        .done(top_15_11_done),
        .in(top_15_11_in),
        .out(top_15_11_out),
        .write_en(top_15_11_write_en)
    );
    std_reg # (
        .width(32)
    ) left_15_11 (
        .clk(left_15_11_clk),
        .done(left_15_11_done),
        .in(left_15_11_in),
        .out(left_15_11_out),
        .write_en(left_15_11_write_en)
    );
    mac_pe pe_15_12 (
        .clk(pe_15_12_clk),
        .done(pe_15_12_done),
        .go(pe_15_12_go),
        .left(pe_15_12_left),
        .out(pe_15_12_out),
        .top(pe_15_12_top)
    );
    std_reg # (
        .width(32)
    ) top_15_12 (
        .clk(top_15_12_clk),
        .done(top_15_12_done),
        .in(top_15_12_in),
        .out(top_15_12_out),
        .write_en(top_15_12_write_en)
    );
    std_reg # (
        .width(32)
    ) left_15_12 (
        .clk(left_15_12_clk),
        .done(left_15_12_done),
        .in(left_15_12_in),
        .out(left_15_12_out),
        .write_en(left_15_12_write_en)
    );
    mac_pe pe_15_13 (
        .clk(pe_15_13_clk),
        .done(pe_15_13_done),
        .go(pe_15_13_go),
        .left(pe_15_13_left),
        .out(pe_15_13_out),
        .top(pe_15_13_top)
    );
    std_reg # (
        .width(32)
    ) top_15_13 (
        .clk(top_15_13_clk),
        .done(top_15_13_done),
        .in(top_15_13_in),
        .out(top_15_13_out),
        .write_en(top_15_13_write_en)
    );
    std_reg # (
        .width(32)
    ) left_15_13 (
        .clk(left_15_13_clk),
        .done(left_15_13_done),
        .in(left_15_13_in),
        .out(left_15_13_out),
        .write_en(left_15_13_write_en)
    );
    mac_pe pe_15_14 (
        .clk(pe_15_14_clk),
        .done(pe_15_14_done),
        .go(pe_15_14_go),
        .left(pe_15_14_left),
        .out(pe_15_14_out),
        .top(pe_15_14_top)
    );
    std_reg # (
        .width(32)
    ) top_15_14 (
        .clk(top_15_14_clk),
        .done(top_15_14_done),
        .in(top_15_14_in),
        .out(top_15_14_out),
        .write_en(top_15_14_write_en)
    );
    std_reg # (
        .width(32)
    ) left_15_14 (
        .clk(left_15_14_clk),
        .done(left_15_14_done),
        .in(left_15_14_in),
        .out(left_15_14_out),
        .write_en(left_15_14_write_en)
    );
    mac_pe pe_15_15 (
        .clk(pe_15_15_clk),
        .done(pe_15_15_done),
        .go(pe_15_15_go),
        .left(pe_15_15_left),
        .out(pe_15_15_out),
        .top(pe_15_15_top)
    );
    std_reg # (
        .width(32)
    ) top_15_15 (
        .clk(top_15_15_clk),
        .done(top_15_15_done),
        .in(top_15_15_in),
        .out(top_15_15_out),
        .write_en(top_15_15_write_en)
    );
    std_reg # (
        .width(32)
    ) left_15_15 (
        .clk(left_15_15_clk),
        .done(left_15_15_done),
        .in(left_15_15_in),
        .out(left_15_15_out),
        .write_en(left_15_15_write_en)
    );
    std_reg # (
        .width(1)
    ) fsm (
        .clk(fsm_clk),
        .done(fsm_done),
        .in(fsm_in),
        .out(fsm_out),
        .write_en(fsm_write_en)
    );
    std_add # (
        .width(1)
    ) incr (
        .left(incr_left),
        .out(incr_out),
        .right(incr_right)
    );
    std_reg # (
        .width(1)
    ) fsm0 (
        .clk(fsm0_clk),
        .done(fsm0_done),
        .in(fsm0_in),
        .out(fsm0_out),
        .write_en(fsm0_write_en)
    );
    std_add # (
        .width(1)
    ) incr0 (
        .left(incr0_left),
        .out(incr0_out),
        .right(incr0_right)
    );
    std_reg # (
        .width(1)
    ) fsm1 (
        .clk(fsm1_clk),
        .done(fsm1_done),
        .in(fsm1_in),
        .out(fsm1_out),
        .write_en(fsm1_write_en)
    );
    std_add # (
        .width(1)
    ) incr1 (
        .left(incr1_left),
        .out(incr1_out),
        .right(incr1_right)
    );
    std_reg # (
        .width(3)
    ) fsm2 (
        .clk(fsm2_clk),
        .done(fsm2_done),
        .in(fsm2_in),
        .out(fsm2_out),
        .write_en(fsm2_write_en)
    );
    std_add # (
        .width(3)
    ) incr2 (
        .left(incr2_left),
        .out(incr2_out),
        .right(incr2_right)
    );
    std_reg # (
        .width(1)
    ) fsm3 (
        .clk(fsm3_clk),
        .done(fsm3_done),
        .in(fsm3_in),
        .out(fsm3_out),
        .write_en(fsm3_write_en)
    );
    std_add # (
        .width(1)
    ) incr3 (
        .left(incr3_left),
        .out(incr3_out),
        .right(incr3_right)
    );
    std_reg # (
        .width(3)
    ) fsm4 (
        .clk(fsm4_clk),
        .done(fsm4_done),
        .in(fsm4_in),
        .out(fsm4_out),
        .write_en(fsm4_write_en)
    );
    std_add # (
        .width(3)
    ) incr4 (
        .left(incr4_left),
        .out(incr4_out),
        .right(incr4_right)
    );
    std_reg # (
        .width(1)
    ) fsm5 (
        .clk(fsm5_clk),
        .done(fsm5_done),
        .in(fsm5_in),
        .out(fsm5_out),
        .write_en(fsm5_write_en)
    );
    std_add # (
        .width(1)
    ) incr5 (
        .left(incr5_left),
        .out(incr5_out),
        .right(incr5_right)
    );
    std_reg # (
        .width(3)
    ) fsm6 (
        .clk(fsm6_clk),
        .done(fsm6_done),
        .in(fsm6_in),
        .out(fsm6_out),
        .write_en(fsm6_write_en)
    );
    std_add # (
        .width(3)
    ) incr6 (
        .left(incr6_left),
        .out(incr6_out),
        .right(incr6_right)
    );
    std_reg # (
        .width(1)
    ) fsm7 (
        .clk(fsm7_clk),
        .done(fsm7_done),
        .in(fsm7_in),
        .out(fsm7_out),
        .write_en(fsm7_write_en)
    );
    std_add # (
        .width(1)
    ) incr7 (
        .left(incr7_left),
        .out(incr7_out),
        .right(incr7_right)
    );
    std_reg # (
        .width(3)
    ) fsm8 (
        .clk(fsm8_clk),
        .done(fsm8_done),
        .in(fsm8_in),
        .out(fsm8_out),
        .write_en(fsm8_write_en)
    );
    std_add # (
        .width(3)
    ) incr8 (
        .left(incr8_left),
        .out(incr8_out),
        .right(incr8_right)
    );
    std_reg # (
        .width(1)
    ) fsm9 (
        .clk(fsm9_clk),
        .done(fsm9_done),
        .in(fsm9_in),
        .out(fsm9_out),
        .write_en(fsm9_write_en)
    );
    std_add # (
        .width(1)
    ) incr9 (
        .left(incr9_left),
        .out(incr9_out),
        .right(incr9_right)
    );
    std_reg # (
        .width(3)
    ) fsm10 (
        .clk(fsm10_clk),
        .done(fsm10_done),
        .in(fsm10_in),
        .out(fsm10_out),
        .write_en(fsm10_write_en)
    );
    std_add # (
        .width(3)
    ) incr10 (
        .left(incr10_left),
        .out(incr10_out),
        .right(incr10_right)
    );
    std_reg # (
        .width(1)
    ) fsm11 (
        .clk(fsm11_clk),
        .done(fsm11_done),
        .in(fsm11_in),
        .out(fsm11_out),
        .write_en(fsm11_write_en)
    );
    std_add # (
        .width(1)
    ) incr11 (
        .left(incr11_left),
        .out(incr11_out),
        .right(incr11_right)
    );
    std_reg # (
        .width(3)
    ) fsm12 (
        .clk(fsm12_clk),
        .done(fsm12_done),
        .in(fsm12_in),
        .out(fsm12_out),
        .write_en(fsm12_write_en)
    );
    std_add # (
        .width(3)
    ) incr12 (
        .left(incr12_left),
        .out(incr12_out),
        .right(incr12_right)
    );
    std_reg # (
        .width(1)
    ) fsm13 (
        .clk(fsm13_clk),
        .done(fsm13_done),
        .in(fsm13_in),
        .out(fsm13_out),
        .write_en(fsm13_write_en)
    );
    std_add # (
        .width(1)
    ) incr13 (
        .left(incr13_left),
        .out(incr13_out),
        .right(incr13_right)
    );
    std_reg # (
        .width(3)
    ) fsm14 (
        .clk(fsm14_clk),
        .done(fsm14_done),
        .in(fsm14_in),
        .out(fsm14_out),
        .write_en(fsm14_write_en)
    );
    std_add # (
        .width(3)
    ) incr14 (
        .left(incr14_left),
        .out(incr14_out),
        .right(incr14_right)
    );
    std_reg # (
        .width(1)
    ) fsm15 (
        .clk(fsm15_clk),
        .done(fsm15_done),
        .in(fsm15_in),
        .out(fsm15_out),
        .write_en(fsm15_write_en)
    );
    std_add # (
        .width(1)
    ) incr15 (
        .left(incr15_left),
        .out(incr15_out),
        .right(incr15_right)
    );
    std_reg # (
        .width(3)
    ) fsm16 (
        .clk(fsm16_clk),
        .done(fsm16_done),
        .in(fsm16_in),
        .out(fsm16_out),
        .write_en(fsm16_write_en)
    );
    std_add # (
        .width(3)
    ) incr16 (
        .left(incr16_left),
        .out(incr16_out),
        .right(incr16_right)
    );
    std_reg # (
        .width(1)
    ) fsm17 (
        .clk(fsm17_clk),
        .done(fsm17_done),
        .in(fsm17_in),
        .out(fsm17_out),
        .write_en(fsm17_write_en)
    );
    std_add # (
        .width(1)
    ) incr17 (
        .left(incr17_left),
        .out(incr17_out),
        .right(incr17_right)
    );
    std_reg # (
        .width(3)
    ) fsm18 (
        .clk(fsm18_clk),
        .done(fsm18_done),
        .in(fsm18_in),
        .out(fsm18_out),
        .write_en(fsm18_write_en)
    );
    std_add # (
        .width(3)
    ) incr18 (
        .left(incr18_left),
        .out(incr18_out),
        .right(incr18_right)
    );
    std_reg # (
        .width(1)
    ) fsm19 (
        .clk(fsm19_clk),
        .done(fsm19_done),
        .in(fsm19_in),
        .out(fsm19_out),
        .write_en(fsm19_write_en)
    );
    std_add # (
        .width(1)
    ) incr19 (
        .left(incr19_left),
        .out(incr19_out),
        .right(incr19_right)
    );
    std_reg # (
        .width(3)
    ) fsm20 (
        .clk(fsm20_clk),
        .done(fsm20_done),
        .in(fsm20_in),
        .out(fsm20_out),
        .write_en(fsm20_write_en)
    );
    std_add # (
        .width(3)
    ) incr20 (
        .left(incr20_left),
        .out(incr20_out),
        .right(incr20_right)
    );
    std_reg # (
        .width(1)
    ) fsm21 (
        .clk(fsm21_clk),
        .done(fsm21_done),
        .in(fsm21_in),
        .out(fsm21_out),
        .write_en(fsm21_write_en)
    );
    std_add # (
        .width(1)
    ) incr21 (
        .left(incr21_left),
        .out(incr21_out),
        .right(incr21_right)
    );
    std_reg # (
        .width(3)
    ) fsm22 (
        .clk(fsm22_clk),
        .done(fsm22_done),
        .in(fsm22_in),
        .out(fsm22_out),
        .write_en(fsm22_write_en)
    );
    std_add # (
        .width(3)
    ) incr22 (
        .left(incr22_left),
        .out(incr22_out),
        .right(incr22_right)
    );
    std_reg # (
        .width(1)
    ) fsm23 (
        .clk(fsm23_clk),
        .done(fsm23_done),
        .in(fsm23_in),
        .out(fsm23_out),
        .write_en(fsm23_write_en)
    );
    std_add # (
        .width(1)
    ) incr23 (
        .left(incr23_left),
        .out(incr23_out),
        .right(incr23_right)
    );
    std_reg # (
        .width(3)
    ) fsm24 (
        .clk(fsm24_clk),
        .done(fsm24_done),
        .in(fsm24_in),
        .out(fsm24_out),
        .write_en(fsm24_write_en)
    );
    std_add # (
        .width(3)
    ) incr24 (
        .left(incr24_left),
        .out(incr24_out),
        .right(incr24_right)
    );
    std_reg # (
        .width(1)
    ) fsm25 (
        .clk(fsm25_clk),
        .done(fsm25_done),
        .in(fsm25_in),
        .out(fsm25_out),
        .write_en(fsm25_write_en)
    );
    std_add # (
        .width(1)
    ) incr25 (
        .left(incr25_left),
        .out(incr25_out),
        .right(incr25_right)
    );
    std_reg # (
        .width(3)
    ) fsm26 (
        .clk(fsm26_clk),
        .done(fsm26_done),
        .in(fsm26_in),
        .out(fsm26_out),
        .write_en(fsm26_write_en)
    );
    std_add # (
        .width(3)
    ) incr26 (
        .left(incr26_left),
        .out(incr26_out),
        .right(incr26_right)
    );
    std_reg # (
        .width(1)
    ) fsm27 (
        .clk(fsm27_clk),
        .done(fsm27_done),
        .in(fsm27_in),
        .out(fsm27_out),
        .write_en(fsm27_write_en)
    );
    std_add # (
        .width(1)
    ) incr27 (
        .left(incr27_left),
        .out(incr27_out),
        .right(incr27_right)
    );
    std_reg # (
        .width(3)
    ) fsm28 (
        .clk(fsm28_clk),
        .done(fsm28_done),
        .in(fsm28_in),
        .out(fsm28_out),
        .write_en(fsm28_write_en)
    );
    std_add # (
        .width(3)
    ) incr28 (
        .left(incr28_left),
        .out(incr28_out),
        .right(incr28_right)
    );
    std_reg # (
        .width(1)
    ) fsm29 (
        .clk(fsm29_clk),
        .done(fsm29_done),
        .in(fsm29_in),
        .out(fsm29_out),
        .write_en(fsm29_write_en)
    );
    std_add # (
        .width(1)
    ) incr29 (
        .left(incr29_left),
        .out(incr29_out),
        .right(incr29_right)
    );
    std_reg # (
        .width(3)
    ) fsm30 (
        .clk(fsm30_clk),
        .done(fsm30_done),
        .in(fsm30_in),
        .out(fsm30_out),
        .write_en(fsm30_write_en)
    );
    std_add # (
        .width(3)
    ) incr30 (
        .left(incr30_left),
        .out(incr30_out),
        .right(incr30_right)
    );
    std_reg # (
        .width(1)
    ) fsm31 (
        .clk(fsm31_clk),
        .done(fsm31_done),
        .in(fsm31_in),
        .out(fsm31_out),
        .write_en(fsm31_write_en)
    );
    std_add # (
        .width(1)
    ) incr31 (
        .left(incr31_left),
        .out(incr31_out),
        .right(incr31_right)
    );
    std_reg # (
        .width(3)
    ) fsm32 (
        .clk(fsm32_clk),
        .done(fsm32_done),
        .in(fsm32_in),
        .out(fsm32_out),
        .write_en(fsm32_write_en)
    );
    std_add # (
        .width(3)
    ) incr32 (
        .left(incr32_left),
        .out(incr32_out),
        .right(incr32_right)
    );
    std_reg # (
        .width(1)
    ) fsm33 (
        .clk(fsm33_clk),
        .done(fsm33_done),
        .in(fsm33_in),
        .out(fsm33_out),
        .write_en(fsm33_write_en)
    );
    std_add # (
        .width(1)
    ) incr33 (
        .left(incr33_left),
        .out(incr33_out),
        .right(incr33_right)
    );
    std_reg # (
        .width(3)
    ) fsm34 (
        .clk(fsm34_clk),
        .done(fsm34_done),
        .in(fsm34_in),
        .out(fsm34_out),
        .write_en(fsm34_write_en)
    );
    std_add # (
        .width(3)
    ) incr34 (
        .left(incr34_left),
        .out(incr34_out),
        .right(incr34_right)
    );
    std_reg # (
        .width(1)
    ) fsm35 (
        .clk(fsm35_clk),
        .done(fsm35_done),
        .in(fsm35_in),
        .out(fsm35_out),
        .write_en(fsm35_write_en)
    );
    std_add # (
        .width(1)
    ) incr35 (
        .left(incr35_left),
        .out(incr35_out),
        .right(incr35_right)
    );
    std_reg # (
        .width(3)
    ) fsm36 (
        .clk(fsm36_clk),
        .done(fsm36_done),
        .in(fsm36_in),
        .out(fsm36_out),
        .write_en(fsm36_write_en)
    );
    std_add # (
        .width(3)
    ) incr36 (
        .left(incr36_left),
        .out(incr36_out),
        .right(incr36_right)
    );
    std_reg # (
        .width(1)
    ) fsm37 (
        .clk(fsm37_clk),
        .done(fsm37_done),
        .in(fsm37_in),
        .out(fsm37_out),
        .write_en(fsm37_write_en)
    );
    std_add # (
        .width(1)
    ) incr37 (
        .left(incr37_left),
        .out(incr37_out),
        .right(incr37_right)
    );
    std_reg # (
        .width(3)
    ) fsm38 (
        .clk(fsm38_clk),
        .done(fsm38_done),
        .in(fsm38_in),
        .out(fsm38_out),
        .write_en(fsm38_write_en)
    );
    std_add # (
        .width(3)
    ) incr38 (
        .left(incr38_left),
        .out(incr38_out),
        .right(incr38_right)
    );
    std_reg # (
        .width(1)
    ) fsm39 (
        .clk(fsm39_clk),
        .done(fsm39_done),
        .in(fsm39_in),
        .out(fsm39_out),
        .write_en(fsm39_write_en)
    );
    std_add # (
        .width(1)
    ) incr39 (
        .left(incr39_left),
        .out(incr39_out),
        .right(incr39_right)
    );
    std_reg # (
        .width(3)
    ) fsm40 (
        .clk(fsm40_clk),
        .done(fsm40_done),
        .in(fsm40_in),
        .out(fsm40_out),
        .write_en(fsm40_write_en)
    );
    std_add # (
        .width(3)
    ) incr40 (
        .left(incr40_left),
        .out(incr40_out),
        .right(incr40_right)
    );
    std_reg # (
        .width(1)
    ) fsm41 (
        .clk(fsm41_clk),
        .done(fsm41_done),
        .in(fsm41_in),
        .out(fsm41_out),
        .write_en(fsm41_write_en)
    );
    std_add # (
        .width(1)
    ) incr41 (
        .left(incr41_left),
        .out(incr41_out),
        .right(incr41_right)
    );
    std_reg # (
        .width(3)
    ) fsm42 (
        .clk(fsm42_clk),
        .done(fsm42_done),
        .in(fsm42_in),
        .out(fsm42_out),
        .write_en(fsm42_write_en)
    );
    std_add # (
        .width(3)
    ) incr42 (
        .left(incr42_left),
        .out(incr42_out),
        .right(incr42_right)
    );
    std_reg # (
        .width(1)
    ) fsm43 (
        .clk(fsm43_clk),
        .done(fsm43_done),
        .in(fsm43_in),
        .out(fsm43_out),
        .write_en(fsm43_write_en)
    );
    std_add # (
        .width(1)
    ) incr43 (
        .left(incr43_left),
        .out(incr43_out),
        .right(incr43_right)
    );
    std_reg # (
        .width(3)
    ) fsm44 (
        .clk(fsm44_clk),
        .done(fsm44_done),
        .in(fsm44_in),
        .out(fsm44_out),
        .write_en(fsm44_write_en)
    );
    std_add # (
        .width(3)
    ) incr44 (
        .left(incr44_left),
        .out(incr44_out),
        .right(incr44_right)
    );
    std_reg # (
        .width(1)
    ) fsm45 (
        .clk(fsm45_clk),
        .done(fsm45_done),
        .in(fsm45_in),
        .out(fsm45_out),
        .write_en(fsm45_write_en)
    );
    std_add # (
        .width(1)
    ) incr45 (
        .left(incr45_left),
        .out(incr45_out),
        .right(incr45_right)
    );
    std_reg # (
        .width(3)
    ) fsm46 (
        .clk(fsm46_clk),
        .done(fsm46_done),
        .in(fsm46_in),
        .out(fsm46_out),
        .write_en(fsm46_write_en)
    );
    std_add # (
        .width(3)
    ) incr46 (
        .left(incr46_left),
        .out(incr46_out),
        .right(incr46_right)
    );
    std_reg # (
        .width(1)
    ) fsm47 (
        .clk(fsm47_clk),
        .done(fsm47_done),
        .in(fsm47_in),
        .out(fsm47_out),
        .write_en(fsm47_write_en)
    );
    std_add # (
        .width(1)
    ) incr47 (
        .left(incr47_left),
        .out(incr47_out),
        .right(incr47_right)
    );
    std_reg # (
        .width(3)
    ) fsm48 (
        .clk(fsm48_clk),
        .done(fsm48_done),
        .in(fsm48_in),
        .out(fsm48_out),
        .write_en(fsm48_write_en)
    );
    std_add # (
        .width(3)
    ) incr48 (
        .left(incr48_left),
        .out(incr48_out),
        .right(incr48_right)
    );
    std_reg # (
        .width(1)
    ) fsm49 (
        .clk(fsm49_clk),
        .done(fsm49_done),
        .in(fsm49_in),
        .out(fsm49_out),
        .write_en(fsm49_write_en)
    );
    std_add # (
        .width(1)
    ) incr49 (
        .left(incr49_left),
        .out(incr49_out),
        .right(incr49_right)
    );
    std_reg # (
        .width(3)
    ) fsm50 (
        .clk(fsm50_clk),
        .done(fsm50_done),
        .in(fsm50_in),
        .out(fsm50_out),
        .write_en(fsm50_write_en)
    );
    std_add # (
        .width(3)
    ) incr50 (
        .left(incr50_left),
        .out(incr50_out),
        .right(incr50_right)
    );
    std_reg # (
        .width(1)
    ) fsm51 (
        .clk(fsm51_clk),
        .done(fsm51_done),
        .in(fsm51_in),
        .out(fsm51_out),
        .write_en(fsm51_write_en)
    );
    std_add # (
        .width(1)
    ) incr51 (
        .left(incr51_left),
        .out(incr51_out),
        .right(incr51_right)
    );
    std_reg # (
        .width(3)
    ) fsm52 (
        .clk(fsm52_clk),
        .done(fsm52_done),
        .in(fsm52_in),
        .out(fsm52_out),
        .write_en(fsm52_write_en)
    );
    std_add # (
        .width(3)
    ) incr52 (
        .left(incr52_left),
        .out(incr52_out),
        .right(incr52_right)
    );
    std_reg # (
        .width(1)
    ) fsm53 (
        .clk(fsm53_clk),
        .done(fsm53_done),
        .in(fsm53_in),
        .out(fsm53_out),
        .write_en(fsm53_write_en)
    );
    std_add # (
        .width(1)
    ) incr53 (
        .left(incr53_left),
        .out(incr53_out),
        .right(incr53_right)
    );
    std_reg # (
        .width(3)
    ) fsm54 (
        .clk(fsm54_clk),
        .done(fsm54_done),
        .in(fsm54_in),
        .out(fsm54_out),
        .write_en(fsm54_write_en)
    );
    std_add # (
        .width(3)
    ) incr54 (
        .left(incr54_left),
        .out(incr54_out),
        .right(incr54_right)
    );
    std_reg # (
        .width(1)
    ) fsm55 (
        .clk(fsm55_clk),
        .done(fsm55_done),
        .in(fsm55_in),
        .out(fsm55_out),
        .write_en(fsm55_write_en)
    );
    std_add # (
        .width(1)
    ) incr55 (
        .left(incr55_left),
        .out(incr55_out),
        .right(incr55_right)
    );
    std_reg # (
        .width(3)
    ) fsm56 (
        .clk(fsm56_clk),
        .done(fsm56_done),
        .in(fsm56_in),
        .out(fsm56_out),
        .write_en(fsm56_write_en)
    );
    std_add # (
        .width(3)
    ) incr56 (
        .left(incr56_left),
        .out(incr56_out),
        .right(incr56_right)
    );
    std_reg # (
        .width(1)
    ) fsm57 (
        .clk(fsm57_clk),
        .done(fsm57_done),
        .in(fsm57_in),
        .out(fsm57_out),
        .write_en(fsm57_write_en)
    );
    std_add # (
        .width(1)
    ) incr57 (
        .left(incr57_left),
        .out(incr57_out),
        .right(incr57_right)
    );
    std_reg # (
        .width(3)
    ) fsm58 (
        .clk(fsm58_clk),
        .done(fsm58_done),
        .in(fsm58_in),
        .out(fsm58_out),
        .write_en(fsm58_write_en)
    );
    std_add # (
        .width(3)
    ) incr58 (
        .left(incr58_left),
        .out(incr58_out),
        .right(incr58_right)
    );
    std_reg # (
        .width(1)
    ) fsm59 (
        .clk(fsm59_clk),
        .done(fsm59_done),
        .in(fsm59_in),
        .out(fsm59_out),
        .write_en(fsm59_write_en)
    );
    std_add # (
        .width(1)
    ) incr59 (
        .left(incr59_left),
        .out(incr59_out),
        .right(incr59_right)
    );
    std_reg # (
        .width(3)
    ) fsm60 (
        .clk(fsm60_clk),
        .done(fsm60_done),
        .in(fsm60_in),
        .out(fsm60_out),
        .write_en(fsm60_write_en)
    );
    std_add # (
        .width(3)
    ) incr60 (
        .left(incr60_left),
        .out(incr60_out),
        .right(incr60_right)
    );
    std_reg # (
        .width(1)
    ) fsm61 (
        .clk(fsm61_clk),
        .done(fsm61_done),
        .in(fsm61_in),
        .out(fsm61_out),
        .write_en(fsm61_write_en)
    );
    std_add # (
        .width(1)
    ) incr61 (
        .left(incr61_left),
        .out(incr61_out),
        .right(incr61_right)
    );
    std_reg # (
        .width(3)
    ) fsm62 (
        .clk(fsm62_clk),
        .done(fsm62_done),
        .in(fsm62_in),
        .out(fsm62_out),
        .write_en(fsm62_write_en)
    );
    std_add # (
        .width(3)
    ) incr62 (
        .left(incr62_left),
        .out(incr62_out),
        .right(incr62_right)
    );
    std_reg # (
        .width(1)
    ) fsm63 (
        .clk(fsm63_clk),
        .done(fsm63_done),
        .in(fsm63_in),
        .out(fsm63_out),
        .write_en(fsm63_write_en)
    );
    std_add # (
        .width(1)
    ) incr63 (
        .left(incr63_left),
        .out(incr63_out),
        .right(incr63_right)
    );
    std_reg # (
        .width(3)
    ) fsm64 (
        .clk(fsm64_clk),
        .done(fsm64_done),
        .in(fsm64_in),
        .out(fsm64_out),
        .write_en(fsm64_write_en)
    );
    std_add # (
        .width(3)
    ) incr64 (
        .left(incr64_left),
        .out(incr64_out),
        .right(incr64_right)
    );
    std_reg # (
        .width(1)
    ) fsm65 (
        .clk(fsm65_clk),
        .done(fsm65_done),
        .in(fsm65_in),
        .out(fsm65_out),
        .write_en(fsm65_write_en)
    );
    std_add # (
        .width(1)
    ) incr65 (
        .left(incr65_left),
        .out(incr65_out),
        .right(incr65_right)
    );
    std_reg # (
        .width(3)
    ) fsm66 (
        .clk(fsm66_clk),
        .done(fsm66_done),
        .in(fsm66_in),
        .out(fsm66_out),
        .write_en(fsm66_write_en)
    );
    std_add # (
        .width(3)
    ) incr66 (
        .left(incr66_left),
        .out(incr66_out),
        .right(incr66_right)
    );
    std_reg # (
        .width(1)
    ) fsm67 (
        .clk(fsm67_clk),
        .done(fsm67_done),
        .in(fsm67_in),
        .out(fsm67_out),
        .write_en(fsm67_write_en)
    );
    std_add # (
        .width(1)
    ) incr67 (
        .left(incr67_left),
        .out(incr67_out),
        .right(incr67_right)
    );
    std_reg # (
        .width(3)
    ) fsm68 (
        .clk(fsm68_clk),
        .done(fsm68_done),
        .in(fsm68_in),
        .out(fsm68_out),
        .write_en(fsm68_write_en)
    );
    std_add # (
        .width(3)
    ) incr68 (
        .left(incr68_left),
        .out(incr68_out),
        .right(incr68_right)
    );
    std_reg # (
        .width(1)
    ) fsm69 (
        .clk(fsm69_clk),
        .done(fsm69_done),
        .in(fsm69_in),
        .out(fsm69_out),
        .write_en(fsm69_write_en)
    );
    std_add # (
        .width(1)
    ) incr69 (
        .left(incr69_left),
        .out(incr69_out),
        .right(incr69_right)
    );
    std_reg # (
        .width(3)
    ) fsm70 (
        .clk(fsm70_clk),
        .done(fsm70_done),
        .in(fsm70_in),
        .out(fsm70_out),
        .write_en(fsm70_write_en)
    );
    std_add # (
        .width(3)
    ) incr70 (
        .left(incr70_left),
        .out(incr70_out),
        .right(incr70_right)
    );
    std_reg # (
        .width(1)
    ) fsm71 (
        .clk(fsm71_clk),
        .done(fsm71_done),
        .in(fsm71_in),
        .out(fsm71_out),
        .write_en(fsm71_write_en)
    );
    std_add # (
        .width(1)
    ) incr71 (
        .left(incr71_left),
        .out(incr71_out),
        .right(incr71_right)
    );
    std_reg # (
        .width(3)
    ) fsm72 (
        .clk(fsm72_clk),
        .done(fsm72_done),
        .in(fsm72_in),
        .out(fsm72_out),
        .write_en(fsm72_write_en)
    );
    std_add # (
        .width(3)
    ) incr72 (
        .left(incr72_left),
        .out(incr72_out),
        .right(incr72_right)
    );
    std_reg # (
        .width(1)
    ) fsm73 (
        .clk(fsm73_clk),
        .done(fsm73_done),
        .in(fsm73_in),
        .out(fsm73_out),
        .write_en(fsm73_write_en)
    );
    std_add # (
        .width(1)
    ) incr73 (
        .left(incr73_left),
        .out(incr73_out),
        .right(incr73_right)
    );
    std_reg # (
        .width(3)
    ) fsm74 (
        .clk(fsm74_clk),
        .done(fsm74_done),
        .in(fsm74_in),
        .out(fsm74_out),
        .write_en(fsm74_write_en)
    );
    std_add # (
        .width(3)
    ) incr74 (
        .left(incr74_left),
        .out(incr74_out),
        .right(incr74_right)
    );
    std_reg # (
        .width(1)
    ) fsm75 (
        .clk(fsm75_clk),
        .done(fsm75_done),
        .in(fsm75_in),
        .out(fsm75_out),
        .write_en(fsm75_write_en)
    );
    std_add # (
        .width(1)
    ) incr75 (
        .left(incr75_left),
        .out(incr75_out),
        .right(incr75_right)
    );
    std_reg # (
        .width(3)
    ) fsm76 (
        .clk(fsm76_clk),
        .done(fsm76_done),
        .in(fsm76_in),
        .out(fsm76_out),
        .write_en(fsm76_write_en)
    );
    std_add # (
        .width(3)
    ) incr76 (
        .left(incr76_left),
        .out(incr76_out),
        .right(incr76_right)
    );
    std_reg # (
        .width(1)
    ) fsm77 (
        .clk(fsm77_clk),
        .done(fsm77_done),
        .in(fsm77_in),
        .out(fsm77_out),
        .write_en(fsm77_write_en)
    );
    std_add # (
        .width(1)
    ) incr77 (
        .left(incr77_left),
        .out(incr77_out),
        .right(incr77_right)
    );
    std_reg # (
        .width(3)
    ) fsm78 (
        .clk(fsm78_clk),
        .done(fsm78_done),
        .in(fsm78_in),
        .out(fsm78_out),
        .write_en(fsm78_write_en)
    );
    std_add # (
        .width(3)
    ) incr78 (
        .left(incr78_left),
        .out(incr78_out),
        .right(incr78_right)
    );
    std_reg # (
        .width(1)
    ) fsm79 (
        .clk(fsm79_clk),
        .done(fsm79_done),
        .in(fsm79_in),
        .out(fsm79_out),
        .write_en(fsm79_write_en)
    );
    std_add # (
        .width(1)
    ) incr79 (
        .left(incr79_left),
        .out(incr79_out),
        .right(incr79_right)
    );
    std_reg # (
        .width(3)
    ) fsm80 (
        .clk(fsm80_clk),
        .done(fsm80_done),
        .in(fsm80_in),
        .out(fsm80_out),
        .write_en(fsm80_write_en)
    );
    std_add # (
        .width(3)
    ) incr80 (
        .left(incr80_left),
        .out(incr80_out),
        .right(incr80_right)
    );
    std_reg # (
        .width(1)
    ) fsm81 (
        .clk(fsm81_clk),
        .done(fsm81_done),
        .in(fsm81_in),
        .out(fsm81_out),
        .write_en(fsm81_write_en)
    );
    std_add # (
        .width(1)
    ) incr81 (
        .left(incr81_left),
        .out(incr81_out),
        .right(incr81_right)
    );
    std_reg # (
        .width(3)
    ) fsm82 (
        .clk(fsm82_clk),
        .done(fsm82_done),
        .in(fsm82_in),
        .out(fsm82_out),
        .write_en(fsm82_write_en)
    );
    std_add # (
        .width(3)
    ) incr82 (
        .left(incr82_left),
        .out(incr82_out),
        .right(incr82_right)
    );
    std_reg # (
        .width(1)
    ) fsm83 (
        .clk(fsm83_clk),
        .done(fsm83_done),
        .in(fsm83_in),
        .out(fsm83_out),
        .write_en(fsm83_write_en)
    );
    std_add # (
        .width(1)
    ) incr83 (
        .left(incr83_left),
        .out(incr83_out),
        .right(incr83_right)
    );
    std_reg # (
        .width(3)
    ) fsm84 (
        .clk(fsm84_clk),
        .done(fsm84_done),
        .in(fsm84_in),
        .out(fsm84_out),
        .write_en(fsm84_write_en)
    );
    std_add # (
        .width(3)
    ) incr84 (
        .left(incr84_left),
        .out(incr84_out),
        .right(incr84_right)
    );
    std_reg # (
        .width(1)
    ) fsm85 (
        .clk(fsm85_clk),
        .done(fsm85_done),
        .in(fsm85_in),
        .out(fsm85_out),
        .write_en(fsm85_write_en)
    );
    std_add # (
        .width(1)
    ) incr85 (
        .left(incr85_left),
        .out(incr85_out),
        .right(incr85_right)
    );
    std_reg # (
        .width(3)
    ) fsm86 (
        .clk(fsm86_clk),
        .done(fsm86_done),
        .in(fsm86_in),
        .out(fsm86_out),
        .write_en(fsm86_write_en)
    );
    std_add # (
        .width(3)
    ) incr86 (
        .left(incr86_left),
        .out(incr86_out),
        .right(incr86_right)
    );
    std_reg # (
        .width(1)
    ) fsm87 (
        .clk(fsm87_clk),
        .done(fsm87_done),
        .in(fsm87_in),
        .out(fsm87_out),
        .write_en(fsm87_write_en)
    );
    std_add # (
        .width(1)
    ) incr87 (
        .left(incr87_left),
        .out(incr87_out),
        .right(incr87_right)
    );
    std_reg # (
        .width(3)
    ) fsm88 (
        .clk(fsm88_clk),
        .done(fsm88_done),
        .in(fsm88_in),
        .out(fsm88_out),
        .write_en(fsm88_write_en)
    );
    std_add # (
        .width(3)
    ) incr88 (
        .left(incr88_left),
        .out(incr88_out),
        .right(incr88_right)
    );
    std_reg # (
        .width(1)
    ) fsm89 (
        .clk(fsm89_clk),
        .done(fsm89_done),
        .in(fsm89_in),
        .out(fsm89_out),
        .write_en(fsm89_write_en)
    );
    std_add # (
        .width(1)
    ) incr89 (
        .left(incr89_left),
        .out(incr89_out),
        .right(incr89_right)
    );
    std_reg # (
        .width(3)
    ) fsm90 (
        .clk(fsm90_clk),
        .done(fsm90_done),
        .in(fsm90_in),
        .out(fsm90_out),
        .write_en(fsm90_write_en)
    );
    std_add # (
        .width(3)
    ) incr90 (
        .left(incr90_left),
        .out(incr90_out),
        .right(incr90_right)
    );
    std_reg # (
        .width(1)
    ) fsm91 (
        .clk(fsm91_clk),
        .done(fsm91_done),
        .in(fsm91_in),
        .out(fsm91_out),
        .write_en(fsm91_write_en)
    );
    std_add # (
        .width(1)
    ) incr91 (
        .left(incr91_left),
        .out(incr91_out),
        .right(incr91_right)
    );
    std_reg # (
        .width(10)
    ) fsm92 (
        .clk(fsm92_clk),
        .done(fsm92_done),
        .in(fsm92_in),
        .out(fsm92_out),
        .write_en(fsm92_write_en)
    );
    std_add # (
        .width(10)
    ) incr92 (
        .left(incr92_left),
        .out(incr92_out),
        .right(incr92_right)
    );
    assign done =
     fsm92_out == 10'd534 ? 1'd1 : 1'd0;
    assign l0_addr0 =
     fsm1_out < 1'd1 & fsm92_out == 10'd2 & go | fsm3_out < 1'd1 & fsm92_out == 10'd8 & go | fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go ? l0_idx_out : 5'd0;
    assign l0_clk =
     1'b1 ? clk : 1'd0;
    assign l10_addr0 =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? l10_idx_out : 5'd0;
    assign l10_clk =
     1'b1 ? clk : 1'd0;
    assign l11_addr0 =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? l11_idx_out : 5'd0;
    assign l11_clk =
     1'b1 ? clk : 1'd0;
    assign l12_addr0 =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? l12_idx_out : 5'd0;
    assign l12_clk =
     1'b1 ? clk : 1'd0;
    assign l13_addr0 =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? l13_idx_out : 5'd0;
    assign l13_clk =
     1'b1 ? clk : 1'd0;
    assign l14_addr0 =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? l14_idx_out : 5'd0;
    assign l14_clk =
     1'b1 ? clk : 1'd0;
    assign l15_addr0 =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? l15_idx_out : 5'd0;
    assign l15_clk =
     1'b1 ? clk : 1'd0;
    assign l1_addr0 =
     fsm3_out < 1'd1 & fsm92_out == 10'd8 & go | fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go ? l1_idx_out : 5'd0;
    assign l1_clk =
     1'b1 ? clk : 1'd0;
    assign l2_addr0 =
     fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go ? l2_idx_out : 5'd0;
    assign l2_clk =
     1'b1 ? clk : 1'd0;
    assign l3_addr0 =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? l3_idx_out : 5'd0;
    assign l3_clk =
     1'b1 ? clk : 1'd0;
    assign l4_addr0 =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? l4_idx_out : 5'd0;
    assign l4_clk =
     1'b1 ? clk : 1'd0;
    assign l5_addr0 =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? l5_idx_out : 5'd0;
    assign l5_clk =
     1'b1 ? clk : 1'd0;
    assign l6_addr0 =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? l6_idx_out : 5'd0;
    assign l6_clk =
     1'b1 ? clk : 1'd0;
    assign l7_addr0 =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? l7_idx_out : 5'd0;
    assign l7_clk =
     1'b1 ? clk : 1'd0;
    assign l8_addr0 =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? l8_idx_out : 5'd0;
    assign l8_clk =
     1'b1 ? clk : 1'd0;
    assign l9_addr0 =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? l9_idx_out : 5'd0;
    assign l9_clk =
     1'b1 ? clk : 1'd0;
    assign out_mem_addr0 =
     fsm92_out == 10'd278 & go | fsm92_out == 10'd279 & go | fsm92_out == 10'd280 & go | fsm92_out == 10'd281 & go | fsm92_out == 10'd282 & go | fsm92_out == 10'd283 & go | fsm92_out == 10'd284 & go | fsm92_out == 10'd285 & go | fsm92_out == 10'd286 & go | fsm92_out == 10'd287 & go | fsm92_out == 10'd288 & go | fsm92_out == 10'd289 & go | fsm92_out == 10'd290 & go | fsm92_out == 10'd291 & go | fsm92_out == 10'd292 & go | fsm92_out == 10'd293 & go ? 5'd0 :
     fsm92_out == 10'd438 & go | fsm92_out == 10'd439 & go | fsm92_out == 10'd440 & go | fsm92_out == 10'd441 & go | fsm92_out == 10'd442 & go | fsm92_out == 10'd443 & go | fsm92_out == 10'd444 & go | fsm92_out == 10'd445 & go | fsm92_out == 10'd446 & go | fsm92_out == 10'd447 & go | fsm92_out == 10'd448 & go | fsm92_out == 10'd449 & go | fsm92_out == 10'd450 & go | fsm92_out == 10'd451 & go | fsm92_out == 10'd452 & go | fsm92_out == 10'd453 & go ? 5'd10 :
     fsm92_out == 10'd454 & go | fsm92_out == 10'd455 & go | fsm92_out == 10'd456 & go | fsm92_out == 10'd457 & go | fsm92_out == 10'd458 & go | fsm92_out == 10'd459 & go | fsm92_out == 10'd460 & go | fsm92_out == 10'd461 & go | fsm92_out == 10'd462 & go | fsm92_out == 10'd463 & go | fsm92_out == 10'd464 & go | fsm92_out == 10'd465 & go | fsm92_out == 10'd466 & go | fsm92_out == 10'd467 & go | fsm92_out == 10'd468 & go | fsm92_out == 10'd469 & go ? 5'd11 :
     fsm92_out == 10'd470 & go | fsm92_out == 10'd471 & go | fsm92_out == 10'd472 & go | fsm92_out == 10'd473 & go | fsm92_out == 10'd474 & go | fsm92_out == 10'd475 & go | fsm92_out == 10'd476 & go | fsm92_out == 10'd477 & go | fsm92_out == 10'd478 & go | fsm92_out == 10'd479 & go | fsm92_out == 10'd480 & go | fsm92_out == 10'd481 & go | fsm92_out == 10'd482 & go | fsm92_out == 10'd483 & go | fsm92_out == 10'd484 & go | fsm92_out == 10'd485 & go ? 5'd12 :
     fsm92_out == 10'd486 & go | fsm92_out == 10'd487 & go | fsm92_out == 10'd488 & go | fsm92_out == 10'd489 & go | fsm92_out == 10'd490 & go | fsm92_out == 10'd491 & go | fsm92_out == 10'd492 & go | fsm92_out == 10'd493 & go | fsm92_out == 10'd494 & go | fsm92_out == 10'd495 & go | fsm92_out == 10'd496 & go | fsm92_out == 10'd497 & go | fsm92_out == 10'd498 & go | fsm92_out == 10'd499 & go | fsm92_out == 10'd500 & go | fsm92_out == 10'd501 & go ? 5'd13 :
     fsm92_out == 10'd502 & go | fsm92_out == 10'd503 & go | fsm92_out == 10'd504 & go | fsm92_out == 10'd505 & go | fsm92_out == 10'd506 & go | fsm92_out == 10'd507 & go | fsm92_out == 10'd508 & go | fsm92_out == 10'd509 & go | fsm92_out == 10'd510 & go | fsm92_out == 10'd511 & go | fsm92_out == 10'd512 & go | fsm92_out == 10'd513 & go | fsm92_out == 10'd514 & go | fsm92_out == 10'd515 & go | fsm92_out == 10'd516 & go | fsm92_out == 10'd517 & go ? 5'd14 :
     fsm92_out == 10'd518 & go | fsm92_out == 10'd519 & go | fsm92_out == 10'd520 & go | fsm92_out == 10'd521 & go | fsm92_out == 10'd522 & go | fsm92_out == 10'd523 & go | fsm92_out == 10'd524 & go | fsm92_out == 10'd525 & go | fsm92_out == 10'd526 & go | fsm92_out == 10'd527 & go | fsm92_out == 10'd528 & go | fsm92_out == 10'd529 & go | fsm92_out == 10'd530 & go | fsm92_out == 10'd531 & go | fsm92_out == 10'd532 & go | fsm92_out == 10'd533 & go ? 5'd15 :
     fsm92_out == 10'd294 & go | fsm92_out == 10'd295 & go | fsm92_out == 10'd296 & go | fsm92_out == 10'd297 & go | fsm92_out == 10'd298 & go | fsm92_out == 10'd299 & go | fsm92_out == 10'd300 & go | fsm92_out == 10'd301 & go | fsm92_out == 10'd302 & go | fsm92_out == 10'd303 & go | fsm92_out == 10'd304 & go | fsm92_out == 10'd305 & go | fsm92_out == 10'd306 & go | fsm92_out == 10'd307 & go | fsm92_out == 10'd308 & go | fsm92_out == 10'd309 & go ? 5'd1 :
     fsm92_out == 10'd310 & go | fsm92_out == 10'd311 & go | fsm92_out == 10'd312 & go | fsm92_out == 10'd313 & go | fsm92_out == 10'd314 & go | fsm92_out == 10'd315 & go | fsm92_out == 10'd316 & go | fsm92_out == 10'd317 & go | fsm92_out == 10'd318 & go | fsm92_out == 10'd319 & go | fsm92_out == 10'd320 & go | fsm92_out == 10'd321 & go | fsm92_out == 10'd322 & go | fsm92_out == 10'd323 & go | fsm92_out == 10'd324 & go | fsm92_out == 10'd325 & go ? 5'd2 :
     fsm92_out == 10'd326 & go | fsm92_out == 10'd327 & go | fsm92_out == 10'd328 & go | fsm92_out == 10'd329 & go | fsm92_out == 10'd330 & go | fsm92_out == 10'd331 & go | fsm92_out == 10'd332 & go | fsm92_out == 10'd333 & go | fsm92_out == 10'd334 & go | fsm92_out == 10'd335 & go | fsm92_out == 10'd336 & go | fsm92_out == 10'd337 & go | fsm92_out == 10'd338 & go | fsm92_out == 10'd339 & go | fsm92_out == 10'd340 & go | fsm92_out == 10'd341 & go ? 5'd3 :
     fsm92_out == 10'd342 & go | fsm92_out == 10'd343 & go | fsm92_out == 10'd344 & go | fsm92_out == 10'd345 & go | fsm92_out == 10'd346 & go | fsm92_out == 10'd347 & go | fsm92_out == 10'd348 & go | fsm92_out == 10'd349 & go | fsm92_out == 10'd350 & go | fsm92_out == 10'd351 & go | fsm92_out == 10'd352 & go | fsm92_out == 10'd353 & go | fsm92_out == 10'd354 & go | fsm92_out == 10'd355 & go | fsm92_out == 10'd356 & go | fsm92_out == 10'd357 & go ? 5'd4 :
     fsm92_out == 10'd358 & go | fsm92_out == 10'd359 & go | fsm92_out == 10'd360 & go | fsm92_out == 10'd361 & go | fsm92_out == 10'd362 & go | fsm92_out == 10'd363 & go | fsm92_out == 10'd364 & go | fsm92_out == 10'd365 & go | fsm92_out == 10'd366 & go | fsm92_out == 10'd367 & go | fsm92_out == 10'd368 & go | fsm92_out == 10'd369 & go | fsm92_out == 10'd370 & go | fsm92_out == 10'd371 & go | fsm92_out == 10'd372 & go | fsm92_out == 10'd373 & go ? 5'd5 :
     fsm92_out == 10'd374 & go | fsm92_out == 10'd375 & go | fsm92_out == 10'd376 & go | fsm92_out == 10'd377 & go | fsm92_out == 10'd378 & go | fsm92_out == 10'd379 & go | fsm92_out == 10'd380 & go | fsm92_out == 10'd381 & go | fsm92_out == 10'd382 & go | fsm92_out == 10'd383 & go | fsm92_out == 10'd384 & go | fsm92_out == 10'd385 & go | fsm92_out == 10'd386 & go | fsm92_out == 10'd387 & go | fsm92_out == 10'd388 & go | fsm92_out == 10'd389 & go ? 5'd6 :
     fsm92_out == 10'd390 & go | fsm92_out == 10'd391 & go | fsm92_out == 10'd392 & go | fsm92_out == 10'd393 & go | fsm92_out == 10'd394 & go | fsm92_out == 10'd395 & go | fsm92_out == 10'd396 & go | fsm92_out == 10'd397 & go | fsm92_out == 10'd398 & go | fsm92_out == 10'd399 & go | fsm92_out == 10'd400 & go | fsm92_out == 10'd401 & go | fsm92_out == 10'd402 & go | fsm92_out == 10'd403 & go | fsm92_out == 10'd404 & go | fsm92_out == 10'd405 & go ? 5'd7 :
     fsm92_out == 10'd406 & go | fsm92_out == 10'd407 & go | fsm92_out == 10'd408 & go | fsm92_out == 10'd409 & go | fsm92_out == 10'd410 & go | fsm92_out == 10'd411 & go | fsm92_out == 10'd412 & go | fsm92_out == 10'd413 & go | fsm92_out == 10'd414 & go | fsm92_out == 10'd415 & go | fsm92_out == 10'd416 & go | fsm92_out == 10'd417 & go | fsm92_out == 10'd418 & go | fsm92_out == 10'd419 & go | fsm92_out == 10'd420 & go | fsm92_out == 10'd421 & go ? 5'd8 :
     fsm92_out == 10'd422 & go | fsm92_out == 10'd423 & go | fsm92_out == 10'd424 & go | fsm92_out == 10'd425 & go | fsm92_out == 10'd426 & go | fsm92_out == 10'd427 & go | fsm92_out == 10'd428 & go | fsm92_out == 10'd429 & go | fsm92_out == 10'd430 & go | fsm92_out == 10'd431 & go | fsm92_out == 10'd432 & go | fsm92_out == 10'd433 & go | fsm92_out == 10'd434 & go | fsm92_out == 10'd435 & go | fsm92_out == 10'd436 & go | fsm92_out == 10'd437 & go ? 5'd9 : 5'd0;
    assign out_mem_addr1 =
     fsm92_out == 10'd278 & go | fsm92_out == 10'd294 & go | fsm92_out == 10'd310 & go | fsm92_out == 10'd326 & go | fsm92_out == 10'd342 & go | fsm92_out == 10'd358 & go | fsm92_out == 10'd374 & go | fsm92_out == 10'd390 & go | fsm92_out == 10'd406 & go | fsm92_out == 10'd422 & go | fsm92_out == 10'd438 & go | fsm92_out == 10'd454 & go | fsm92_out == 10'd470 & go | fsm92_out == 10'd486 & go | fsm92_out == 10'd502 & go | fsm92_out == 10'd518 & go ? 5'd0 :
     fsm92_out == 10'd288 & go | fsm92_out == 10'd304 & go | fsm92_out == 10'd320 & go | fsm92_out == 10'd336 & go | fsm92_out == 10'd352 & go | fsm92_out == 10'd368 & go | fsm92_out == 10'd384 & go | fsm92_out == 10'd400 & go | fsm92_out == 10'd416 & go | fsm92_out == 10'd432 & go | fsm92_out == 10'd448 & go | fsm92_out == 10'd464 & go | fsm92_out == 10'd480 & go | fsm92_out == 10'd496 & go | fsm92_out == 10'd512 & go | fsm92_out == 10'd528 & go ? 5'd10 :
     fsm92_out == 10'd289 & go | fsm92_out == 10'd305 & go | fsm92_out == 10'd321 & go | fsm92_out == 10'd337 & go | fsm92_out == 10'd353 & go | fsm92_out == 10'd369 & go | fsm92_out == 10'd385 & go | fsm92_out == 10'd401 & go | fsm92_out == 10'd417 & go | fsm92_out == 10'd433 & go | fsm92_out == 10'd449 & go | fsm92_out == 10'd465 & go | fsm92_out == 10'd481 & go | fsm92_out == 10'd497 & go | fsm92_out == 10'd513 & go | fsm92_out == 10'd529 & go ? 5'd11 :
     fsm92_out == 10'd290 & go | fsm92_out == 10'd306 & go | fsm92_out == 10'd322 & go | fsm92_out == 10'd338 & go | fsm92_out == 10'd354 & go | fsm92_out == 10'd370 & go | fsm92_out == 10'd386 & go | fsm92_out == 10'd402 & go | fsm92_out == 10'd418 & go | fsm92_out == 10'd434 & go | fsm92_out == 10'd450 & go | fsm92_out == 10'd466 & go | fsm92_out == 10'd482 & go | fsm92_out == 10'd498 & go | fsm92_out == 10'd514 & go | fsm92_out == 10'd530 & go ? 5'd12 :
     fsm92_out == 10'd291 & go | fsm92_out == 10'd307 & go | fsm92_out == 10'd323 & go | fsm92_out == 10'd339 & go | fsm92_out == 10'd355 & go | fsm92_out == 10'd371 & go | fsm92_out == 10'd387 & go | fsm92_out == 10'd403 & go | fsm92_out == 10'd419 & go | fsm92_out == 10'd435 & go | fsm92_out == 10'd451 & go | fsm92_out == 10'd467 & go | fsm92_out == 10'd483 & go | fsm92_out == 10'd499 & go | fsm92_out == 10'd515 & go | fsm92_out == 10'd531 & go ? 5'd13 :
     fsm92_out == 10'd292 & go | fsm92_out == 10'd308 & go | fsm92_out == 10'd324 & go | fsm92_out == 10'd340 & go | fsm92_out == 10'd356 & go | fsm92_out == 10'd372 & go | fsm92_out == 10'd388 & go | fsm92_out == 10'd404 & go | fsm92_out == 10'd420 & go | fsm92_out == 10'd436 & go | fsm92_out == 10'd452 & go | fsm92_out == 10'd468 & go | fsm92_out == 10'd484 & go | fsm92_out == 10'd500 & go | fsm92_out == 10'd516 & go | fsm92_out == 10'd532 & go ? 5'd14 :
     fsm92_out == 10'd293 & go | fsm92_out == 10'd309 & go | fsm92_out == 10'd325 & go | fsm92_out == 10'd341 & go | fsm92_out == 10'd357 & go | fsm92_out == 10'd373 & go | fsm92_out == 10'd389 & go | fsm92_out == 10'd405 & go | fsm92_out == 10'd421 & go | fsm92_out == 10'd437 & go | fsm92_out == 10'd453 & go | fsm92_out == 10'd469 & go | fsm92_out == 10'd485 & go | fsm92_out == 10'd501 & go | fsm92_out == 10'd517 & go | fsm92_out == 10'd533 & go ? 5'd15 :
     fsm92_out == 10'd279 & go | fsm92_out == 10'd295 & go | fsm92_out == 10'd311 & go | fsm92_out == 10'd327 & go | fsm92_out == 10'd343 & go | fsm92_out == 10'd359 & go | fsm92_out == 10'd375 & go | fsm92_out == 10'd391 & go | fsm92_out == 10'd407 & go | fsm92_out == 10'd423 & go | fsm92_out == 10'd439 & go | fsm92_out == 10'd455 & go | fsm92_out == 10'd471 & go | fsm92_out == 10'd487 & go | fsm92_out == 10'd503 & go | fsm92_out == 10'd519 & go ? 5'd1 :
     fsm92_out == 10'd280 & go | fsm92_out == 10'd296 & go | fsm92_out == 10'd312 & go | fsm92_out == 10'd328 & go | fsm92_out == 10'd344 & go | fsm92_out == 10'd360 & go | fsm92_out == 10'd376 & go | fsm92_out == 10'd392 & go | fsm92_out == 10'd408 & go | fsm92_out == 10'd424 & go | fsm92_out == 10'd440 & go | fsm92_out == 10'd456 & go | fsm92_out == 10'd472 & go | fsm92_out == 10'd488 & go | fsm92_out == 10'd504 & go | fsm92_out == 10'd520 & go ? 5'd2 :
     fsm92_out == 10'd281 & go | fsm92_out == 10'd297 & go | fsm92_out == 10'd313 & go | fsm92_out == 10'd329 & go | fsm92_out == 10'd345 & go | fsm92_out == 10'd361 & go | fsm92_out == 10'd377 & go | fsm92_out == 10'd393 & go | fsm92_out == 10'd409 & go | fsm92_out == 10'd425 & go | fsm92_out == 10'd441 & go | fsm92_out == 10'd457 & go | fsm92_out == 10'd473 & go | fsm92_out == 10'd489 & go | fsm92_out == 10'd505 & go | fsm92_out == 10'd521 & go ? 5'd3 :
     fsm92_out == 10'd282 & go | fsm92_out == 10'd298 & go | fsm92_out == 10'd314 & go | fsm92_out == 10'd330 & go | fsm92_out == 10'd346 & go | fsm92_out == 10'd362 & go | fsm92_out == 10'd378 & go | fsm92_out == 10'd394 & go | fsm92_out == 10'd410 & go | fsm92_out == 10'd426 & go | fsm92_out == 10'd442 & go | fsm92_out == 10'd458 & go | fsm92_out == 10'd474 & go | fsm92_out == 10'd490 & go | fsm92_out == 10'd506 & go | fsm92_out == 10'd522 & go ? 5'd4 :
     fsm92_out == 10'd283 & go | fsm92_out == 10'd299 & go | fsm92_out == 10'd315 & go | fsm92_out == 10'd331 & go | fsm92_out == 10'd347 & go | fsm92_out == 10'd363 & go | fsm92_out == 10'd379 & go | fsm92_out == 10'd395 & go | fsm92_out == 10'd411 & go | fsm92_out == 10'd427 & go | fsm92_out == 10'd443 & go | fsm92_out == 10'd459 & go | fsm92_out == 10'd475 & go | fsm92_out == 10'd491 & go | fsm92_out == 10'd507 & go | fsm92_out == 10'd523 & go ? 5'd5 :
     fsm92_out == 10'd284 & go | fsm92_out == 10'd300 & go | fsm92_out == 10'd316 & go | fsm92_out == 10'd332 & go | fsm92_out == 10'd348 & go | fsm92_out == 10'd364 & go | fsm92_out == 10'd380 & go | fsm92_out == 10'd396 & go | fsm92_out == 10'd412 & go | fsm92_out == 10'd428 & go | fsm92_out == 10'd444 & go | fsm92_out == 10'd460 & go | fsm92_out == 10'd476 & go | fsm92_out == 10'd492 & go | fsm92_out == 10'd508 & go | fsm92_out == 10'd524 & go ? 5'd6 :
     fsm92_out == 10'd285 & go | fsm92_out == 10'd301 & go | fsm92_out == 10'd317 & go | fsm92_out == 10'd333 & go | fsm92_out == 10'd349 & go | fsm92_out == 10'd365 & go | fsm92_out == 10'd381 & go | fsm92_out == 10'd397 & go | fsm92_out == 10'd413 & go | fsm92_out == 10'd429 & go | fsm92_out == 10'd445 & go | fsm92_out == 10'd461 & go | fsm92_out == 10'd477 & go | fsm92_out == 10'd493 & go | fsm92_out == 10'd509 & go | fsm92_out == 10'd525 & go ? 5'd7 :
     fsm92_out == 10'd286 & go | fsm92_out == 10'd302 & go | fsm92_out == 10'd318 & go | fsm92_out == 10'd334 & go | fsm92_out == 10'd350 & go | fsm92_out == 10'd366 & go | fsm92_out == 10'd382 & go | fsm92_out == 10'd398 & go | fsm92_out == 10'd414 & go | fsm92_out == 10'd430 & go | fsm92_out == 10'd446 & go | fsm92_out == 10'd462 & go | fsm92_out == 10'd478 & go | fsm92_out == 10'd494 & go | fsm92_out == 10'd510 & go | fsm92_out == 10'd526 & go ? 5'd8 :
     fsm92_out == 10'd287 & go | fsm92_out == 10'd303 & go | fsm92_out == 10'd319 & go | fsm92_out == 10'd335 & go | fsm92_out == 10'd351 & go | fsm92_out == 10'd367 & go | fsm92_out == 10'd383 & go | fsm92_out == 10'd399 & go | fsm92_out == 10'd415 & go | fsm92_out == 10'd431 & go | fsm92_out == 10'd447 & go | fsm92_out == 10'd463 & go | fsm92_out == 10'd479 & go | fsm92_out == 10'd495 & go | fsm92_out == 10'd511 & go | fsm92_out == 10'd527 & go ? 5'd9 : 5'd0;
    assign out_mem_clk =
     1'b1 ? clk : 1'd0;
    assign out_mem_write_data =
     fsm92_out == 10'd278 & go ? pe_0_0_out :
     fsm92_out == 10'd279 & go ? pe_0_1_out :
     fsm92_out == 10'd288 & go ? pe_0_10_out :
     fsm92_out == 10'd289 & go ? pe_0_11_out :
     fsm92_out == 10'd290 & go ? pe_0_12_out :
     fsm92_out == 10'd291 & go ? pe_0_13_out :
     fsm92_out == 10'd292 & go ? pe_0_14_out :
     fsm92_out == 10'd293 & go ? pe_0_15_out :
     fsm92_out == 10'd280 & go ? pe_0_2_out :
     fsm92_out == 10'd281 & go ? pe_0_3_out :
     fsm92_out == 10'd282 & go ? pe_0_4_out :
     fsm92_out == 10'd283 & go ? pe_0_5_out :
     fsm92_out == 10'd284 & go ? pe_0_6_out :
     fsm92_out == 10'd285 & go ? pe_0_7_out :
     fsm92_out == 10'd286 & go ? pe_0_8_out :
     fsm92_out == 10'd287 & go ? pe_0_9_out :
     fsm92_out == 10'd438 & go ? pe_10_0_out :
     fsm92_out == 10'd439 & go ? pe_10_1_out :
     fsm92_out == 10'd448 & go ? pe_10_10_out :
     fsm92_out == 10'd449 & go ? pe_10_11_out :
     fsm92_out == 10'd450 & go ? pe_10_12_out :
     fsm92_out == 10'd451 & go ? pe_10_13_out :
     fsm92_out == 10'd452 & go ? pe_10_14_out :
     fsm92_out == 10'd453 & go ? pe_10_15_out :
     fsm92_out == 10'd440 & go ? pe_10_2_out :
     fsm92_out == 10'd441 & go ? pe_10_3_out :
     fsm92_out == 10'd442 & go ? pe_10_4_out :
     fsm92_out == 10'd443 & go ? pe_10_5_out :
     fsm92_out == 10'd444 & go ? pe_10_6_out :
     fsm92_out == 10'd445 & go ? pe_10_7_out :
     fsm92_out == 10'd446 & go ? pe_10_8_out :
     fsm92_out == 10'd447 & go ? pe_10_9_out :
     fsm92_out == 10'd454 & go ? pe_11_0_out :
     fsm92_out == 10'd455 & go ? pe_11_1_out :
     fsm92_out == 10'd464 & go ? pe_11_10_out :
     fsm92_out == 10'd465 & go ? pe_11_11_out :
     fsm92_out == 10'd466 & go ? pe_11_12_out :
     fsm92_out == 10'd467 & go ? pe_11_13_out :
     fsm92_out == 10'd468 & go ? pe_11_14_out :
     fsm92_out == 10'd469 & go ? pe_11_15_out :
     fsm92_out == 10'd456 & go ? pe_11_2_out :
     fsm92_out == 10'd457 & go ? pe_11_3_out :
     fsm92_out == 10'd458 & go ? pe_11_4_out :
     fsm92_out == 10'd459 & go ? pe_11_5_out :
     fsm92_out == 10'd460 & go ? pe_11_6_out :
     fsm92_out == 10'd461 & go ? pe_11_7_out :
     fsm92_out == 10'd462 & go ? pe_11_8_out :
     fsm92_out == 10'd463 & go ? pe_11_9_out :
     fsm92_out == 10'd470 & go ? pe_12_0_out :
     fsm92_out == 10'd471 & go ? pe_12_1_out :
     fsm92_out == 10'd480 & go ? pe_12_10_out :
     fsm92_out == 10'd481 & go ? pe_12_11_out :
     fsm92_out == 10'd482 & go ? pe_12_12_out :
     fsm92_out == 10'd483 & go ? pe_12_13_out :
     fsm92_out == 10'd484 & go ? pe_12_14_out :
     fsm92_out == 10'd485 & go ? pe_12_15_out :
     fsm92_out == 10'd472 & go ? pe_12_2_out :
     fsm92_out == 10'd473 & go ? pe_12_3_out :
     fsm92_out == 10'd474 & go ? pe_12_4_out :
     fsm92_out == 10'd475 & go ? pe_12_5_out :
     fsm92_out == 10'd476 & go ? pe_12_6_out :
     fsm92_out == 10'd477 & go ? pe_12_7_out :
     fsm92_out == 10'd478 & go ? pe_12_8_out :
     fsm92_out == 10'd479 & go ? pe_12_9_out :
     fsm92_out == 10'd486 & go ? pe_13_0_out :
     fsm92_out == 10'd487 & go ? pe_13_1_out :
     fsm92_out == 10'd496 & go ? pe_13_10_out :
     fsm92_out == 10'd497 & go ? pe_13_11_out :
     fsm92_out == 10'd498 & go ? pe_13_12_out :
     fsm92_out == 10'd499 & go ? pe_13_13_out :
     fsm92_out == 10'd500 & go ? pe_13_14_out :
     fsm92_out == 10'd501 & go ? pe_13_15_out :
     fsm92_out == 10'd488 & go ? pe_13_2_out :
     fsm92_out == 10'd489 & go ? pe_13_3_out :
     fsm92_out == 10'd490 & go ? pe_13_4_out :
     fsm92_out == 10'd491 & go ? pe_13_5_out :
     fsm92_out == 10'd492 & go ? pe_13_6_out :
     fsm92_out == 10'd493 & go ? pe_13_7_out :
     fsm92_out == 10'd494 & go ? pe_13_8_out :
     fsm92_out == 10'd495 & go ? pe_13_9_out :
     fsm92_out == 10'd502 & go ? pe_14_0_out :
     fsm92_out == 10'd503 & go ? pe_14_1_out :
     fsm92_out == 10'd512 & go ? pe_14_10_out :
     fsm92_out == 10'd513 & go ? pe_14_11_out :
     fsm92_out == 10'd514 & go ? pe_14_12_out :
     fsm92_out == 10'd515 & go ? pe_14_13_out :
     fsm92_out == 10'd516 & go ? pe_14_14_out :
     fsm92_out == 10'd517 & go ? pe_14_15_out :
     fsm92_out == 10'd504 & go ? pe_14_2_out :
     fsm92_out == 10'd505 & go ? pe_14_3_out :
     fsm92_out == 10'd506 & go ? pe_14_4_out :
     fsm92_out == 10'd507 & go ? pe_14_5_out :
     fsm92_out == 10'd508 & go ? pe_14_6_out :
     fsm92_out == 10'd509 & go ? pe_14_7_out :
     fsm92_out == 10'd510 & go ? pe_14_8_out :
     fsm92_out == 10'd511 & go ? pe_14_9_out :
     fsm92_out == 10'd518 & go ? pe_15_0_out :
     fsm92_out == 10'd519 & go ? pe_15_1_out :
     fsm92_out == 10'd528 & go ? pe_15_10_out :
     fsm92_out == 10'd529 & go ? pe_15_11_out :
     fsm92_out == 10'd530 & go ? pe_15_12_out :
     fsm92_out == 10'd531 & go ? pe_15_13_out :
     fsm92_out == 10'd532 & go ? pe_15_14_out :
     fsm92_out == 10'd533 & go ? pe_15_15_out :
     fsm92_out == 10'd520 & go ? pe_15_2_out :
     fsm92_out == 10'd521 & go ? pe_15_3_out :
     fsm92_out == 10'd522 & go ? pe_15_4_out :
     fsm92_out == 10'd523 & go ? pe_15_5_out :
     fsm92_out == 10'd524 & go ? pe_15_6_out :
     fsm92_out == 10'd525 & go ? pe_15_7_out :
     fsm92_out == 10'd526 & go ? pe_15_8_out :
     fsm92_out == 10'd527 & go ? pe_15_9_out :
     fsm92_out == 10'd294 & go ? pe_1_0_out :
     fsm92_out == 10'd295 & go ? pe_1_1_out :
     fsm92_out == 10'd304 & go ? pe_1_10_out :
     fsm92_out == 10'd305 & go ? pe_1_11_out :
     fsm92_out == 10'd306 & go ? pe_1_12_out :
     fsm92_out == 10'd307 & go ? pe_1_13_out :
     fsm92_out == 10'd308 & go ? pe_1_14_out :
     fsm92_out == 10'd309 & go ? pe_1_15_out :
     fsm92_out == 10'd296 & go ? pe_1_2_out :
     fsm92_out == 10'd297 & go ? pe_1_3_out :
     fsm92_out == 10'd298 & go ? pe_1_4_out :
     fsm92_out == 10'd299 & go ? pe_1_5_out :
     fsm92_out == 10'd300 & go ? pe_1_6_out :
     fsm92_out == 10'd301 & go ? pe_1_7_out :
     fsm92_out == 10'd302 & go ? pe_1_8_out :
     fsm92_out == 10'd303 & go ? pe_1_9_out :
     fsm92_out == 10'd310 & go ? pe_2_0_out :
     fsm92_out == 10'd311 & go ? pe_2_1_out :
     fsm92_out == 10'd320 & go ? pe_2_10_out :
     fsm92_out == 10'd321 & go ? pe_2_11_out :
     fsm92_out == 10'd322 & go ? pe_2_12_out :
     fsm92_out == 10'd323 & go ? pe_2_13_out :
     fsm92_out == 10'd324 & go ? pe_2_14_out :
     fsm92_out == 10'd325 & go ? pe_2_15_out :
     fsm92_out == 10'd312 & go ? pe_2_2_out :
     fsm92_out == 10'd313 & go ? pe_2_3_out :
     fsm92_out == 10'd314 & go ? pe_2_4_out :
     fsm92_out == 10'd315 & go ? pe_2_5_out :
     fsm92_out == 10'd316 & go ? pe_2_6_out :
     fsm92_out == 10'd317 & go ? pe_2_7_out :
     fsm92_out == 10'd318 & go ? pe_2_8_out :
     fsm92_out == 10'd319 & go ? pe_2_9_out :
     fsm92_out == 10'd326 & go ? pe_3_0_out :
     fsm92_out == 10'd327 & go ? pe_3_1_out :
     fsm92_out == 10'd336 & go ? pe_3_10_out :
     fsm92_out == 10'd337 & go ? pe_3_11_out :
     fsm92_out == 10'd338 & go ? pe_3_12_out :
     fsm92_out == 10'd339 & go ? pe_3_13_out :
     fsm92_out == 10'd340 & go ? pe_3_14_out :
     fsm92_out == 10'd341 & go ? pe_3_15_out :
     fsm92_out == 10'd328 & go ? pe_3_2_out :
     fsm92_out == 10'd329 & go ? pe_3_3_out :
     fsm92_out == 10'd330 & go ? pe_3_4_out :
     fsm92_out == 10'd331 & go ? pe_3_5_out :
     fsm92_out == 10'd332 & go ? pe_3_6_out :
     fsm92_out == 10'd333 & go ? pe_3_7_out :
     fsm92_out == 10'd334 & go ? pe_3_8_out :
     fsm92_out == 10'd335 & go ? pe_3_9_out :
     fsm92_out == 10'd342 & go ? pe_4_0_out :
     fsm92_out == 10'd343 & go ? pe_4_1_out :
     fsm92_out == 10'd352 & go ? pe_4_10_out :
     fsm92_out == 10'd353 & go ? pe_4_11_out :
     fsm92_out == 10'd354 & go ? pe_4_12_out :
     fsm92_out == 10'd355 & go ? pe_4_13_out :
     fsm92_out == 10'd356 & go ? pe_4_14_out :
     fsm92_out == 10'd357 & go ? pe_4_15_out :
     fsm92_out == 10'd344 & go ? pe_4_2_out :
     fsm92_out == 10'd345 & go ? pe_4_3_out :
     fsm92_out == 10'd346 & go ? pe_4_4_out :
     fsm92_out == 10'd347 & go ? pe_4_5_out :
     fsm92_out == 10'd348 & go ? pe_4_6_out :
     fsm92_out == 10'd349 & go ? pe_4_7_out :
     fsm92_out == 10'd350 & go ? pe_4_8_out :
     fsm92_out == 10'd351 & go ? pe_4_9_out :
     fsm92_out == 10'd358 & go ? pe_5_0_out :
     fsm92_out == 10'd359 & go ? pe_5_1_out :
     fsm92_out == 10'd368 & go ? pe_5_10_out :
     fsm92_out == 10'd369 & go ? pe_5_11_out :
     fsm92_out == 10'd370 & go ? pe_5_12_out :
     fsm92_out == 10'd371 & go ? pe_5_13_out :
     fsm92_out == 10'd372 & go ? pe_5_14_out :
     fsm92_out == 10'd373 & go ? pe_5_15_out :
     fsm92_out == 10'd360 & go ? pe_5_2_out :
     fsm92_out == 10'd361 & go ? pe_5_3_out :
     fsm92_out == 10'd362 & go ? pe_5_4_out :
     fsm92_out == 10'd363 & go ? pe_5_5_out :
     fsm92_out == 10'd364 & go ? pe_5_6_out :
     fsm92_out == 10'd365 & go ? pe_5_7_out :
     fsm92_out == 10'd366 & go ? pe_5_8_out :
     fsm92_out == 10'd367 & go ? pe_5_9_out :
     fsm92_out == 10'd374 & go ? pe_6_0_out :
     fsm92_out == 10'd375 & go ? pe_6_1_out :
     fsm92_out == 10'd384 & go ? pe_6_10_out :
     fsm92_out == 10'd385 & go ? pe_6_11_out :
     fsm92_out == 10'd386 & go ? pe_6_12_out :
     fsm92_out == 10'd387 & go ? pe_6_13_out :
     fsm92_out == 10'd388 & go ? pe_6_14_out :
     fsm92_out == 10'd389 & go ? pe_6_15_out :
     fsm92_out == 10'd376 & go ? pe_6_2_out :
     fsm92_out == 10'd377 & go ? pe_6_3_out :
     fsm92_out == 10'd378 & go ? pe_6_4_out :
     fsm92_out == 10'd379 & go ? pe_6_5_out :
     fsm92_out == 10'd380 & go ? pe_6_6_out :
     fsm92_out == 10'd381 & go ? pe_6_7_out :
     fsm92_out == 10'd382 & go ? pe_6_8_out :
     fsm92_out == 10'd383 & go ? pe_6_9_out :
     fsm92_out == 10'd390 & go ? pe_7_0_out :
     fsm92_out == 10'd391 & go ? pe_7_1_out :
     fsm92_out == 10'd400 & go ? pe_7_10_out :
     fsm92_out == 10'd401 & go ? pe_7_11_out :
     fsm92_out == 10'd402 & go ? pe_7_12_out :
     fsm92_out == 10'd403 & go ? pe_7_13_out :
     fsm92_out == 10'd404 & go ? pe_7_14_out :
     fsm92_out == 10'd405 & go ? pe_7_15_out :
     fsm92_out == 10'd392 & go ? pe_7_2_out :
     fsm92_out == 10'd393 & go ? pe_7_3_out :
     fsm92_out == 10'd394 & go ? pe_7_4_out :
     fsm92_out == 10'd395 & go ? pe_7_5_out :
     fsm92_out == 10'd396 & go ? pe_7_6_out :
     fsm92_out == 10'd397 & go ? pe_7_7_out :
     fsm92_out == 10'd398 & go ? pe_7_8_out :
     fsm92_out == 10'd399 & go ? pe_7_9_out :
     fsm92_out == 10'd406 & go ? pe_8_0_out :
     fsm92_out == 10'd407 & go ? pe_8_1_out :
     fsm92_out == 10'd416 & go ? pe_8_10_out :
     fsm92_out == 10'd417 & go ? pe_8_11_out :
     fsm92_out == 10'd418 & go ? pe_8_12_out :
     fsm92_out == 10'd419 & go ? pe_8_13_out :
     fsm92_out == 10'd420 & go ? pe_8_14_out :
     fsm92_out == 10'd421 & go ? pe_8_15_out :
     fsm92_out == 10'd408 & go ? pe_8_2_out :
     fsm92_out == 10'd409 & go ? pe_8_3_out :
     fsm92_out == 10'd410 & go ? pe_8_4_out :
     fsm92_out == 10'd411 & go ? pe_8_5_out :
     fsm92_out == 10'd412 & go ? pe_8_6_out :
     fsm92_out == 10'd413 & go ? pe_8_7_out :
     fsm92_out == 10'd414 & go ? pe_8_8_out :
     fsm92_out == 10'd415 & go ? pe_8_9_out :
     fsm92_out == 10'd422 & go ? pe_9_0_out :
     fsm92_out == 10'd423 & go ? pe_9_1_out :
     fsm92_out == 10'd432 & go ? pe_9_10_out :
     fsm92_out == 10'd433 & go ? pe_9_11_out :
     fsm92_out == 10'd434 & go ? pe_9_12_out :
     fsm92_out == 10'd435 & go ? pe_9_13_out :
     fsm92_out == 10'd436 & go ? pe_9_14_out :
     fsm92_out == 10'd437 & go ? pe_9_15_out :
     fsm92_out == 10'd424 & go ? pe_9_2_out :
     fsm92_out == 10'd425 & go ? pe_9_3_out :
     fsm92_out == 10'd426 & go ? pe_9_4_out :
     fsm92_out == 10'd427 & go ? pe_9_5_out :
     fsm92_out == 10'd428 & go ? pe_9_6_out :
     fsm92_out == 10'd429 & go ? pe_9_7_out :
     fsm92_out == 10'd430 & go ? pe_9_8_out :
     fsm92_out == 10'd431 & go ? pe_9_9_out : 32'd0;
    assign out_mem_write_en =
     fsm92_out == 10'd278 & go | fsm92_out == 10'd279 & go | fsm92_out == 10'd280 & go | fsm92_out == 10'd281 & go | fsm92_out == 10'd282 & go | fsm92_out == 10'd283 & go | fsm92_out == 10'd284 & go | fsm92_out == 10'd285 & go | fsm92_out == 10'd286 & go | fsm92_out == 10'd287 & go | fsm92_out == 10'd288 & go | fsm92_out == 10'd289 & go | fsm92_out == 10'd290 & go | fsm92_out == 10'd291 & go | fsm92_out == 10'd292 & go | fsm92_out == 10'd293 & go | fsm92_out == 10'd294 & go | fsm92_out == 10'd295 & go | fsm92_out == 10'd296 & go | fsm92_out == 10'd297 & go | fsm92_out == 10'd298 & go | fsm92_out == 10'd299 & go | fsm92_out == 10'd300 & go | fsm92_out == 10'd301 & go | fsm92_out == 10'd302 & go | fsm92_out == 10'd303 & go | fsm92_out == 10'd304 & go | fsm92_out == 10'd305 & go | fsm92_out == 10'd306 & go | fsm92_out == 10'd307 & go | fsm92_out == 10'd308 & go | fsm92_out == 10'd309 & go | fsm92_out == 10'd310 & go | fsm92_out == 10'd311 & go | fsm92_out == 10'd312 & go | fsm92_out == 10'd313 & go | fsm92_out == 10'd314 & go | fsm92_out == 10'd315 & go | fsm92_out == 10'd316 & go | fsm92_out == 10'd317 & go | fsm92_out == 10'd318 & go | fsm92_out == 10'd319 & go | fsm92_out == 10'd320 & go | fsm92_out == 10'd321 & go | fsm92_out == 10'd322 & go | fsm92_out == 10'd323 & go | fsm92_out == 10'd324 & go | fsm92_out == 10'd325 & go | fsm92_out == 10'd326 & go | fsm92_out == 10'd327 & go | fsm92_out == 10'd328 & go | fsm92_out == 10'd329 & go | fsm92_out == 10'd330 & go | fsm92_out == 10'd331 & go | fsm92_out == 10'd332 & go | fsm92_out == 10'd333 & go | fsm92_out == 10'd334 & go | fsm92_out == 10'd335 & go | fsm92_out == 10'd336 & go | fsm92_out == 10'd337 & go | fsm92_out == 10'd338 & go | fsm92_out == 10'd339 & go | fsm92_out == 10'd340 & go | fsm92_out == 10'd341 & go | fsm92_out == 10'd342 & go | fsm92_out == 10'd343 & go | fsm92_out == 10'd344 & go | fsm92_out == 10'd345 & go | fsm92_out == 10'd346 & go | fsm92_out == 10'd347 & go | fsm92_out == 10'd348 & go | fsm92_out == 10'd349 & go | fsm92_out == 10'd350 & go | fsm92_out == 10'd351 & go | fsm92_out == 10'd352 & go | fsm92_out == 10'd353 & go | fsm92_out == 10'd354 & go | fsm92_out == 10'd355 & go | fsm92_out == 10'd356 & go | fsm92_out == 10'd357 & go | fsm92_out == 10'd358 & go | fsm92_out == 10'd359 & go | fsm92_out == 10'd360 & go | fsm92_out == 10'd361 & go | fsm92_out == 10'd362 & go | fsm92_out == 10'd363 & go | fsm92_out == 10'd364 & go | fsm92_out == 10'd365 & go | fsm92_out == 10'd366 & go | fsm92_out == 10'd367 & go | fsm92_out == 10'd368 & go | fsm92_out == 10'd369 & go | fsm92_out == 10'd370 & go | fsm92_out == 10'd371 & go | fsm92_out == 10'd372 & go | fsm92_out == 10'd373 & go | fsm92_out == 10'd374 & go | fsm92_out == 10'd375 & go | fsm92_out == 10'd376 & go | fsm92_out == 10'd377 & go | fsm92_out == 10'd378 & go | fsm92_out == 10'd379 & go | fsm92_out == 10'd380 & go | fsm92_out == 10'd381 & go | fsm92_out == 10'd382 & go | fsm92_out == 10'd383 & go | fsm92_out == 10'd384 & go | fsm92_out == 10'd385 & go | fsm92_out == 10'd386 & go | fsm92_out == 10'd387 & go | fsm92_out == 10'd388 & go | fsm92_out == 10'd389 & go | fsm92_out == 10'd390 & go | fsm92_out == 10'd391 & go | fsm92_out == 10'd392 & go | fsm92_out == 10'd393 & go | fsm92_out == 10'd394 & go | fsm92_out == 10'd395 & go | fsm92_out == 10'd396 & go | fsm92_out == 10'd397 & go | fsm92_out == 10'd398 & go | fsm92_out == 10'd399 & go | fsm92_out == 10'd400 & go | fsm92_out == 10'd401 & go | fsm92_out == 10'd402 & go | fsm92_out == 10'd403 & go | fsm92_out == 10'd404 & go | fsm92_out == 10'd405 & go | fsm92_out == 10'd406 & go | fsm92_out == 10'd407 & go | fsm92_out == 10'd408 & go | fsm92_out == 10'd409 & go | fsm92_out == 10'd410 & go | fsm92_out == 10'd411 & go | fsm92_out == 10'd412 & go | fsm92_out == 10'd413 & go | fsm92_out == 10'd414 & go | fsm92_out == 10'd415 & go | fsm92_out == 10'd416 & go | fsm92_out == 10'd417 & go | fsm92_out == 10'd418 & go | fsm92_out == 10'd419 & go | fsm92_out == 10'd420 & go | fsm92_out == 10'd421 & go | fsm92_out == 10'd422 & go | fsm92_out == 10'd423 & go | fsm92_out == 10'd424 & go | fsm92_out == 10'd425 & go | fsm92_out == 10'd426 & go | fsm92_out == 10'd427 & go | fsm92_out == 10'd428 & go | fsm92_out == 10'd429 & go | fsm92_out == 10'd430 & go | fsm92_out == 10'd431 & go | fsm92_out == 10'd432 & go | fsm92_out == 10'd433 & go | fsm92_out == 10'd434 & go | fsm92_out == 10'd435 & go | fsm92_out == 10'd436 & go | fsm92_out == 10'd437 & go | fsm92_out == 10'd438 & go | fsm92_out == 10'd439 & go | fsm92_out == 10'd440 & go | fsm92_out == 10'd441 & go | fsm92_out == 10'd442 & go | fsm92_out == 10'd443 & go | fsm92_out == 10'd444 & go | fsm92_out == 10'd445 & go | fsm92_out == 10'd446 & go | fsm92_out == 10'd447 & go | fsm92_out == 10'd448 & go | fsm92_out == 10'd449 & go | fsm92_out == 10'd450 & go | fsm92_out == 10'd451 & go | fsm92_out == 10'd452 & go | fsm92_out == 10'd453 & go | fsm92_out == 10'd454 & go | fsm92_out == 10'd455 & go | fsm92_out == 10'd456 & go | fsm92_out == 10'd457 & go | fsm92_out == 10'd458 & go | fsm92_out == 10'd459 & go | fsm92_out == 10'd460 & go | fsm92_out == 10'd461 & go | fsm92_out == 10'd462 & go | fsm92_out == 10'd463 & go | fsm92_out == 10'd464 & go | fsm92_out == 10'd465 & go | fsm92_out == 10'd466 & go | fsm92_out == 10'd467 & go | fsm92_out == 10'd468 & go | fsm92_out == 10'd469 & go | fsm92_out == 10'd470 & go | fsm92_out == 10'd471 & go | fsm92_out == 10'd472 & go | fsm92_out == 10'd473 & go | fsm92_out == 10'd474 & go | fsm92_out == 10'd475 & go | fsm92_out == 10'd476 & go | fsm92_out == 10'd477 & go | fsm92_out == 10'd478 & go | fsm92_out == 10'd479 & go | fsm92_out == 10'd480 & go | fsm92_out == 10'd481 & go | fsm92_out == 10'd482 & go | fsm92_out == 10'd483 & go | fsm92_out == 10'd484 & go | fsm92_out == 10'd485 & go | fsm92_out == 10'd486 & go | fsm92_out == 10'd487 & go | fsm92_out == 10'd488 & go | fsm92_out == 10'd489 & go | fsm92_out == 10'd490 & go | fsm92_out == 10'd491 & go | fsm92_out == 10'd492 & go | fsm92_out == 10'd493 & go | fsm92_out == 10'd494 & go | fsm92_out == 10'd495 & go | fsm92_out == 10'd496 & go | fsm92_out == 10'd497 & go | fsm92_out == 10'd498 & go | fsm92_out == 10'd499 & go | fsm92_out == 10'd500 & go | fsm92_out == 10'd501 & go | fsm92_out == 10'd502 & go | fsm92_out == 10'd503 & go | fsm92_out == 10'd504 & go | fsm92_out == 10'd505 & go | fsm92_out == 10'd506 & go | fsm92_out == 10'd507 & go | fsm92_out == 10'd508 & go | fsm92_out == 10'd509 & go | fsm92_out == 10'd510 & go | fsm92_out == 10'd511 & go | fsm92_out == 10'd512 & go | fsm92_out == 10'd513 & go | fsm92_out == 10'd514 & go | fsm92_out == 10'd515 & go | fsm92_out == 10'd516 & go | fsm92_out == 10'd517 & go | fsm92_out == 10'd518 & go | fsm92_out == 10'd519 & go | fsm92_out == 10'd520 & go | fsm92_out == 10'd521 & go | fsm92_out == 10'd522 & go | fsm92_out == 10'd523 & go | fsm92_out == 10'd524 & go | fsm92_out == 10'd525 & go | fsm92_out == 10'd526 & go | fsm92_out == 10'd527 & go | fsm92_out == 10'd528 & go | fsm92_out == 10'd529 & go | fsm92_out == 10'd530 & go | fsm92_out == 10'd531 & go | fsm92_out == 10'd532 & go | fsm92_out == 10'd533 & go ? 1'd1 : 1'd0;
    assign t0_addr0 =
     fsm1_out < 1'd1 & fsm92_out == 10'd2 & go | fsm3_out < 1'd1 & fsm92_out == 10'd8 & go | fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go ? t0_idx_out : 5'd0;
    assign t0_clk =
     1'b1 ? clk : 1'd0;
    assign t10_addr0 =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? t10_idx_out : 5'd0;
    assign t10_clk =
     1'b1 ? clk : 1'd0;
    assign t11_addr0 =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? t11_idx_out : 5'd0;
    assign t11_clk =
     1'b1 ? clk : 1'd0;
    assign t12_addr0 =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? t12_idx_out : 5'd0;
    assign t12_clk =
     1'b1 ? clk : 1'd0;
    assign t13_addr0 =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? t13_idx_out : 5'd0;
    assign t13_clk =
     1'b1 ? clk : 1'd0;
    assign t14_addr0 =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? t14_idx_out : 5'd0;
    assign t14_clk =
     1'b1 ? clk : 1'd0;
    assign t15_addr0 =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? t15_idx_out : 5'd0;
    assign t15_clk =
     1'b1 ? clk : 1'd0;
    assign t1_addr0 =
     fsm3_out < 1'd1 & fsm92_out == 10'd8 & go | fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go ? t1_idx_out : 5'd0;
    assign t1_clk =
     1'b1 ? clk : 1'd0;
    assign t2_addr0 =
     fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go ? t2_idx_out : 5'd0;
    assign t2_clk =
     1'b1 ? clk : 1'd0;
    assign t3_addr0 =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? t3_idx_out : 5'd0;
    assign t3_clk =
     1'b1 ? clk : 1'd0;
    assign t4_addr0 =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? t4_idx_out : 5'd0;
    assign t4_clk =
     1'b1 ? clk : 1'd0;
    assign t5_addr0 =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? t5_idx_out : 5'd0;
    assign t5_clk =
     1'b1 ? clk : 1'd0;
    assign t6_addr0 =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? t6_idx_out : 5'd0;
    assign t6_clk =
     1'b1 ? clk : 1'd0;
    assign t7_addr0 =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? t7_idx_out : 5'd0;
    assign t7_clk =
     1'b1 ? clk : 1'd0;
    assign t8_addr0 =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? t8_idx_out : 5'd0;
    assign t8_clk =
     1'b1 ? clk : 1'd0;
    assign t9_addr0 =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? t9_idx_out : 5'd0;
    assign t9_clk =
     1'b1 ? clk : 1'd0;
    assign fsm_clk =
     1'b1 ? clk : 1'd0;
    assign fsm_in =
     fsm_out == 1'd1 ? 1'd0 :
     fsm_out != 1'd1 & fsm92_out == 10'd0 & go ? incr_out : 1'd0;
    assign fsm_write_en =
     fsm_out != 1'd1 & fsm92_out == 10'd0 & go | fsm_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm0_clk =
     1'b1 ? clk : 1'd0;
    assign fsm0_in =
     fsm0_out == 1'd1 ? 1'd0 :
     fsm0_out != 1'd1 & fsm92_out == 10'd1 & go ? incr0_out : 1'd0;
    assign fsm0_write_en =
     fsm0_out != 1'd1 & fsm92_out == 10'd1 & go | fsm0_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm1_clk =
     1'b1 ? clk : 1'd0;
    assign fsm1_in =
     fsm1_out == 1'd1 ? 1'd0 :
     fsm1_out != 1'd1 & fsm92_out == 10'd2 & go ? incr1_out : 1'd0;
    assign fsm1_write_en =
     fsm1_out != 1'd1 & fsm92_out == 10'd2 & go | fsm1_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm10_clk =
     1'b1 ? clk : 1'd0;
    assign fsm10_in =
     fsm10_out == 3'd5 ? 3'd0 :
     fsm10_out != 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go ? incr10_out : 3'd0;
    assign fsm10_write_en =
     fsm10_out != 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm10_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm11_clk =
     1'b1 ? clk : 1'd0;
    assign fsm11_in =
     fsm11_out == 1'd1 ? 1'd0 :
     fsm11_out != 1'd1 & fsm92_out == 10'd32 & go ? incr11_out : 1'd0;
    assign fsm11_write_en =
     fsm11_out != 1'd1 & fsm92_out == 10'd32 & go | fsm11_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm12_clk =
     1'b1 ? clk : 1'd0;
    assign fsm12_in =
     fsm12_out == 3'd5 ? 3'd0 :
     fsm12_out != 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go ? incr12_out : 3'd0;
    assign fsm12_write_en =
     fsm12_out != 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm12_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm13_clk =
     1'b1 ? clk : 1'd0;
    assign fsm13_in =
     fsm13_out == 1'd1 ? 1'd0 :
     fsm13_out != 1'd1 & fsm92_out == 10'd38 & go ? incr13_out : 1'd0;
    assign fsm13_write_en =
     fsm13_out != 1'd1 & fsm92_out == 10'd38 & go | fsm13_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm14_clk =
     1'b1 ? clk : 1'd0;
    assign fsm14_in =
     fsm14_out == 3'd5 ? 3'd0 :
     fsm14_out != 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go ? incr14_out : 3'd0;
    assign fsm14_write_en =
     fsm14_out != 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm14_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm15_clk =
     1'b1 ? clk : 1'd0;
    assign fsm15_in =
     fsm15_out == 1'd1 ? 1'd0 :
     fsm15_out != 1'd1 & fsm92_out == 10'd44 & go ? incr15_out : 1'd0;
    assign fsm15_write_en =
     fsm15_out != 1'd1 & fsm92_out == 10'd44 & go | fsm15_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm16_clk =
     1'b1 ? clk : 1'd0;
    assign fsm16_in =
     fsm16_out == 3'd5 ? 3'd0 :
     fsm16_out != 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go ? incr16_out : 3'd0;
    assign fsm16_write_en =
     fsm16_out != 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm16_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm17_clk =
     1'b1 ? clk : 1'd0;
    assign fsm17_in =
     fsm17_out == 1'd1 ? 1'd0 :
     fsm17_out != 1'd1 & fsm92_out == 10'd50 & go ? incr17_out : 1'd0;
    assign fsm17_write_en =
     fsm17_out != 1'd1 & fsm92_out == 10'd50 & go | fsm17_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm18_clk =
     1'b1 ? clk : 1'd0;
    assign fsm18_in =
     fsm18_out == 3'd5 ? 3'd0 :
     fsm18_out != 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go ? incr18_out : 3'd0;
    assign fsm18_write_en =
     fsm18_out != 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm18_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm19_clk =
     1'b1 ? clk : 1'd0;
    assign fsm19_in =
     fsm19_out == 1'd1 ? 1'd0 :
     fsm19_out != 1'd1 & fsm92_out == 10'd56 & go ? incr19_out : 1'd0;
    assign fsm19_write_en =
     fsm19_out != 1'd1 & fsm92_out == 10'd56 & go | fsm19_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm2_clk =
     1'b1 ? clk : 1'd0;
    assign fsm2_in =
     fsm2_out == 3'd5 ? 3'd0 :
     fsm2_out != 3'd5 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go ? incr2_out : 3'd0;
    assign fsm2_write_en =
     fsm2_out != 3'd5 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm2_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm20_clk =
     1'b1 ? clk : 1'd0;
    assign fsm20_in =
     fsm20_out == 3'd5 ? 3'd0 :
     fsm20_out != 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go ? incr20_out : 3'd0;
    assign fsm20_write_en =
     fsm20_out != 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm20_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm21_clk =
     1'b1 ? clk : 1'd0;
    assign fsm21_in =
     fsm21_out == 1'd1 ? 1'd0 :
     fsm21_out != 1'd1 & fsm92_out == 10'd62 & go ? incr21_out : 1'd0;
    assign fsm21_write_en =
     fsm21_out != 1'd1 & fsm92_out == 10'd62 & go | fsm21_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm22_clk =
     1'b1 ? clk : 1'd0;
    assign fsm22_in =
     fsm22_out == 3'd5 ? 3'd0 :
     fsm22_out != 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go ? incr22_out : 3'd0;
    assign fsm22_write_en =
     fsm22_out != 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm22_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm23_clk =
     1'b1 ? clk : 1'd0;
    assign fsm23_in =
     fsm23_out == 1'd1 ? 1'd0 :
     fsm23_out != 1'd1 & fsm92_out == 10'd68 & go ? incr23_out : 1'd0;
    assign fsm23_write_en =
     fsm23_out != 1'd1 & fsm92_out == 10'd68 & go | fsm23_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm24_clk =
     1'b1 ? clk : 1'd0;
    assign fsm24_in =
     fsm24_out == 3'd5 ? 3'd0 :
     fsm24_out != 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go ? incr24_out : 3'd0;
    assign fsm24_write_en =
     fsm24_out != 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm24_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm25_clk =
     1'b1 ? clk : 1'd0;
    assign fsm25_in =
     fsm25_out == 1'd1 ? 1'd0 :
     fsm25_out != 1'd1 & fsm92_out == 10'd74 & go ? incr25_out : 1'd0;
    assign fsm25_write_en =
     fsm25_out != 1'd1 & fsm92_out == 10'd74 & go | fsm25_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm26_clk =
     1'b1 ? clk : 1'd0;
    assign fsm26_in =
     fsm26_out == 3'd5 ? 3'd0 :
     fsm26_out != 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go ? incr26_out : 3'd0;
    assign fsm26_write_en =
     fsm26_out != 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm26_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm27_clk =
     1'b1 ? clk : 1'd0;
    assign fsm27_in =
     fsm27_out == 1'd1 ? 1'd0 :
     fsm27_out != 1'd1 & fsm92_out == 10'd80 & go ? incr27_out : 1'd0;
    assign fsm27_write_en =
     fsm27_out != 1'd1 & fsm92_out == 10'd80 & go | fsm27_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm28_clk =
     1'b1 ? clk : 1'd0;
    assign fsm28_in =
     fsm28_out == 3'd5 ? 3'd0 :
     fsm28_out != 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go ? incr28_out : 3'd0;
    assign fsm28_write_en =
     fsm28_out != 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm28_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm29_clk =
     1'b1 ? clk : 1'd0;
    assign fsm29_in =
     fsm29_out == 1'd1 ? 1'd0 :
     fsm29_out != 1'd1 & fsm92_out == 10'd86 & go ? incr29_out : 1'd0;
    assign fsm29_write_en =
     fsm29_out != 1'd1 & fsm92_out == 10'd86 & go | fsm29_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm3_clk =
     1'b1 ? clk : 1'd0;
    assign fsm3_in =
     fsm3_out == 1'd1 ? 1'd0 :
     fsm3_out != 1'd1 & fsm92_out == 10'd8 & go ? incr3_out : 1'd0;
    assign fsm3_write_en =
     fsm3_out != 1'd1 & fsm92_out == 10'd8 & go | fsm3_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm30_clk =
     1'b1 ? clk : 1'd0;
    assign fsm30_in =
     fsm30_out == 3'd5 ? 3'd0 :
     fsm30_out != 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go ? incr30_out : 3'd0;
    assign fsm30_write_en =
     fsm30_out != 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm30_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm31_clk =
     1'b1 ? clk : 1'd0;
    assign fsm31_in =
     fsm31_out == 1'd1 ? 1'd0 :
     fsm31_out != 1'd1 & fsm92_out == 10'd92 & go ? incr31_out : 1'd0;
    assign fsm31_write_en =
     fsm31_out != 1'd1 & fsm92_out == 10'd92 & go | fsm31_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm32_clk =
     1'b1 ? clk : 1'd0;
    assign fsm32_in =
     fsm32_out == 3'd5 ? 3'd0 :
     fsm32_out != 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go ? incr32_out : 3'd0;
    assign fsm32_write_en =
     fsm32_out != 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm32_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm33_clk =
     1'b1 ? clk : 1'd0;
    assign fsm33_in =
     fsm33_out == 1'd1 ? 1'd0 :
     fsm33_out != 1'd1 & fsm92_out == 10'd98 & go ? incr33_out : 1'd0;
    assign fsm33_write_en =
     fsm33_out != 1'd1 & fsm92_out == 10'd98 & go | fsm33_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm34_clk =
     1'b1 ? clk : 1'd0;
    assign fsm34_in =
     fsm34_out == 3'd5 ? 3'd0 :
     fsm34_out != 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? incr34_out : 3'd0;
    assign fsm34_write_en =
     fsm34_out != 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm34_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm35_clk =
     1'b1 ? clk : 1'd0;
    assign fsm35_in =
     fsm35_out == 1'd1 ? 1'd0 :
     fsm35_out != 1'd1 & fsm92_out == 10'd104 & go ? incr35_out : 1'd0;
    assign fsm35_write_en =
     fsm35_out != 1'd1 & fsm92_out == 10'd104 & go | fsm35_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm36_clk =
     1'b1 ? clk : 1'd0;
    assign fsm36_in =
     fsm36_out == 3'd5 ? 3'd0 :
     fsm36_out != 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? incr36_out : 3'd0;
    assign fsm36_write_en =
     fsm36_out != 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm36_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm37_clk =
     1'b1 ? clk : 1'd0;
    assign fsm37_in =
     fsm37_out == 1'd1 ? 1'd0 :
     fsm37_out != 1'd1 & fsm92_out == 10'd110 & go ? incr37_out : 1'd0;
    assign fsm37_write_en =
     fsm37_out != 1'd1 & fsm92_out == 10'd110 & go | fsm37_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm38_clk =
     1'b1 ? clk : 1'd0;
    assign fsm38_in =
     fsm38_out == 3'd5 ? 3'd0 :
     fsm38_out != 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? incr38_out : 3'd0;
    assign fsm38_write_en =
     fsm38_out != 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm38_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm39_clk =
     1'b1 ? clk : 1'd0;
    assign fsm39_in =
     fsm39_out == 1'd1 ? 1'd0 :
     fsm39_out != 1'd1 & fsm92_out == 10'd116 & go ? incr39_out : 1'd0;
    assign fsm39_write_en =
     fsm39_out != 1'd1 & fsm92_out == 10'd116 & go | fsm39_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm4_clk =
     1'b1 ? clk : 1'd0;
    assign fsm4_in =
     fsm4_out == 3'd5 ? 3'd0 :
     fsm4_out != 3'd5 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go ? incr4_out : 3'd0;
    assign fsm4_write_en =
     fsm4_out != 3'd5 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm4_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm40_clk =
     1'b1 ? clk : 1'd0;
    assign fsm40_in =
     fsm40_out == 3'd5 ? 3'd0 :
     fsm40_out != 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? incr40_out : 3'd0;
    assign fsm40_write_en =
     fsm40_out != 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm40_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm41_clk =
     1'b1 ? clk : 1'd0;
    assign fsm41_in =
     fsm41_out == 1'd1 ? 1'd0 :
     fsm41_out != 1'd1 & fsm92_out == 10'd122 & go ? incr41_out : 1'd0;
    assign fsm41_write_en =
     fsm41_out != 1'd1 & fsm92_out == 10'd122 & go | fsm41_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm42_clk =
     1'b1 ? clk : 1'd0;
    assign fsm42_in =
     fsm42_out == 3'd5 ? 3'd0 :
     fsm42_out != 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? incr42_out : 3'd0;
    assign fsm42_write_en =
     fsm42_out != 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm42_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm43_clk =
     1'b1 ? clk : 1'd0;
    assign fsm43_in =
     fsm43_out == 1'd1 ? 1'd0 :
     fsm43_out != 1'd1 & fsm92_out == 10'd128 & go ? incr43_out : 1'd0;
    assign fsm43_write_en =
     fsm43_out != 1'd1 & fsm92_out == 10'd128 & go | fsm43_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm44_clk =
     1'b1 ? clk : 1'd0;
    assign fsm44_in =
     fsm44_out == 3'd5 ? 3'd0 :
     fsm44_out != 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? incr44_out : 3'd0;
    assign fsm44_write_en =
     fsm44_out != 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm44_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm45_clk =
     1'b1 ? clk : 1'd0;
    assign fsm45_in =
     fsm45_out == 1'd1 ? 1'd0 :
     fsm45_out != 1'd1 & fsm92_out == 10'd134 & go ? incr45_out : 1'd0;
    assign fsm45_write_en =
     fsm45_out != 1'd1 & fsm92_out == 10'd134 & go | fsm45_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm46_clk =
     1'b1 ? clk : 1'd0;
    assign fsm46_in =
     fsm46_out == 3'd5 ? 3'd0 :
     fsm46_out != 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? incr46_out : 3'd0;
    assign fsm46_write_en =
     fsm46_out != 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm46_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm47_clk =
     1'b1 ? clk : 1'd0;
    assign fsm47_in =
     fsm47_out == 1'd1 ? 1'd0 :
     fsm47_out != 1'd1 & fsm92_out == 10'd140 & go ? incr47_out : 1'd0;
    assign fsm47_write_en =
     fsm47_out != 1'd1 & fsm92_out == 10'd140 & go | fsm47_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm48_clk =
     1'b1 ? clk : 1'd0;
    assign fsm48_in =
     fsm48_out == 3'd5 ? 3'd0 :
     fsm48_out != 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? incr48_out : 3'd0;
    assign fsm48_write_en =
     fsm48_out != 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm48_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm49_clk =
     1'b1 ? clk : 1'd0;
    assign fsm49_in =
     fsm49_out == 1'd1 ? 1'd0 :
     fsm49_out != 1'd1 & fsm92_out == 10'd146 & go ? incr49_out : 1'd0;
    assign fsm49_write_en =
     fsm49_out != 1'd1 & fsm92_out == 10'd146 & go | fsm49_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm5_clk =
     1'b1 ? clk : 1'd0;
    assign fsm5_in =
     fsm5_out == 1'd1 ? 1'd0 :
     fsm5_out != 1'd1 & fsm92_out == 10'd14 & go ? incr5_out : 1'd0;
    assign fsm5_write_en =
     fsm5_out != 1'd1 & fsm92_out == 10'd14 & go | fsm5_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm50_clk =
     1'b1 ? clk : 1'd0;
    assign fsm50_in =
     fsm50_out == 3'd5 ? 3'd0 :
     fsm50_out != 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? incr50_out : 3'd0;
    assign fsm50_write_en =
     fsm50_out != 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm50_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm51_clk =
     1'b1 ? clk : 1'd0;
    assign fsm51_in =
     fsm51_out == 1'd1 ? 1'd0 :
     fsm51_out != 1'd1 & fsm92_out == 10'd152 & go ? incr51_out : 1'd0;
    assign fsm51_write_en =
     fsm51_out != 1'd1 & fsm92_out == 10'd152 & go | fsm51_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm52_clk =
     1'b1 ? clk : 1'd0;
    assign fsm52_in =
     fsm52_out == 3'd5 ? 3'd0 :
     fsm52_out != 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? incr52_out : 3'd0;
    assign fsm52_write_en =
     fsm52_out != 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm52_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm53_clk =
     1'b1 ? clk : 1'd0;
    assign fsm53_in =
     fsm53_out == 1'd1 ? 1'd0 :
     fsm53_out != 1'd1 & fsm92_out == 10'd158 & go ? incr53_out : 1'd0;
    assign fsm53_write_en =
     fsm53_out != 1'd1 & fsm92_out == 10'd158 & go | fsm53_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm54_clk =
     1'b1 ? clk : 1'd0;
    assign fsm54_in =
     fsm54_out == 3'd5 ? 3'd0 :
     fsm54_out != 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? incr54_out : 3'd0;
    assign fsm54_write_en =
     fsm54_out != 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm54_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm55_clk =
     1'b1 ? clk : 1'd0;
    assign fsm55_in =
     fsm55_out == 1'd1 ? 1'd0 :
     fsm55_out != 1'd1 & fsm92_out == 10'd164 & go ? incr55_out : 1'd0;
    assign fsm55_write_en =
     fsm55_out != 1'd1 & fsm92_out == 10'd164 & go | fsm55_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm56_clk =
     1'b1 ? clk : 1'd0;
    assign fsm56_in =
     fsm56_out == 3'd5 ? 3'd0 :
     fsm56_out != 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? incr56_out : 3'd0;
    assign fsm56_write_en =
     fsm56_out != 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm56_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm57_clk =
     1'b1 ? clk : 1'd0;
    assign fsm57_in =
     fsm57_out == 1'd1 ? 1'd0 :
     fsm57_out != 1'd1 & fsm92_out == 10'd170 & go ? incr57_out : 1'd0;
    assign fsm57_write_en =
     fsm57_out != 1'd1 & fsm92_out == 10'd170 & go | fsm57_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm58_clk =
     1'b1 ? clk : 1'd0;
    assign fsm58_in =
     fsm58_out == 3'd5 ? 3'd0 :
     fsm58_out != 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? incr58_out : 3'd0;
    assign fsm58_write_en =
     fsm58_out != 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm58_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm59_clk =
     1'b1 ? clk : 1'd0;
    assign fsm59_in =
     fsm59_out == 1'd1 ? 1'd0 :
     fsm59_out != 1'd1 & fsm92_out == 10'd176 & go ? incr59_out : 1'd0;
    assign fsm59_write_en =
     fsm59_out != 1'd1 & fsm92_out == 10'd176 & go | fsm59_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm6_clk =
     1'b1 ? clk : 1'd0;
    assign fsm6_in =
     fsm6_out == 3'd5 ? 3'd0 :
     fsm6_out != 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go ? incr6_out : 3'd0;
    assign fsm6_write_en =
     fsm6_out != 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm6_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm60_clk =
     1'b1 ? clk : 1'd0;
    assign fsm60_in =
     fsm60_out == 3'd5 ? 3'd0 :
     fsm60_out != 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? incr60_out : 3'd0;
    assign fsm60_write_en =
     fsm60_out != 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm60_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm61_clk =
     1'b1 ? clk : 1'd0;
    assign fsm61_in =
     fsm61_out == 1'd1 ? 1'd0 :
     fsm61_out != 1'd1 & fsm92_out == 10'd182 & go ? incr61_out : 1'd0;
    assign fsm61_write_en =
     fsm61_out != 1'd1 & fsm92_out == 10'd182 & go | fsm61_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm62_clk =
     1'b1 ? clk : 1'd0;
    assign fsm62_in =
     fsm62_out == 3'd5 ? 3'd0 :
     fsm62_out != 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? incr62_out : 3'd0;
    assign fsm62_write_en =
     fsm62_out != 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm62_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm63_clk =
     1'b1 ? clk : 1'd0;
    assign fsm63_in =
     fsm63_out == 1'd1 ? 1'd0 :
     fsm63_out != 1'd1 & fsm92_out == 10'd188 & go ? incr63_out : 1'd0;
    assign fsm63_write_en =
     fsm63_out != 1'd1 & fsm92_out == 10'd188 & go | fsm63_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm64_clk =
     1'b1 ? clk : 1'd0;
    assign fsm64_in =
     fsm64_out == 3'd5 ? 3'd0 :
     fsm64_out != 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? incr64_out : 3'd0;
    assign fsm64_write_en =
     fsm64_out != 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm64_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm65_clk =
     1'b1 ? clk : 1'd0;
    assign fsm65_in =
     fsm65_out == 1'd1 ? 1'd0 :
     fsm65_out != 1'd1 & fsm92_out == 10'd194 & go ? incr65_out : 1'd0;
    assign fsm65_write_en =
     fsm65_out != 1'd1 & fsm92_out == 10'd194 & go | fsm65_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm66_clk =
     1'b1 ? clk : 1'd0;
    assign fsm66_in =
     fsm66_out == 3'd5 ? 3'd0 :
     fsm66_out != 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? incr66_out : 3'd0;
    assign fsm66_write_en =
     fsm66_out != 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm66_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm67_clk =
     1'b1 ? clk : 1'd0;
    assign fsm67_in =
     fsm67_out == 1'd1 ? 1'd0 :
     fsm67_out != 1'd1 & fsm92_out == 10'd200 & go ? incr67_out : 1'd0;
    assign fsm67_write_en =
     fsm67_out != 1'd1 & fsm92_out == 10'd200 & go | fsm67_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm68_clk =
     1'b1 ? clk : 1'd0;
    assign fsm68_in =
     fsm68_out == 3'd5 ? 3'd0 :
     fsm68_out != 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? incr68_out : 3'd0;
    assign fsm68_write_en =
     fsm68_out != 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm68_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm69_clk =
     1'b1 ? clk : 1'd0;
    assign fsm69_in =
     fsm69_out == 1'd1 ? 1'd0 :
     fsm69_out != 1'd1 & fsm92_out == 10'd206 & go ? incr69_out : 1'd0;
    assign fsm69_write_en =
     fsm69_out != 1'd1 & fsm92_out == 10'd206 & go | fsm69_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm7_clk =
     1'b1 ? clk : 1'd0;
    assign fsm7_in =
     fsm7_out == 1'd1 ? 1'd0 :
     fsm7_out != 1'd1 & fsm92_out == 10'd20 & go ? incr7_out : 1'd0;
    assign fsm7_write_en =
     fsm7_out != 1'd1 & fsm92_out == 10'd20 & go | fsm7_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm70_clk =
     1'b1 ? clk : 1'd0;
    assign fsm70_in =
     fsm70_out == 3'd5 ? 3'd0 :
     fsm70_out != 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? incr70_out : 3'd0;
    assign fsm70_write_en =
     fsm70_out != 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm70_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm71_clk =
     1'b1 ? clk : 1'd0;
    assign fsm71_in =
     fsm71_out == 1'd1 ? 1'd0 :
     fsm71_out != 1'd1 & fsm92_out == 10'd212 & go ? incr71_out : 1'd0;
    assign fsm71_write_en =
     fsm71_out != 1'd1 & fsm92_out == 10'd212 & go | fsm71_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm72_clk =
     1'b1 ? clk : 1'd0;
    assign fsm72_in =
     fsm72_out == 3'd5 ? 3'd0 :
     fsm72_out != 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? incr72_out : 3'd0;
    assign fsm72_write_en =
     fsm72_out != 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm72_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm73_clk =
     1'b1 ? clk : 1'd0;
    assign fsm73_in =
     fsm73_out == 1'd1 ? 1'd0 :
     fsm73_out != 1'd1 & fsm92_out == 10'd218 & go ? incr73_out : 1'd0;
    assign fsm73_write_en =
     fsm73_out != 1'd1 & fsm92_out == 10'd218 & go | fsm73_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm74_clk =
     1'b1 ? clk : 1'd0;
    assign fsm74_in =
     fsm74_out == 3'd5 ? 3'd0 :
     fsm74_out != 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? incr74_out : 3'd0;
    assign fsm74_write_en =
     fsm74_out != 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm74_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm75_clk =
     1'b1 ? clk : 1'd0;
    assign fsm75_in =
     fsm75_out == 1'd1 ? 1'd0 :
     fsm75_out != 1'd1 & fsm92_out == 10'd224 & go ? incr75_out : 1'd0;
    assign fsm75_write_en =
     fsm75_out != 1'd1 & fsm92_out == 10'd224 & go | fsm75_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm76_clk =
     1'b1 ? clk : 1'd0;
    assign fsm76_in =
     fsm76_out == 3'd5 ? 3'd0 :
     fsm76_out != 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? incr76_out : 3'd0;
    assign fsm76_write_en =
     fsm76_out != 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm76_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm77_clk =
     1'b1 ? clk : 1'd0;
    assign fsm77_in =
     fsm77_out == 1'd1 ? 1'd0 :
     fsm77_out != 1'd1 & fsm92_out == 10'd230 & go ? incr77_out : 1'd0;
    assign fsm77_write_en =
     fsm77_out != 1'd1 & fsm92_out == 10'd230 & go | fsm77_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm78_clk =
     1'b1 ? clk : 1'd0;
    assign fsm78_in =
     fsm78_out == 3'd5 ? 3'd0 :
     fsm78_out != 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? incr78_out : 3'd0;
    assign fsm78_write_en =
     fsm78_out != 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm78_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm79_clk =
     1'b1 ? clk : 1'd0;
    assign fsm79_in =
     fsm79_out == 1'd1 ? 1'd0 :
     fsm79_out != 1'd1 & fsm92_out == 10'd236 & go ? incr79_out : 1'd0;
    assign fsm79_write_en =
     fsm79_out != 1'd1 & fsm92_out == 10'd236 & go | fsm79_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm8_clk =
     1'b1 ? clk : 1'd0;
    assign fsm8_in =
     fsm8_out == 3'd5 ? 3'd0 :
     fsm8_out != 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go ? incr8_out : 3'd0;
    assign fsm8_write_en =
     fsm8_out != 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm8_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm80_clk =
     1'b1 ? clk : 1'd0;
    assign fsm80_in =
     fsm80_out == 3'd5 ? 3'd0 :
     fsm80_out != 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? incr80_out : 3'd0;
    assign fsm80_write_en =
     fsm80_out != 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm80_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm81_clk =
     1'b1 ? clk : 1'd0;
    assign fsm81_in =
     fsm81_out == 1'd1 ? 1'd0 :
     fsm81_out != 1'd1 & fsm92_out == 10'd242 & go ? incr81_out : 1'd0;
    assign fsm81_write_en =
     fsm81_out != 1'd1 & fsm92_out == 10'd242 & go | fsm81_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm82_clk =
     1'b1 ? clk : 1'd0;
    assign fsm82_in =
     fsm82_out == 3'd5 ? 3'd0 :
     fsm82_out != 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? incr82_out : 3'd0;
    assign fsm82_write_en =
     fsm82_out != 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm82_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm83_clk =
     1'b1 ? clk : 1'd0;
    assign fsm83_in =
     fsm83_out == 1'd1 ? 1'd0 :
     fsm83_out != 1'd1 & fsm92_out == 10'd248 & go ? incr83_out : 1'd0;
    assign fsm83_write_en =
     fsm83_out != 1'd1 & fsm92_out == 10'd248 & go | fsm83_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm84_clk =
     1'b1 ? clk : 1'd0;
    assign fsm84_in =
     fsm84_out == 3'd5 ? 3'd0 :
     fsm84_out != 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? incr84_out : 3'd0;
    assign fsm84_write_en =
     fsm84_out != 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm84_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm85_clk =
     1'b1 ? clk : 1'd0;
    assign fsm85_in =
     fsm85_out == 1'd1 ? 1'd0 :
     fsm85_out != 1'd1 & fsm92_out == 10'd254 & go ? incr85_out : 1'd0;
    assign fsm85_write_en =
     fsm85_out != 1'd1 & fsm92_out == 10'd254 & go | fsm85_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm86_clk =
     1'b1 ? clk : 1'd0;
    assign fsm86_in =
     fsm86_out == 3'd5 ? 3'd0 :
     fsm86_out != 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go ? incr86_out : 3'd0;
    assign fsm86_write_en =
     fsm86_out != 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm86_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm87_clk =
     1'b1 ? clk : 1'd0;
    assign fsm87_in =
     fsm87_out == 1'd1 ? 1'd0 :
     fsm87_out != 1'd1 & fsm92_out == 10'd260 & go ? incr87_out : 1'd0;
    assign fsm87_write_en =
     fsm87_out != 1'd1 & fsm92_out == 10'd260 & go | fsm87_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm88_clk =
     1'b1 ? clk : 1'd0;
    assign fsm88_in =
     fsm88_out == 3'd5 ? 3'd0 :
     fsm88_out != 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go ? incr88_out : 3'd0;
    assign fsm88_write_en =
     fsm88_out != 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go | fsm88_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm89_clk =
     1'b1 ? clk : 1'd0;
    assign fsm89_in =
     fsm89_out == 1'd1 ? 1'd0 :
     fsm89_out != 1'd1 & fsm92_out == 10'd266 & go ? incr89_out : 1'd0;
    assign fsm89_write_en =
     fsm89_out != 1'd1 & fsm92_out == 10'd266 & go | fsm89_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm9_clk =
     1'b1 ? clk : 1'd0;
    assign fsm9_in =
     fsm9_out == 1'd1 ? 1'd0 :
     fsm9_out != 1'd1 & fsm92_out == 10'd26 & go ? incr9_out : 1'd0;
    assign fsm9_write_en =
     fsm9_out != 1'd1 & fsm92_out == 10'd26 & go | fsm9_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm90_clk =
     1'b1 ? clk : 1'd0;
    assign fsm90_in =
     fsm90_out == 3'd5 ? 3'd0 :
     fsm90_out != 3'd5 & fsm92_out >= 10'd267 & fsm92_out < 10'd272 & go ? incr90_out : 3'd0;
    assign fsm90_write_en =
     fsm90_out != 3'd5 & fsm92_out >= 10'd267 & fsm92_out < 10'd272 & go | fsm90_out == 3'd5 ? 1'd1 : 1'd0;
    assign fsm91_clk =
     1'b1 ? clk : 1'd0;
    assign fsm91_in =
     fsm91_out == 1'd1 ? 1'd0 :
     fsm91_out != 1'd1 & fsm92_out == 10'd272 & go ? incr91_out : 1'd0;
    assign fsm91_write_en =
     fsm91_out != 1'd1 & fsm92_out == 10'd272 & go | fsm91_out == 1'd1 ? 1'd1 : 1'd0;
    assign fsm92_clk =
     1'b1 ? clk : 1'd0;
    assign fsm92_in =
     fsm92_out == 10'd534 ? 10'd0 :
     fsm92_out != 10'd534 & go ? incr92_out : 10'd0;
    assign fsm92_write_en =
     fsm92_out != 10'd534 & go | fsm92_out == 10'd534 ? 1'd1 : 1'd0;
    assign incr_left =
     fsm92_out == 10'd0 & go ? 1'd1 : 1'd0;
    assign incr_right =
     fsm92_out == 10'd0 & go ? fsm_out : 1'd0;
    assign incr0_left =
     fsm92_out == 10'd1 & go ? 1'd1 : 1'd0;
    assign incr0_right =
     fsm92_out == 10'd1 & go ? fsm0_out : 1'd0;
    assign incr1_left =
     fsm92_out == 10'd2 & go ? 1'd1 : 1'd0;
    assign incr1_right =
     fsm92_out == 10'd2 & go ? fsm1_out : 1'd0;
    assign incr10_left =
     fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go ? 3'd1 : 3'd0;
    assign incr10_right =
     fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go ? fsm10_out : 3'd0;
    assign incr11_left =
     fsm92_out == 10'd32 & go ? 1'd1 : 1'd0;
    assign incr11_right =
     fsm92_out == 10'd32 & go ? fsm11_out : 1'd0;
    assign incr12_left =
     fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go ? 3'd1 : 3'd0;
    assign incr12_right =
     fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go ? fsm12_out : 3'd0;
    assign incr13_left =
     fsm92_out == 10'd38 & go ? 1'd1 : 1'd0;
    assign incr13_right =
     fsm92_out == 10'd38 & go ? fsm13_out : 1'd0;
    assign incr14_left =
     fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go ? 3'd1 : 3'd0;
    assign incr14_right =
     fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go ? fsm14_out : 3'd0;
    assign incr15_left =
     fsm92_out == 10'd44 & go ? 1'd1 : 1'd0;
    assign incr15_right =
     fsm92_out == 10'd44 & go ? fsm15_out : 1'd0;
    assign incr16_left =
     fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go ? 3'd1 : 3'd0;
    assign incr16_right =
     fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go ? fsm16_out : 3'd0;
    assign incr17_left =
     fsm92_out == 10'd50 & go ? 1'd1 : 1'd0;
    assign incr17_right =
     fsm92_out == 10'd50 & go ? fsm17_out : 1'd0;
    assign incr18_left =
     fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go ? 3'd1 : 3'd0;
    assign incr18_right =
     fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go ? fsm18_out : 3'd0;
    assign incr19_left =
     fsm92_out == 10'd56 & go ? 1'd1 : 1'd0;
    assign incr19_right =
     fsm92_out == 10'd56 & go ? fsm19_out : 1'd0;
    assign incr2_left =
     fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go ? 3'd1 : 3'd0;
    assign incr2_right =
     fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go ? fsm2_out : 3'd0;
    assign incr20_left =
     fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go ? 3'd1 : 3'd0;
    assign incr20_right =
     fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go ? fsm20_out : 3'd0;
    assign incr21_left =
     fsm92_out == 10'd62 & go ? 1'd1 : 1'd0;
    assign incr21_right =
     fsm92_out == 10'd62 & go ? fsm21_out : 1'd0;
    assign incr22_left =
     fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go ? 3'd1 : 3'd0;
    assign incr22_right =
     fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go ? fsm22_out : 3'd0;
    assign incr23_left =
     fsm92_out == 10'd68 & go ? 1'd1 : 1'd0;
    assign incr23_right =
     fsm92_out == 10'd68 & go ? fsm23_out : 1'd0;
    assign incr24_left =
     fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go ? 3'd1 : 3'd0;
    assign incr24_right =
     fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go ? fsm24_out : 3'd0;
    assign incr25_left =
     fsm92_out == 10'd74 & go ? 1'd1 : 1'd0;
    assign incr25_right =
     fsm92_out == 10'd74 & go ? fsm25_out : 1'd0;
    assign incr26_left =
     fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go ? 3'd1 : 3'd0;
    assign incr26_right =
     fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go ? fsm26_out : 3'd0;
    assign incr27_left =
     fsm92_out == 10'd80 & go ? 1'd1 : 1'd0;
    assign incr27_right =
     fsm92_out == 10'd80 & go ? fsm27_out : 1'd0;
    assign incr28_left =
     fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go ? 3'd1 : 3'd0;
    assign incr28_right =
     fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go ? fsm28_out : 3'd0;
    assign incr29_left =
     fsm92_out == 10'd86 & go ? 1'd1 : 1'd0;
    assign incr29_right =
     fsm92_out == 10'd86 & go ? fsm29_out : 1'd0;
    assign incr3_left =
     fsm92_out == 10'd8 & go ? 1'd1 : 1'd0;
    assign incr3_right =
     fsm92_out == 10'd8 & go ? fsm3_out : 1'd0;
    assign incr30_left =
     fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go ? 3'd1 : 3'd0;
    assign incr30_right =
     fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go ? fsm30_out : 3'd0;
    assign incr31_left =
     fsm92_out == 10'd92 & go ? 1'd1 : 1'd0;
    assign incr31_right =
     fsm92_out == 10'd92 & go ? fsm31_out : 1'd0;
    assign incr32_left =
     fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go ? 3'd1 : 3'd0;
    assign incr32_right =
     fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go ? fsm32_out : 3'd0;
    assign incr33_left =
     fsm92_out == 10'd98 & go ? 1'd1 : 1'd0;
    assign incr33_right =
     fsm92_out == 10'd98 & go ? fsm33_out : 1'd0;
    assign incr34_left =
     fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? 3'd1 : 3'd0;
    assign incr34_right =
     fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? fsm34_out : 3'd0;
    assign incr35_left =
     fsm92_out == 10'd104 & go ? 1'd1 : 1'd0;
    assign incr35_right =
     fsm92_out == 10'd104 & go ? fsm35_out : 1'd0;
    assign incr36_left =
     fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? 3'd1 : 3'd0;
    assign incr36_right =
     fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? fsm36_out : 3'd0;
    assign incr37_left =
     fsm92_out == 10'd110 & go ? 1'd1 : 1'd0;
    assign incr37_right =
     fsm92_out == 10'd110 & go ? fsm37_out : 1'd0;
    assign incr38_left =
     fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? 3'd1 : 3'd0;
    assign incr38_right =
     fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? fsm38_out : 3'd0;
    assign incr39_left =
     fsm92_out == 10'd116 & go ? 1'd1 : 1'd0;
    assign incr39_right =
     fsm92_out == 10'd116 & go ? fsm39_out : 1'd0;
    assign incr4_left =
     fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go ? 3'd1 : 3'd0;
    assign incr4_right =
     fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go ? fsm4_out : 3'd0;
    assign incr40_left =
     fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? 3'd1 : 3'd0;
    assign incr40_right =
     fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? fsm40_out : 3'd0;
    assign incr41_left =
     fsm92_out == 10'd122 & go ? 1'd1 : 1'd0;
    assign incr41_right =
     fsm92_out == 10'd122 & go ? fsm41_out : 1'd0;
    assign incr42_left =
     fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? 3'd1 : 3'd0;
    assign incr42_right =
     fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? fsm42_out : 3'd0;
    assign incr43_left =
     fsm92_out == 10'd128 & go ? 1'd1 : 1'd0;
    assign incr43_right =
     fsm92_out == 10'd128 & go ? fsm43_out : 1'd0;
    assign incr44_left =
     fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? 3'd1 : 3'd0;
    assign incr44_right =
     fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? fsm44_out : 3'd0;
    assign incr45_left =
     fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign incr45_right =
     fsm92_out == 10'd134 & go ? fsm45_out : 1'd0;
    assign incr46_left =
     fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? 3'd1 : 3'd0;
    assign incr46_right =
     fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? fsm46_out : 3'd0;
    assign incr47_left =
     fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign incr47_right =
     fsm92_out == 10'd140 & go ? fsm47_out : 1'd0;
    assign incr48_left =
     fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? 3'd1 : 3'd0;
    assign incr48_right =
     fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? fsm48_out : 3'd0;
    assign incr49_left =
     fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign incr49_right =
     fsm92_out == 10'd146 & go ? fsm49_out : 1'd0;
    assign incr5_left =
     fsm92_out == 10'd14 & go ? 1'd1 : 1'd0;
    assign incr5_right =
     fsm92_out == 10'd14 & go ? fsm5_out : 1'd0;
    assign incr50_left =
     fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? 3'd1 : 3'd0;
    assign incr50_right =
     fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? fsm50_out : 3'd0;
    assign incr51_left =
     fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign incr51_right =
     fsm92_out == 10'd152 & go ? fsm51_out : 1'd0;
    assign incr52_left =
     fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? 3'd1 : 3'd0;
    assign incr52_right =
     fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? fsm52_out : 3'd0;
    assign incr53_left =
     fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign incr53_right =
     fsm92_out == 10'd158 & go ? fsm53_out : 1'd0;
    assign incr54_left =
     fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 3'd1 : 3'd0;
    assign incr54_right =
     fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? fsm54_out : 3'd0;
    assign incr55_left =
     fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign incr55_right =
     fsm92_out == 10'd164 & go ? fsm55_out : 1'd0;
    assign incr56_left =
     fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 3'd1 : 3'd0;
    assign incr56_right =
     fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? fsm56_out : 3'd0;
    assign incr57_left =
     fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign incr57_right =
     fsm92_out == 10'd170 & go ? fsm57_out : 1'd0;
    assign incr58_left =
     fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 3'd1 : 3'd0;
    assign incr58_right =
     fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? fsm58_out : 3'd0;
    assign incr59_left =
     fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign incr59_right =
     fsm92_out == 10'd176 & go ? fsm59_out : 1'd0;
    assign incr6_left =
     fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go ? 3'd1 : 3'd0;
    assign incr6_right =
     fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go ? fsm6_out : 3'd0;
    assign incr60_left =
     fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 3'd1 : 3'd0;
    assign incr60_right =
     fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? fsm60_out : 3'd0;
    assign incr61_left =
     fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign incr61_right =
     fsm92_out == 10'd182 & go ? fsm61_out : 1'd0;
    assign incr62_left =
     fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 3'd1 : 3'd0;
    assign incr62_right =
     fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? fsm62_out : 3'd0;
    assign incr63_left =
     fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign incr63_right =
     fsm92_out == 10'd188 & go ? fsm63_out : 1'd0;
    assign incr64_left =
     fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? 3'd1 : 3'd0;
    assign incr64_right =
     fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? fsm64_out : 3'd0;
    assign incr65_left =
     fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign incr65_right =
     fsm92_out == 10'd194 & go ? fsm65_out : 1'd0;
    assign incr66_left =
     fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? 3'd1 : 3'd0;
    assign incr66_right =
     fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? fsm66_out : 3'd0;
    assign incr67_left =
     fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign incr67_right =
     fsm92_out == 10'd200 & go ? fsm67_out : 1'd0;
    assign incr68_left =
     fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? 3'd1 : 3'd0;
    assign incr68_right =
     fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? fsm68_out : 3'd0;
    assign incr69_left =
     fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign incr69_right =
     fsm92_out == 10'd206 & go ? fsm69_out : 1'd0;
    assign incr7_left =
     fsm92_out == 10'd20 & go ? 1'd1 : 1'd0;
    assign incr7_right =
     fsm92_out == 10'd20 & go ? fsm7_out : 1'd0;
    assign incr70_left =
     fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? 3'd1 : 3'd0;
    assign incr70_right =
     fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? fsm70_out : 3'd0;
    assign incr71_left =
     fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign incr71_right =
     fsm92_out == 10'd212 & go ? fsm71_out : 1'd0;
    assign incr72_left =
     fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? 3'd1 : 3'd0;
    assign incr72_right =
     fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? fsm72_out : 3'd0;
    assign incr73_left =
     fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign incr73_right =
     fsm92_out == 10'd218 & go ? fsm73_out : 1'd0;
    assign incr74_left =
     fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? 3'd1 : 3'd0;
    assign incr74_right =
     fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? fsm74_out : 3'd0;
    assign incr75_left =
     fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign incr75_right =
     fsm92_out == 10'd224 & go ? fsm75_out : 1'd0;
    assign incr76_left =
     fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? 3'd1 : 3'd0;
    assign incr76_right =
     fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? fsm76_out : 3'd0;
    assign incr77_left =
     fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign incr77_right =
     fsm92_out == 10'd230 & go ? fsm77_out : 1'd0;
    assign incr78_left =
     fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? 3'd1 : 3'd0;
    assign incr78_right =
     fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? fsm78_out : 3'd0;
    assign incr79_left =
     fsm92_out == 10'd236 & go ? 1'd1 : 1'd0;
    assign incr79_right =
     fsm92_out == 10'd236 & go ? fsm79_out : 1'd0;
    assign incr8_left =
     fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go ? 3'd1 : 3'd0;
    assign incr8_right =
     fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go ? fsm8_out : 3'd0;
    assign incr80_left =
     fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? 3'd1 : 3'd0;
    assign incr80_right =
     fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? fsm80_out : 3'd0;
    assign incr81_left =
     fsm92_out == 10'd242 & go ? 1'd1 : 1'd0;
    assign incr81_right =
     fsm92_out == 10'd242 & go ? fsm81_out : 1'd0;
    assign incr82_left =
     fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? 3'd1 : 3'd0;
    assign incr82_right =
     fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? fsm82_out : 3'd0;
    assign incr83_left =
     fsm92_out == 10'd248 & go ? 1'd1 : 1'd0;
    assign incr83_right =
     fsm92_out == 10'd248 & go ? fsm83_out : 1'd0;
    assign incr84_left =
     fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? 3'd1 : 3'd0;
    assign incr84_right =
     fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? fsm84_out : 3'd0;
    assign incr85_left =
     fsm92_out == 10'd254 & go ? 1'd1 : 1'd0;
    assign incr85_right =
     fsm92_out == 10'd254 & go ? fsm85_out : 1'd0;
    assign incr86_left =
     fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go ? 3'd1 : 3'd0;
    assign incr86_right =
     fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go ? fsm86_out : 3'd0;
    assign incr87_left =
     fsm92_out == 10'd260 & go ? 1'd1 : 1'd0;
    assign incr87_right =
     fsm92_out == 10'd260 & go ? fsm87_out : 1'd0;
    assign incr88_left =
     fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go ? 3'd1 : 3'd0;
    assign incr88_right =
     fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go ? fsm88_out : 3'd0;
    assign incr89_left =
     fsm92_out == 10'd266 & go ? 1'd1 : 1'd0;
    assign incr89_right =
     fsm92_out == 10'd266 & go ? fsm89_out : 1'd0;
    assign incr9_left =
     fsm92_out == 10'd26 & go ? 1'd1 : 1'd0;
    assign incr9_right =
     fsm92_out == 10'd26 & go ? fsm9_out : 1'd0;
    assign incr90_left =
     fsm92_out >= 10'd267 & fsm92_out < 10'd272 & go ? 3'd1 : 3'd0;
    assign incr90_right =
     fsm92_out >= 10'd267 & fsm92_out < 10'd272 & go ? fsm90_out : 3'd0;
    assign incr91_left =
     fsm92_out == 10'd272 & go ? 1'd1 : 1'd0;
    assign incr91_right =
     fsm92_out == 10'd272 & go ? fsm91_out : 1'd0;
    assign incr92_left =
     go ? 10'd1 : 10'd0;
    assign incr92_right =
     go ? fsm92_out : 10'd0;
    assign l0_add_left =
     fsm0_out < 1'd1 & fsm92_out == 10'd1 & go | fsm2_out < 3'd1 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go ? 5'd1 : 5'd0;
    assign l0_add_right =
     fsm0_out < 1'd1 & fsm92_out == 10'd1 & go | fsm2_out < 3'd1 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go ? l0_idx_out : 5'd0;
    assign l0_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l0_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm0_out < 1'd1 & fsm92_out == 10'd1 & go | fsm2_out < 3'd1 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go ? l0_add_out : 5'd0;
    assign l0_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm0_out < 1'd1 & fsm92_out == 10'd1 & go | fsm2_out < 3'd1 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go ? 1'd1 : 1'd0;
    assign l10_add_left =
     fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? 5'd1 : 5'd0;
    assign l10_add_right =
     fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? l10_idx_out : 5'd0;
    assign l10_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l10_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? l10_add_out : 5'd0;
    assign l10_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? 1'd1 : 1'd0;
    assign l11_add_left =
     fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? 5'd1 : 5'd0;
    assign l11_add_right =
     fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? l11_idx_out : 5'd0;
    assign l11_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l11_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? l11_add_out : 5'd0;
    assign l11_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? 1'd1 : 1'd0;
    assign l12_add_left =
     fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 5'd1 : 5'd0;
    assign l12_add_right =
     fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? l12_idx_out : 5'd0;
    assign l12_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l12_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? l12_add_out : 5'd0;
    assign l12_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 1'd1 : 1'd0;
    assign l13_add_left =
     fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 5'd1 : 5'd0;
    assign l13_add_right =
     fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? l13_idx_out : 5'd0;
    assign l13_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l13_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? l13_add_out : 5'd0;
    assign l13_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 1'd1 : 1'd0;
    assign l14_add_left =
     fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd1 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 5'd1 : 5'd0;
    assign l14_add_right =
     fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd1 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? l14_idx_out : 5'd0;
    assign l14_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l14_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd1 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? l14_add_out : 5'd0;
    assign l14_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd1 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 1'd1 : 1'd0;
    assign l15_add_left =
     fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd1 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd1 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 5'd1 : 5'd0;
    assign l15_add_right =
     fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd1 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd1 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? l15_idx_out : 5'd0;
    assign l15_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l15_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd1 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd1 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? l15_add_out : 5'd0;
    assign l15_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd1 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd1 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign l1_add_left =
     fsm2_out < 3'd1 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go ? 5'd1 : 5'd0;
    assign l1_add_right =
     fsm2_out < 3'd1 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go ? l1_idx_out : 5'd0;
    assign l1_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l1_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm2_out < 3'd1 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go ? l1_add_out : 5'd0;
    assign l1_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm2_out < 3'd1 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go ? 1'd1 : 1'd0;
    assign l2_add_left =
     fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? 5'd1 : 5'd0;
    assign l2_add_right =
     fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? l2_idx_out : 5'd0;
    assign l2_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l2_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? l2_add_out : 5'd0;
    assign l2_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? 1'd1 : 1'd0;
    assign l3_add_left =
     fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? 5'd1 : 5'd0;
    assign l3_add_right =
     fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? l3_idx_out : 5'd0;
    assign l3_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l3_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? l3_add_out : 5'd0;
    assign l3_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? 1'd1 : 1'd0;
    assign l4_add_left =
     fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? 5'd1 : 5'd0;
    assign l4_add_right =
     fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? l4_idx_out : 5'd0;
    assign l4_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l4_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? l4_add_out : 5'd0;
    assign l4_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? 1'd1 : 1'd0;
    assign l5_add_left =
     fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? 5'd1 : 5'd0;
    assign l5_add_right =
     fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? l5_idx_out : 5'd0;
    assign l5_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l5_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? l5_add_out : 5'd0;
    assign l5_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? 1'd1 : 1'd0;
    assign l6_add_left =
     fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? 5'd1 : 5'd0;
    assign l6_add_right =
     fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? l6_idx_out : 5'd0;
    assign l6_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l6_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? l6_add_out : 5'd0;
    assign l6_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? 1'd1 : 1'd0;
    assign l7_add_left =
     fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? 5'd1 : 5'd0;
    assign l7_add_right =
     fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? l7_idx_out : 5'd0;
    assign l7_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l7_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? l7_add_out : 5'd0;
    assign l7_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? 1'd1 : 1'd0;
    assign l8_add_left =
     fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? 5'd1 : 5'd0;
    assign l8_add_right =
     fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? l8_idx_out : 5'd0;
    assign l8_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l8_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? l8_add_out : 5'd0;
    assign l8_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? 1'd1 : 1'd0;
    assign l9_add_left =
     fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? 5'd1 : 5'd0;
    assign l9_add_right =
     fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? l9_idx_out : 5'd0;
    assign l9_idx_clk =
     1'b1 ? clk : 1'd0;
    assign l9_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? l9_add_out : 5'd0;
    assign l9_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? 1'd1 : 1'd0;
    assign left_0_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_0_in =
     fsm1_out < 1'd1 & fsm92_out == 10'd2 & go | fsm3_out < 1'd1 & fsm92_out == 10'd8 & go | fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go ? l0_read_data : 32'd0;
    assign left_0_0_write_en =
     fsm1_out < 1'd1 & fsm92_out == 10'd2 & go | fsm3_out < 1'd1 & fsm92_out == 10'd8 & go | fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go ? 1'd1 : 1'd0;
    assign left_0_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_1_in =
     fsm3_out < 1'd1 & fsm92_out == 10'd8 & go | fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go ? left_0_0_out : 32'd0;
    assign left_0_1_write_en =
     fsm3_out < 1'd1 & fsm92_out == 10'd8 & go | fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go ? 1'd1 : 1'd0;
    assign left_0_10_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_10_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? left_0_9_out : 32'd0;
    assign left_0_10_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign left_0_11_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_11_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? left_0_10_out : 32'd0;
    assign left_0_11_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign left_0_12_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_12_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? left_0_11_out : 32'd0;
    assign left_0_12_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign left_0_13_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_13_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? left_0_12_out : 32'd0;
    assign left_0_13_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign left_0_14_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_14_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? left_0_13_out : 32'd0;
    assign left_0_14_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign left_0_15_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_15_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? left_0_14_out : 32'd0;
    assign left_0_15_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign left_0_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_2_in =
     fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go ? left_0_1_out : 32'd0;
    assign left_0_2_write_en =
     fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go ? 1'd1 : 1'd0;
    assign left_0_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_3_in =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? left_0_2_out : 32'd0;
    assign left_0_3_write_en =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? 1'd1 : 1'd0;
    assign left_0_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_4_in =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? left_0_3_out : 32'd0;
    assign left_0_4_write_en =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? 1'd1 : 1'd0;
    assign left_0_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_5_in =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? left_0_4_out : 32'd0;
    assign left_0_5_write_en =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? 1'd1 : 1'd0;
    assign left_0_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_6_in =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? left_0_5_out : 32'd0;
    assign left_0_6_write_en =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? 1'd1 : 1'd0;
    assign left_0_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_7_in =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? left_0_6_out : 32'd0;
    assign left_0_7_write_en =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign left_0_8_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_8_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? left_0_7_out : 32'd0;
    assign left_0_8_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign left_0_9_clk =
     1'b1 ? clk : 1'd0;
    assign left_0_9_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? left_0_8_out : 32'd0;
    assign left_0_9_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign left_10_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_10_0_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? l10_read_data : 32'd0;
    assign left_10_0_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign left_10_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_10_1_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? left_10_0_out : 32'd0;
    assign left_10_1_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign left_10_10_clk =
     1'b1 ? clk : 1'd0;
    assign left_10_10_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? left_10_9_out : 32'd0;
    assign left_10_10_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign left_10_11_clk =
     1'b1 ? clk : 1'd0;
    assign left_10_11_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? left_10_10_out : 32'd0;
    assign left_10_11_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign left_10_12_clk =
     1'b1 ? clk : 1'd0;
    assign left_10_12_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? left_10_11_out : 32'd0;
    assign left_10_12_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign left_10_13_clk =
     1'b1 ? clk : 1'd0;
    assign left_10_13_in =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? left_10_12_out : 32'd0;
    assign left_10_13_write_en =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign left_10_14_clk =
     1'b1 ? clk : 1'd0;
    assign left_10_14_in =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? left_10_13_out : 32'd0;
    assign left_10_14_write_en =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? 1'd1 : 1'd0;
    assign left_10_15_clk =
     1'b1 ? clk : 1'd0;
    assign left_10_15_in =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? left_10_14_out : 32'd0;
    assign left_10_15_write_en =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? 1'd1 : 1'd0;
    assign left_10_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_10_2_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? left_10_1_out : 32'd0;
    assign left_10_2_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign left_10_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_10_3_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? left_10_2_out : 32'd0;
    assign left_10_3_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign left_10_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_10_4_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? left_10_3_out : 32'd0;
    assign left_10_4_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign left_10_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_10_5_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? left_10_4_out : 32'd0;
    assign left_10_5_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign left_10_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_10_6_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? left_10_5_out : 32'd0;
    assign left_10_6_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign left_10_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_10_7_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? left_10_6_out : 32'd0;
    assign left_10_7_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign left_10_8_clk =
     1'b1 ? clk : 1'd0;
    assign left_10_8_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? left_10_7_out : 32'd0;
    assign left_10_8_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign left_10_9_clk =
     1'b1 ? clk : 1'd0;
    assign left_10_9_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? left_10_8_out : 32'd0;
    assign left_10_9_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign left_11_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_11_0_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? l11_read_data : 32'd0;
    assign left_11_0_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign left_11_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_11_1_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? left_11_0_out : 32'd0;
    assign left_11_1_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign left_11_10_clk =
     1'b1 ? clk : 1'd0;
    assign left_11_10_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? left_11_9_out : 32'd0;
    assign left_11_10_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign left_11_11_clk =
     1'b1 ? clk : 1'd0;
    assign left_11_11_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? left_11_10_out : 32'd0;
    assign left_11_11_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign left_11_12_clk =
     1'b1 ? clk : 1'd0;
    assign left_11_12_in =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? left_11_11_out : 32'd0;
    assign left_11_12_write_en =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign left_11_13_clk =
     1'b1 ? clk : 1'd0;
    assign left_11_13_in =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? left_11_12_out : 32'd0;
    assign left_11_13_write_en =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? 1'd1 : 1'd0;
    assign left_11_14_clk =
     1'b1 ? clk : 1'd0;
    assign left_11_14_in =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? left_11_13_out : 32'd0;
    assign left_11_14_write_en =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? 1'd1 : 1'd0;
    assign left_11_15_clk =
     1'b1 ? clk : 1'd0;
    assign left_11_15_in =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? left_11_14_out : 32'd0;
    assign left_11_15_write_en =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? 1'd1 : 1'd0;
    assign left_11_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_11_2_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? left_11_1_out : 32'd0;
    assign left_11_2_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign left_11_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_11_3_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? left_11_2_out : 32'd0;
    assign left_11_3_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign left_11_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_11_4_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? left_11_3_out : 32'd0;
    assign left_11_4_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign left_11_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_11_5_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? left_11_4_out : 32'd0;
    assign left_11_5_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign left_11_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_11_6_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? left_11_5_out : 32'd0;
    assign left_11_6_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign left_11_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_11_7_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? left_11_6_out : 32'd0;
    assign left_11_7_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign left_11_8_clk =
     1'b1 ? clk : 1'd0;
    assign left_11_8_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? left_11_7_out : 32'd0;
    assign left_11_8_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign left_11_9_clk =
     1'b1 ? clk : 1'd0;
    assign left_11_9_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? left_11_8_out : 32'd0;
    assign left_11_9_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign left_12_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_12_0_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? l12_read_data : 32'd0;
    assign left_12_0_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign left_12_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_12_1_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? left_12_0_out : 32'd0;
    assign left_12_1_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign left_12_10_clk =
     1'b1 ? clk : 1'd0;
    assign left_12_10_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? left_12_9_out : 32'd0;
    assign left_12_10_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign left_12_11_clk =
     1'b1 ? clk : 1'd0;
    assign left_12_11_in =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? left_12_10_out : 32'd0;
    assign left_12_11_write_en =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign left_12_12_clk =
     1'b1 ? clk : 1'd0;
    assign left_12_12_in =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? left_12_11_out : 32'd0;
    assign left_12_12_write_en =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? 1'd1 : 1'd0;
    assign left_12_13_clk =
     1'b1 ? clk : 1'd0;
    assign left_12_13_in =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? left_12_12_out : 32'd0;
    assign left_12_13_write_en =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? 1'd1 : 1'd0;
    assign left_12_14_clk =
     1'b1 ? clk : 1'd0;
    assign left_12_14_in =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? left_12_13_out : 32'd0;
    assign left_12_14_write_en =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? 1'd1 : 1'd0;
    assign left_12_15_clk =
     1'b1 ? clk : 1'd0;
    assign left_12_15_in =
     fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go ? left_12_14_out : 32'd0;
    assign left_12_15_write_en =
     fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go ? 1'd1 : 1'd0;
    assign left_12_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_12_2_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? left_12_1_out : 32'd0;
    assign left_12_2_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign left_12_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_12_3_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? left_12_2_out : 32'd0;
    assign left_12_3_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign left_12_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_12_4_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? left_12_3_out : 32'd0;
    assign left_12_4_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign left_12_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_12_5_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? left_12_4_out : 32'd0;
    assign left_12_5_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign left_12_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_12_6_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? left_12_5_out : 32'd0;
    assign left_12_6_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign left_12_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_12_7_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? left_12_6_out : 32'd0;
    assign left_12_7_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign left_12_8_clk =
     1'b1 ? clk : 1'd0;
    assign left_12_8_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? left_12_7_out : 32'd0;
    assign left_12_8_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign left_12_9_clk =
     1'b1 ? clk : 1'd0;
    assign left_12_9_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? left_12_8_out : 32'd0;
    assign left_12_9_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign left_13_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_13_0_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? l13_read_data : 32'd0;
    assign left_13_0_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign left_13_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_13_1_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? left_13_0_out : 32'd0;
    assign left_13_1_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign left_13_10_clk =
     1'b1 ? clk : 1'd0;
    assign left_13_10_in =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? left_13_9_out : 32'd0;
    assign left_13_10_write_en =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign left_13_11_clk =
     1'b1 ? clk : 1'd0;
    assign left_13_11_in =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? left_13_10_out : 32'd0;
    assign left_13_11_write_en =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? 1'd1 : 1'd0;
    assign left_13_12_clk =
     1'b1 ? clk : 1'd0;
    assign left_13_12_in =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? left_13_11_out : 32'd0;
    assign left_13_12_write_en =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? 1'd1 : 1'd0;
    assign left_13_13_clk =
     1'b1 ? clk : 1'd0;
    assign left_13_13_in =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? left_13_12_out : 32'd0;
    assign left_13_13_write_en =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? 1'd1 : 1'd0;
    assign left_13_14_clk =
     1'b1 ? clk : 1'd0;
    assign left_13_14_in =
     fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go ? left_13_13_out : 32'd0;
    assign left_13_14_write_en =
     fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go ? 1'd1 : 1'd0;
    assign left_13_15_clk =
     1'b1 ? clk : 1'd0;
    assign left_13_15_in =
     fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go ? left_13_14_out : 32'd0;
    assign left_13_15_write_en =
     fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go ? 1'd1 : 1'd0;
    assign left_13_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_13_2_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? left_13_1_out : 32'd0;
    assign left_13_2_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign left_13_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_13_3_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? left_13_2_out : 32'd0;
    assign left_13_3_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign left_13_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_13_4_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? left_13_3_out : 32'd0;
    assign left_13_4_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign left_13_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_13_5_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? left_13_4_out : 32'd0;
    assign left_13_5_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign left_13_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_13_6_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? left_13_5_out : 32'd0;
    assign left_13_6_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign left_13_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_13_7_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? left_13_6_out : 32'd0;
    assign left_13_7_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign left_13_8_clk =
     1'b1 ? clk : 1'd0;
    assign left_13_8_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? left_13_7_out : 32'd0;
    assign left_13_8_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign left_13_9_clk =
     1'b1 ? clk : 1'd0;
    assign left_13_9_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? left_13_8_out : 32'd0;
    assign left_13_9_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign left_14_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_14_0_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? l14_read_data : 32'd0;
    assign left_14_0_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign left_14_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_14_1_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? left_14_0_out : 32'd0;
    assign left_14_1_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign left_14_10_clk =
     1'b1 ? clk : 1'd0;
    assign left_14_10_in =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? left_14_9_out : 32'd0;
    assign left_14_10_write_en =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? 1'd1 : 1'd0;
    assign left_14_11_clk =
     1'b1 ? clk : 1'd0;
    assign left_14_11_in =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? left_14_10_out : 32'd0;
    assign left_14_11_write_en =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? 1'd1 : 1'd0;
    assign left_14_12_clk =
     1'b1 ? clk : 1'd0;
    assign left_14_12_in =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? left_14_11_out : 32'd0;
    assign left_14_12_write_en =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? 1'd1 : 1'd0;
    assign left_14_13_clk =
     1'b1 ? clk : 1'd0;
    assign left_14_13_in =
     fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go ? left_14_12_out : 32'd0;
    assign left_14_13_write_en =
     fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go ? 1'd1 : 1'd0;
    assign left_14_14_clk =
     1'b1 ? clk : 1'd0;
    assign left_14_14_in =
     fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go ? left_14_13_out : 32'd0;
    assign left_14_14_write_en =
     fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go ? 1'd1 : 1'd0;
    assign left_14_15_clk =
     1'b1 ? clk : 1'd0;
    assign left_14_15_in =
     fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go | fsm89_out < 1'd1 & fsm92_out == 10'd266 & go ? left_14_14_out : 32'd0;
    assign left_14_15_write_en =
     fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go | fsm89_out < 1'd1 & fsm92_out == 10'd266 & go ? 1'd1 : 1'd0;
    assign left_14_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_14_2_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? left_14_1_out : 32'd0;
    assign left_14_2_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign left_14_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_14_3_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? left_14_2_out : 32'd0;
    assign left_14_3_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign left_14_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_14_4_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? left_14_3_out : 32'd0;
    assign left_14_4_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign left_14_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_14_5_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? left_14_4_out : 32'd0;
    assign left_14_5_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign left_14_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_14_6_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? left_14_5_out : 32'd0;
    assign left_14_6_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign left_14_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_14_7_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? left_14_6_out : 32'd0;
    assign left_14_7_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign left_14_8_clk =
     1'b1 ? clk : 1'd0;
    assign left_14_8_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? left_14_7_out : 32'd0;
    assign left_14_8_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign left_14_9_clk =
     1'b1 ? clk : 1'd0;
    assign left_14_9_in =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? left_14_8_out : 32'd0;
    assign left_14_9_write_en =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign left_15_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_15_0_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? l15_read_data : 32'd0;
    assign left_15_0_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign left_15_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_15_1_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? left_15_0_out : 32'd0;
    assign left_15_1_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign left_15_10_clk =
     1'b1 ? clk : 1'd0;
    assign left_15_10_in =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? left_15_9_out : 32'd0;
    assign left_15_10_write_en =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? 1'd1 : 1'd0;
    assign left_15_11_clk =
     1'b1 ? clk : 1'd0;
    assign left_15_11_in =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? left_15_10_out : 32'd0;
    assign left_15_11_write_en =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? 1'd1 : 1'd0;
    assign left_15_12_clk =
     1'b1 ? clk : 1'd0;
    assign left_15_12_in =
     fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go ? left_15_11_out : 32'd0;
    assign left_15_12_write_en =
     fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go ? 1'd1 : 1'd0;
    assign left_15_13_clk =
     1'b1 ? clk : 1'd0;
    assign left_15_13_in =
     fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go ? left_15_12_out : 32'd0;
    assign left_15_13_write_en =
     fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go ? 1'd1 : 1'd0;
    assign left_15_14_clk =
     1'b1 ? clk : 1'd0;
    assign left_15_14_in =
     fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go | fsm89_out < 1'd1 & fsm92_out == 10'd266 & go ? left_15_13_out : 32'd0;
    assign left_15_14_write_en =
     fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go | fsm89_out < 1'd1 & fsm92_out == 10'd266 & go ? 1'd1 : 1'd0;
    assign left_15_15_clk =
     1'b1 ? clk : 1'd0;
    assign left_15_15_in =
     fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go | fsm89_out < 1'd1 & fsm92_out == 10'd266 & go | fsm91_out < 1'd1 & fsm92_out == 10'd272 & go ? left_15_14_out : 32'd0;
    assign left_15_15_write_en =
     fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go | fsm89_out < 1'd1 & fsm92_out == 10'd266 & go | fsm91_out < 1'd1 & fsm92_out == 10'd272 & go ? 1'd1 : 1'd0;
    assign left_15_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_15_2_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? left_15_1_out : 32'd0;
    assign left_15_2_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign left_15_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_15_3_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? left_15_2_out : 32'd0;
    assign left_15_3_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign left_15_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_15_4_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? left_15_3_out : 32'd0;
    assign left_15_4_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign left_15_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_15_5_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? left_15_4_out : 32'd0;
    assign left_15_5_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign left_15_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_15_6_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? left_15_5_out : 32'd0;
    assign left_15_6_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign left_15_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_15_7_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? left_15_6_out : 32'd0;
    assign left_15_7_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign left_15_8_clk =
     1'b1 ? clk : 1'd0;
    assign left_15_8_in =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? left_15_7_out : 32'd0;
    assign left_15_8_write_en =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign left_15_9_clk =
     1'b1 ? clk : 1'd0;
    assign left_15_9_in =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? left_15_8_out : 32'd0;
    assign left_15_9_write_en =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? 1'd1 : 1'd0;
    assign left_1_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_0_in =
     fsm3_out < 1'd1 & fsm92_out == 10'd8 & go | fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go ? l1_read_data : 32'd0;
    assign left_1_0_write_en =
     fsm3_out < 1'd1 & fsm92_out == 10'd8 & go | fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go ? 1'd1 : 1'd0;
    assign left_1_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_1_in =
     fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go ? left_1_0_out : 32'd0;
    assign left_1_1_write_en =
     fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go ? 1'd1 : 1'd0;
    assign left_1_10_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_10_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? left_1_9_out : 32'd0;
    assign left_1_10_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign left_1_11_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_11_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? left_1_10_out : 32'd0;
    assign left_1_11_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign left_1_12_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_12_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? left_1_11_out : 32'd0;
    assign left_1_12_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign left_1_13_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_13_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? left_1_12_out : 32'd0;
    assign left_1_13_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign left_1_14_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_14_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? left_1_13_out : 32'd0;
    assign left_1_14_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign left_1_15_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_15_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? left_1_14_out : 32'd0;
    assign left_1_15_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign left_1_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_2_in =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? left_1_1_out : 32'd0;
    assign left_1_2_write_en =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? 1'd1 : 1'd0;
    assign left_1_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_3_in =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? left_1_2_out : 32'd0;
    assign left_1_3_write_en =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? 1'd1 : 1'd0;
    assign left_1_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_4_in =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? left_1_3_out : 32'd0;
    assign left_1_4_write_en =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? 1'd1 : 1'd0;
    assign left_1_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_5_in =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? left_1_4_out : 32'd0;
    assign left_1_5_write_en =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? 1'd1 : 1'd0;
    assign left_1_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_6_in =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? left_1_5_out : 32'd0;
    assign left_1_6_write_en =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign left_1_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_7_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? left_1_6_out : 32'd0;
    assign left_1_7_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign left_1_8_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_8_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? left_1_7_out : 32'd0;
    assign left_1_8_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign left_1_9_clk =
     1'b1 ? clk : 1'd0;
    assign left_1_9_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? left_1_8_out : 32'd0;
    assign left_1_9_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign left_2_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_0_in =
     fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go ? l2_read_data : 32'd0;
    assign left_2_0_write_en =
     fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go ? 1'd1 : 1'd0;
    assign left_2_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_1_in =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? left_2_0_out : 32'd0;
    assign left_2_1_write_en =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? 1'd1 : 1'd0;
    assign left_2_10_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_10_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? left_2_9_out : 32'd0;
    assign left_2_10_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign left_2_11_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_11_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? left_2_10_out : 32'd0;
    assign left_2_11_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign left_2_12_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_12_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? left_2_11_out : 32'd0;
    assign left_2_12_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign left_2_13_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_13_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? left_2_12_out : 32'd0;
    assign left_2_13_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign left_2_14_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_14_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? left_2_13_out : 32'd0;
    assign left_2_14_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign left_2_15_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_15_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? left_2_14_out : 32'd0;
    assign left_2_15_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign left_2_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_2_in =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? left_2_1_out : 32'd0;
    assign left_2_2_write_en =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? 1'd1 : 1'd0;
    assign left_2_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_3_in =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? left_2_2_out : 32'd0;
    assign left_2_3_write_en =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? 1'd1 : 1'd0;
    assign left_2_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_4_in =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? left_2_3_out : 32'd0;
    assign left_2_4_write_en =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? 1'd1 : 1'd0;
    assign left_2_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_5_in =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? left_2_4_out : 32'd0;
    assign left_2_5_write_en =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign left_2_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_6_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? left_2_5_out : 32'd0;
    assign left_2_6_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign left_2_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_7_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? left_2_6_out : 32'd0;
    assign left_2_7_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign left_2_8_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_8_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? left_2_7_out : 32'd0;
    assign left_2_8_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign left_2_9_clk =
     1'b1 ? clk : 1'd0;
    assign left_2_9_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? left_2_8_out : 32'd0;
    assign left_2_9_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign left_3_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_0_in =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? l3_read_data : 32'd0;
    assign left_3_0_write_en =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? 1'd1 : 1'd0;
    assign left_3_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_1_in =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? left_3_0_out : 32'd0;
    assign left_3_1_write_en =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? 1'd1 : 1'd0;
    assign left_3_10_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_10_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? left_3_9_out : 32'd0;
    assign left_3_10_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign left_3_11_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_11_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? left_3_10_out : 32'd0;
    assign left_3_11_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign left_3_12_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_12_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? left_3_11_out : 32'd0;
    assign left_3_12_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign left_3_13_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_13_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? left_3_12_out : 32'd0;
    assign left_3_13_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign left_3_14_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_14_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? left_3_13_out : 32'd0;
    assign left_3_14_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign left_3_15_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_15_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? left_3_14_out : 32'd0;
    assign left_3_15_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign left_3_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_2_in =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? left_3_1_out : 32'd0;
    assign left_3_2_write_en =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? 1'd1 : 1'd0;
    assign left_3_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_3_in =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? left_3_2_out : 32'd0;
    assign left_3_3_write_en =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? 1'd1 : 1'd0;
    assign left_3_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_4_in =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? left_3_3_out : 32'd0;
    assign left_3_4_write_en =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign left_3_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_5_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? left_3_4_out : 32'd0;
    assign left_3_5_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign left_3_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_6_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? left_3_5_out : 32'd0;
    assign left_3_6_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign left_3_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_7_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? left_3_6_out : 32'd0;
    assign left_3_7_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign left_3_8_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_8_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? left_3_7_out : 32'd0;
    assign left_3_8_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign left_3_9_clk =
     1'b1 ? clk : 1'd0;
    assign left_3_9_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? left_3_8_out : 32'd0;
    assign left_3_9_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign left_4_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_0_in =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? l4_read_data : 32'd0;
    assign left_4_0_write_en =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? 1'd1 : 1'd0;
    assign left_4_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_1_in =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? left_4_0_out : 32'd0;
    assign left_4_1_write_en =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? 1'd1 : 1'd0;
    assign left_4_10_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_10_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? left_4_9_out : 32'd0;
    assign left_4_10_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign left_4_11_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_11_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? left_4_10_out : 32'd0;
    assign left_4_11_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign left_4_12_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_12_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? left_4_11_out : 32'd0;
    assign left_4_12_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign left_4_13_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_13_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? left_4_12_out : 32'd0;
    assign left_4_13_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign left_4_14_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_14_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? left_4_13_out : 32'd0;
    assign left_4_14_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign left_4_15_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_15_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? left_4_14_out : 32'd0;
    assign left_4_15_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign left_4_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_2_in =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? left_4_1_out : 32'd0;
    assign left_4_2_write_en =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? 1'd1 : 1'd0;
    assign left_4_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_3_in =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? left_4_2_out : 32'd0;
    assign left_4_3_write_en =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign left_4_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_4_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? left_4_3_out : 32'd0;
    assign left_4_4_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign left_4_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_5_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? left_4_4_out : 32'd0;
    assign left_4_5_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign left_4_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_6_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? left_4_5_out : 32'd0;
    assign left_4_6_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign left_4_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_7_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? left_4_6_out : 32'd0;
    assign left_4_7_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign left_4_8_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_8_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? left_4_7_out : 32'd0;
    assign left_4_8_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign left_4_9_clk =
     1'b1 ? clk : 1'd0;
    assign left_4_9_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? left_4_8_out : 32'd0;
    assign left_4_9_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign left_5_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_0_in =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? l5_read_data : 32'd0;
    assign left_5_0_write_en =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? 1'd1 : 1'd0;
    assign left_5_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_1_in =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? left_5_0_out : 32'd0;
    assign left_5_1_write_en =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? 1'd1 : 1'd0;
    assign left_5_10_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_10_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? left_5_9_out : 32'd0;
    assign left_5_10_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign left_5_11_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_11_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? left_5_10_out : 32'd0;
    assign left_5_11_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign left_5_12_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_12_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? left_5_11_out : 32'd0;
    assign left_5_12_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign left_5_13_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_13_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? left_5_12_out : 32'd0;
    assign left_5_13_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign left_5_14_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_14_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? left_5_13_out : 32'd0;
    assign left_5_14_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign left_5_15_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_15_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? left_5_14_out : 32'd0;
    assign left_5_15_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign left_5_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_2_in =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? left_5_1_out : 32'd0;
    assign left_5_2_write_en =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign left_5_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_3_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? left_5_2_out : 32'd0;
    assign left_5_3_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign left_5_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_4_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? left_5_3_out : 32'd0;
    assign left_5_4_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign left_5_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_5_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? left_5_4_out : 32'd0;
    assign left_5_5_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign left_5_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_6_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? left_5_5_out : 32'd0;
    assign left_5_6_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign left_5_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_7_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? left_5_6_out : 32'd0;
    assign left_5_7_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign left_5_8_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_8_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? left_5_7_out : 32'd0;
    assign left_5_8_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign left_5_9_clk =
     1'b1 ? clk : 1'd0;
    assign left_5_9_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? left_5_8_out : 32'd0;
    assign left_5_9_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign left_6_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_0_in =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? l6_read_data : 32'd0;
    assign left_6_0_write_en =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? 1'd1 : 1'd0;
    assign left_6_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_1_in =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? left_6_0_out : 32'd0;
    assign left_6_1_write_en =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign left_6_10_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_10_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? left_6_9_out : 32'd0;
    assign left_6_10_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign left_6_11_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_11_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? left_6_10_out : 32'd0;
    assign left_6_11_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign left_6_12_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_12_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? left_6_11_out : 32'd0;
    assign left_6_12_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign left_6_13_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_13_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? left_6_12_out : 32'd0;
    assign left_6_13_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign left_6_14_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_14_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? left_6_13_out : 32'd0;
    assign left_6_14_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign left_6_15_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_15_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? left_6_14_out : 32'd0;
    assign left_6_15_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign left_6_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_2_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? left_6_1_out : 32'd0;
    assign left_6_2_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign left_6_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_3_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? left_6_2_out : 32'd0;
    assign left_6_3_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign left_6_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_4_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? left_6_3_out : 32'd0;
    assign left_6_4_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign left_6_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_5_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? left_6_4_out : 32'd0;
    assign left_6_5_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign left_6_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_6_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? left_6_5_out : 32'd0;
    assign left_6_6_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign left_6_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_7_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? left_6_6_out : 32'd0;
    assign left_6_7_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign left_6_8_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_8_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? left_6_7_out : 32'd0;
    assign left_6_8_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign left_6_9_clk =
     1'b1 ? clk : 1'd0;
    assign left_6_9_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? left_6_8_out : 32'd0;
    assign left_6_9_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign left_7_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_0_in =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? l7_read_data : 32'd0;
    assign left_7_0_write_en =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign left_7_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_1_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? left_7_0_out : 32'd0;
    assign left_7_1_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign left_7_10_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_10_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? left_7_9_out : 32'd0;
    assign left_7_10_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign left_7_11_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_11_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? left_7_10_out : 32'd0;
    assign left_7_11_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign left_7_12_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_12_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? left_7_11_out : 32'd0;
    assign left_7_12_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign left_7_13_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_13_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? left_7_12_out : 32'd0;
    assign left_7_13_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign left_7_14_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_14_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? left_7_13_out : 32'd0;
    assign left_7_14_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign left_7_15_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_15_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? left_7_14_out : 32'd0;
    assign left_7_15_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign left_7_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_2_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? left_7_1_out : 32'd0;
    assign left_7_2_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign left_7_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_3_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? left_7_2_out : 32'd0;
    assign left_7_3_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign left_7_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_4_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? left_7_3_out : 32'd0;
    assign left_7_4_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign left_7_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_5_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? left_7_4_out : 32'd0;
    assign left_7_5_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign left_7_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_6_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? left_7_5_out : 32'd0;
    assign left_7_6_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign left_7_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_7_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? left_7_6_out : 32'd0;
    assign left_7_7_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign left_7_8_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_8_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? left_7_7_out : 32'd0;
    assign left_7_8_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign left_7_9_clk =
     1'b1 ? clk : 1'd0;
    assign left_7_9_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? left_7_8_out : 32'd0;
    assign left_7_9_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign left_8_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_8_0_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? l8_read_data : 32'd0;
    assign left_8_0_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign left_8_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_8_1_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? left_8_0_out : 32'd0;
    assign left_8_1_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign left_8_10_clk =
     1'b1 ? clk : 1'd0;
    assign left_8_10_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? left_8_9_out : 32'd0;
    assign left_8_10_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign left_8_11_clk =
     1'b1 ? clk : 1'd0;
    assign left_8_11_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? left_8_10_out : 32'd0;
    assign left_8_11_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign left_8_12_clk =
     1'b1 ? clk : 1'd0;
    assign left_8_12_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? left_8_11_out : 32'd0;
    assign left_8_12_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign left_8_13_clk =
     1'b1 ? clk : 1'd0;
    assign left_8_13_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? left_8_12_out : 32'd0;
    assign left_8_13_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign left_8_14_clk =
     1'b1 ? clk : 1'd0;
    assign left_8_14_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? left_8_13_out : 32'd0;
    assign left_8_14_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign left_8_15_clk =
     1'b1 ? clk : 1'd0;
    assign left_8_15_in =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? left_8_14_out : 32'd0;
    assign left_8_15_write_en =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign left_8_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_8_2_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? left_8_1_out : 32'd0;
    assign left_8_2_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign left_8_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_8_3_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? left_8_2_out : 32'd0;
    assign left_8_3_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign left_8_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_8_4_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? left_8_3_out : 32'd0;
    assign left_8_4_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign left_8_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_8_5_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? left_8_4_out : 32'd0;
    assign left_8_5_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign left_8_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_8_6_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? left_8_5_out : 32'd0;
    assign left_8_6_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign left_8_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_8_7_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? left_8_6_out : 32'd0;
    assign left_8_7_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign left_8_8_clk =
     1'b1 ? clk : 1'd0;
    assign left_8_8_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? left_8_7_out : 32'd0;
    assign left_8_8_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign left_8_9_clk =
     1'b1 ? clk : 1'd0;
    assign left_8_9_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? left_8_8_out : 32'd0;
    assign left_8_9_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign left_9_0_clk =
     1'b1 ? clk : 1'd0;
    assign left_9_0_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? l9_read_data : 32'd0;
    assign left_9_0_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign left_9_1_clk =
     1'b1 ? clk : 1'd0;
    assign left_9_1_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? left_9_0_out : 32'd0;
    assign left_9_1_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign left_9_10_clk =
     1'b1 ? clk : 1'd0;
    assign left_9_10_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? left_9_9_out : 32'd0;
    assign left_9_10_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign left_9_11_clk =
     1'b1 ? clk : 1'd0;
    assign left_9_11_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? left_9_10_out : 32'd0;
    assign left_9_11_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign left_9_12_clk =
     1'b1 ? clk : 1'd0;
    assign left_9_12_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? left_9_11_out : 32'd0;
    assign left_9_12_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign left_9_13_clk =
     1'b1 ? clk : 1'd0;
    assign left_9_13_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? left_9_12_out : 32'd0;
    assign left_9_13_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign left_9_14_clk =
     1'b1 ? clk : 1'd0;
    assign left_9_14_in =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? left_9_13_out : 32'd0;
    assign left_9_14_write_en =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign left_9_15_clk =
     1'b1 ? clk : 1'd0;
    assign left_9_15_in =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? left_9_14_out : 32'd0;
    assign left_9_15_write_en =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? 1'd1 : 1'd0;
    assign left_9_2_clk =
     1'b1 ? clk : 1'd0;
    assign left_9_2_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? left_9_1_out : 32'd0;
    assign left_9_2_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign left_9_3_clk =
     1'b1 ? clk : 1'd0;
    assign left_9_3_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? left_9_2_out : 32'd0;
    assign left_9_3_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign left_9_4_clk =
     1'b1 ? clk : 1'd0;
    assign left_9_4_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? left_9_3_out : 32'd0;
    assign left_9_4_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign left_9_5_clk =
     1'b1 ? clk : 1'd0;
    assign left_9_5_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? left_9_4_out : 32'd0;
    assign left_9_5_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign left_9_6_clk =
     1'b1 ? clk : 1'd0;
    assign left_9_6_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? left_9_5_out : 32'd0;
    assign left_9_6_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign left_9_7_clk =
     1'b1 ? clk : 1'd0;
    assign left_9_7_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? left_9_6_out : 32'd0;
    assign left_9_7_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign left_9_8_clk =
     1'b1 ? clk : 1'd0;
    assign left_9_8_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? left_9_7_out : 32'd0;
    assign left_9_8_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign left_9_9_clk =
     1'b1 ? clk : 1'd0;
    assign left_9_9_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? left_9_8_out : 32'd0;
    assign left_9_9_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign pe_0_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_0_go =
     fsm2_out < 3'd5 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd5 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go ? 1'd1 : 1'd0;
    assign pe_0_0_left =
     fsm2_out < 3'd5 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd5 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go ? left_0_0_out : 32'd0;
    assign pe_0_0_top =
     fsm2_out < 3'd5 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd5 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go ? top_0_0_out : 32'd0;
    assign pe_0_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_1_go =
     fsm4_out < 3'd5 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? 1'd1 : 1'd0;
    assign pe_0_1_left =
     fsm4_out < 3'd5 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? left_0_1_out : 32'd0;
    assign pe_0_1_top =
     fsm4_out < 3'd5 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? top_0_1_out : 32'd0;
    assign pe_0_10_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_10_go =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? 1'd1 : 1'd0;
    assign pe_0_10_left =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? left_0_10_out : 32'd0;
    assign pe_0_10_top =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? top_0_10_out : 32'd0;
    assign pe_0_11_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_11_go =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 1'd1 : 1'd0;
    assign pe_0_11_left =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? left_0_11_out : 32'd0;
    assign pe_0_11_top =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? top_0_11_out : 32'd0;
    assign pe_0_12_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_12_go =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 1'd1 : 1'd0;
    assign pe_0_12_left =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? left_0_12_out : 32'd0;
    assign pe_0_12_top =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? top_0_12_out : 32'd0;
    assign pe_0_13_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_13_go =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 1'd1 : 1'd0;
    assign pe_0_13_left =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? left_0_13_out : 32'd0;
    assign pe_0_13_top =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? top_0_13_out : 32'd0;
    assign pe_0_14_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_14_go =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign pe_0_14_left =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? left_0_14_out : 32'd0;
    assign pe_0_14_top =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? top_0_14_out : 32'd0;
    assign pe_0_15_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_15_go =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 1'd1 : 1'd0;
    assign pe_0_15_left =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? left_0_15_out : 32'd0;
    assign pe_0_15_top =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? top_0_15_out : 32'd0;
    assign pe_0_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_2_go =
     fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? 1'd1 : 1'd0;
    assign pe_0_2_left =
     fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? left_0_2_out : 32'd0;
    assign pe_0_2_top =
     fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? top_0_2_out : 32'd0;
    assign pe_0_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_3_go =
     fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? 1'd1 : 1'd0;
    assign pe_0_3_left =
     fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? left_0_3_out : 32'd0;
    assign pe_0_3_top =
     fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? top_0_3_out : 32'd0;
    assign pe_0_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_4_go =
     fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? 1'd1 : 1'd0;
    assign pe_0_4_left =
     fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? left_0_4_out : 32'd0;
    assign pe_0_4_top =
     fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? top_0_4_out : 32'd0;
    assign pe_0_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_5_go =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? 1'd1 : 1'd0;
    assign pe_0_5_left =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? left_0_5_out : 32'd0;
    assign pe_0_5_top =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? top_0_5_out : 32'd0;
    assign pe_0_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_6_go =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? 1'd1 : 1'd0;
    assign pe_0_6_left =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? left_0_6_out : 32'd0;
    assign pe_0_6_top =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? top_0_6_out : 32'd0;
    assign pe_0_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_7_go =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? 1'd1 : 1'd0;
    assign pe_0_7_left =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? left_0_7_out : 32'd0;
    assign pe_0_7_top =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? top_0_7_out : 32'd0;
    assign pe_0_8_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_8_go =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? 1'd1 : 1'd0;
    assign pe_0_8_left =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? left_0_8_out : 32'd0;
    assign pe_0_8_top =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? top_0_8_out : 32'd0;
    assign pe_0_9_clk =
     1'b1 ? clk : 1'd0;
    assign pe_0_9_go =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? 1'd1 : 1'd0;
    assign pe_0_9_left =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? left_0_9_out : 32'd0;
    assign pe_0_9_top =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? top_0_9_out : 32'd0;
    assign pe_10_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_10_0_go =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? 1'd1 : 1'd0;
    assign pe_10_0_left =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? left_10_0_out : 32'd0;
    assign pe_10_0_top =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? top_10_0_out : 32'd0;
    assign pe_10_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_10_1_go =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 1'd1 : 1'd0;
    assign pe_10_1_left =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? left_10_1_out : 32'd0;
    assign pe_10_1_top =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? top_10_1_out : 32'd0;
    assign pe_10_10_clk =
     1'b1 ? clk : 1'd0;
    assign pe_10_10_go =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? 1'd1 : 1'd0;
    assign pe_10_10_left =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? left_10_10_out : 32'd0;
    assign pe_10_10_top =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? top_10_10_out : 32'd0;
    assign pe_10_11_clk =
     1'b1 ? clk : 1'd0;
    assign pe_10_11_go =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? 1'd1 : 1'd0;
    assign pe_10_11_left =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? left_10_11_out : 32'd0;
    assign pe_10_11_top =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? top_10_11_out : 32'd0;
    assign pe_10_12_clk =
     1'b1 ? clk : 1'd0;
    assign pe_10_12_go =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? 1'd1 : 1'd0;
    assign pe_10_12_left =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? left_10_12_out : 32'd0;
    assign pe_10_12_top =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? top_10_12_out : 32'd0;
    assign pe_10_13_clk =
     1'b1 ? clk : 1'd0;
    assign pe_10_13_go =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? 1'd1 : 1'd0;
    assign pe_10_13_left =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? left_10_13_out : 32'd0;
    assign pe_10_13_top =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? top_10_13_out : 32'd0;
    assign pe_10_14_clk =
     1'b1 ? clk : 1'd0;
    assign pe_10_14_go =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? 1'd1 : 1'd0;
    assign pe_10_14_left =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? left_10_14_out : 32'd0;
    assign pe_10_14_top =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? top_10_14_out : 32'd0;
    assign pe_10_15_clk =
     1'b1 ? clk : 1'd0;
    assign pe_10_15_go =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? 1'd1 : 1'd0;
    assign pe_10_15_left =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? left_10_15_out : 32'd0;
    assign pe_10_15_top =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? top_10_15_out : 32'd0;
    assign pe_10_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_10_2_go =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 1'd1 : 1'd0;
    assign pe_10_2_left =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? left_10_2_out : 32'd0;
    assign pe_10_2_top =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? top_10_2_out : 32'd0;
    assign pe_10_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_10_3_go =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 1'd1 : 1'd0;
    assign pe_10_3_left =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? left_10_3_out : 32'd0;
    assign pe_10_3_top =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? top_10_3_out : 32'd0;
    assign pe_10_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_10_4_go =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign pe_10_4_left =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? left_10_4_out : 32'd0;
    assign pe_10_4_top =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? top_10_4_out : 32'd0;
    assign pe_10_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_10_5_go =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 1'd1 : 1'd0;
    assign pe_10_5_left =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? left_10_5_out : 32'd0;
    assign pe_10_5_top =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? top_10_5_out : 32'd0;
    assign pe_10_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_10_6_go =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? 1'd1 : 1'd0;
    assign pe_10_6_left =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? left_10_6_out : 32'd0;
    assign pe_10_6_top =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? top_10_6_out : 32'd0;
    assign pe_10_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_10_7_go =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? 1'd1 : 1'd0;
    assign pe_10_7_left =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? left_10_7_out : 32'd0;
    assign pe_10_7_top =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? top_10_7_out : 32'd0;
    assign pe_10_8_clk =
     1'b1 ? clk : 1'd0;
    assign pe_10_8_go =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? 1'd1 : 1'd0;
    assign pe_10_8_left =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? left_10_8_out : 32'd0;
    assign pe_10_8_top =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? top_10_8_out : 32'd0;
    assign pe_10_9_clk =
     1'b1 ? clk : 1'd0;
    assign pe_10_9_go =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? 1'd1 : 1'd0;
    assign pe_10_9_left =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? left_10_9_out : 32'd0;
    assign pe_10_9_top =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? top_10_9_out : 32'd0;
    assign pe_11_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_11_0_go =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 1'd1 : 1'd0;
    assign pe_11_0_left =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? left_11_0_out : 32'd0;
    assign pe_11_0_top =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? top_11_0_out : 32'd0;
    assign pe_11_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_11_1_go =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 1'd1 : 1'd0;
    assign pe_11_1_left =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? left_11_1_out : 32'd0;
    assign pe_11_1_top =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? top_11_1_out : 32'd0;
    assign pe_11_10_clk =
     1'b1 ? clk : 1'd0;
    assign pe_11_10_go =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? 1'd1 : 1'd0;
    assign pe_11_10_left =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? left_11_10_out : 32'd0;
    assign pe_11_10_top =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? top_11_10_out : 32'd0;
    assign pe_11_11_clk =
     1'b1 ? clk : 1'd0;
    assign pe_11_11_go =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? 1'd1 : 1'd0;
    assign pe_11_11_left =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? left_11_11_out : 32'd0;
    assign pe_11_11_top =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? top_11_11_out : 32'd0;
    assign pe_11_12_clk =
     1'b1 ? clk : 1'd0;
    assign pe_11_12_go =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? 1'd1 : 1'd0;
    assign pe_11_12_left =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? left_11_12_out : 32'd0;
    assign pe_11_12_top =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? top_11_12_out : 32'd0;
    assign pe_11_13_clk =
     1'b1 ? clk : 1'd0;
    assign pe_11_13_go =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? 1'd1 : 1'd0;
    assign pe_11_13_left =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? left_11_13_out : 32'd0;
    assign pe_11_13_top =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? top_11_13_out : 32'd0;
    assign pe_11_14_clk =
     1'b1 ? clk : 1'd0;
    assign pe_11_14_go =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? 1'd1 : 1'd0;
    assign pe_11_14_left =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? left_11_14_out : 32'd0;
    assign pe_11_14_top =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? top_11_14_out : 32'd0;
    assign pe_11_15_clk =
     1'b1 ? clk : 1'd0;
    assign pe_11_15_go =
     fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? 1'd1 : 1'd0;
    assign pe_11_15_left =
     fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? left_11_15_out : 32'd0;
    assign pe_11_15_top =
     fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? top_11_15_out : 32'd0;
    assign pe_11_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_11_2_go =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 1'd1 : 1'd0;
    assign pe_11_2_left =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? left_11_2_out : 32'd0;
    assign pe_11_2_top =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? top_11_2_out : 32'd0;
    assign pe_11_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_11_3_go =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign pe_11_3_left =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? left_11_3_out : 32'd0;
    assign pe_11_3_top =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? top_11_3_out : 32'd0;
    assign pe_11_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_11_4_go =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 1'd1 : 1'd0;
    assign pe_11_4_left =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? left_11_4_out : 32'd0;
    assign pe_11_4_top =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? top_11_4_out : 32'd0;
    assign pe_11_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_11_5_go =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? 1'd1 : 1'd0;
    assign pe_11_5_left =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? left_11_5_out : 32'd0;
    assign pe_11_5_top =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? top_11_5_out : 32'd0;
    assign pe_11_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_11_6_go =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? 1'd1 : 1'd0;
    assign pe_11_6_left =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? left_11_6_out : 32'd0;
    assign pe_11_6_top =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? top_11_6_out : 32'd0;
    assign pe_11_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_11_7_go =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? 1'd1 : 1'd0;
    assign pe_11_7_left =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? left_11_7_out : 32'd0;
    assign pe_11_7_top =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? top_11_7_out : 32'd0;
    assign pe_11_8_clk =
     1'b1 ? clk : 1'd0;
    assign pe_11_8_go =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? 1'd1 : 1'd0;
    assign pe_11_8_left =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? left_11_8_out : 32'd0;
    assign pe_11_8_top =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? top_11_8_out : 32'd0;
    assign pe_11_9_clk =
     1'b1 ? clk : 1'd0;
    assign pe_11_9_go =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? 1'd1 : 1'd0;
    assign pe_11_9_left =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? left_11_9_out : 32'd0;
    assign pe_11_9_top =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? top_11_9_out : 32'd0;
    assign pe_12_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_12_0_go =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 1'd1 : 1'd0;
    assign pe_12_0_left =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? left_12_0_out : 32'd0;
    assign pe_12_0_top =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? top_12_0_out : 32'd0;
    assign pe_12_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_12_1_go =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 1'd1 : 1'd0;
    assign pe_12_1_left =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? left_12_1_out : 32'd0;
    assign pe_12_1_top =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? top_12_1_out : 32'd0;
    assign pe_12_10_clk =
     1'b1 ? clk : 1'd0;
    assign pe_12_10_go =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? 1'd1 : 1'd0;
    assign pe_12_10_left =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? left_12_10_out : 32'd0;
    assign pe_12_10_top =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? top_12_10_out : 32'd0;
    assign pe_12_11_clk =
     1'b1 ? clk : 1'd0;
    assign pe_12_11_go =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? 1'd1 : 1'd0;
    assign pe_12_11_left =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? left_12_11_out : 32'd0;
    assign pe_12_11_top =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? top_12_11_out : 32'd0;
    assign pe_12_12_clk =
     1'b1 ? clk : 1'd0;
    assign pe_12_12_go =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? 1'd1 : 1'd0;
    assign pe_12_12_left =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? left_12_12_out : 32'd0;
    assign pe_12_12_top =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? top_12_12_out : 32'd0;
    assign pe_12_13_clk =
     1'b1 ? clk : 1'd0;
    assign pe_12_13_go =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? 1'd1 : 1'd0;
    assign pe_12_13_left =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? left_12_13_out : 32'd0;
    assign pe_12_13_top =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? top_12_13_out : 32'd0;
    assign pe_12_14_clk =
     1'b1 ? clk : 1'd0;
    assign pe_12_14_go =
     fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? 1'd1 : 1'd0;
    assign pe_12_14_left =
     fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? left_12_14_out : 32'd0;
    assign pe_12_14_top =
     fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? top_12_14_out : 32'd0;
    assign pe_12_15_clk =
     1'b1 ? clk : 1'd0;
    assign pe_12_15_go =
     fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go ? 1'd1 : 1'd0;
    assign pe_12_15_left =
     fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go ? left_12_15_out : 32'd0;
    assign pe_12_15_top =
     fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go ? top_12_15_out : 32'd0;
    assign pe_12_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_12_2_go =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign pe_12_2_left =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? left_12_2_out : 32'd0;
    assign pe_12_2_top =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? top_12_2_out : 32'd0;
    assign pe_12_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_12_3_go =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 1'd1 : 1'd0;
    assign pe_12_3_left =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? left_12_3_out : 32'd0;
    assign pe_12_3_top =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? top_12_3_out : 32'd0;
    assign pe_12_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_12_4_go =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? 1'd1 : 1'd0;
    assign pe_12_4_left =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? left_12_4_out : 32'd0;
    assign pe_12_4_top =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? top_12_4_out : 32'd0;
    assign pe_12_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_12_5_go =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? 1'd1 : 1'd0;
    assign pe_12_5_left =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? left_12_5_out : 32'd0;
    assign pe_12_5_top =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? top_12_5_out : 32'd0;
    assign pe_12_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_12_6_go =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? 1'd1 : 1'd0;
    assign pe_12_6_left =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? left_12_6_out : 32'd0;
    assign pe_12_6_top =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? top_12_6_out : 32'd0;
    assign pe_12_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_12_7_go =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? 1'd1 : 1'd0;
    assign pe_12_7_left =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? left_12_7_out : 32'd0;
    assign pe_12_7_top =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? top_12_7_out : 32'd0;
    assign pe_12_8_clk =
     1'b1 ? clk : 1'd0;
    assign pe_12_8_go =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? 1'd1 : 1'd0;
    assign pe_12_8_left =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? left_12_8_out : 32'd0;
    assign pe_12_8_top =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? top_12_8_out : 32'd0;
    assign pe_12_9_clk =
     1'b1 ? clk : 1'd0;
    assign pe_12_9_go =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? 1'd1 : 1'd0;
    assign pe_12_9_left =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? left_12_9_out : 32'd0;
    assign pe_12_9_top =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? top_12_9_out : 32'd0;
    assign pe_13_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_13_0_go =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 1'd1 : 1'd0;
    assign pe_13_0_left =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? left_13_0_out : 32'd0;
    assign pe_13_0_top =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? top_13_0_out : 32'd0;
    assign pe_13_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_13_1_go =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign pe_13_1_left =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? left_13_1_out : 32'd0;
    assign pe_13_1_top =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? top_13_1_out : 32'd0;
    assign pe_13_10_clk =
     1'b1 ? clk : 1'd0;
    assign pe_13_10_go =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? 1'd1 : 1'd0;
    assign pe_13_10_left =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? left_13_10_out : 32'd0;
    assign pe_13_10_top =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? top_13_10_out : 32'd0;
    assign pe_13_11_clk =
     1'b1 ? clk : 1'd0;
    assign pe_13_11_go =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? 1'd1 : 1'd0;
    assign pe_13_11_left =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? left_13_11_out : 32'd0;
    assign pe_13_11_top =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? top_13_11_out : 32'd0;
    assign pe_13_12_clk =
     1'b1 ? clk : 1'd0;
    assign pe_13_12_go =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? 1'd1 : 1'd0;
    assign pe_13_12_left =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? left_13_12_out : 32'd0;
    assign pe_13_12_top =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? top_13_12_out : 32'd0;
    assign pe_13_13_clk =
     1'b1 ? clk : 1'd0;
    assign pe_13_13_go =
     fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? 1'd1 : 1'd0;
    assign pe_13_13_left =
     fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? left_13_13_out : 32'd0;
    assign pe_13_13_top =
     fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? top_13_13_out : 32'd0;
    assign pe_13_14_clk =
     1'b1 ? clk : 1'd0;
    assign pe_13_14_go =
     fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go ? 1'd1 : 1'd0;
    assign pe_13_14_left =
     fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go ? left_13_14_out : 32'd0;
    assign pe_13_14_top =
     fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go ? top_13_14_out : 32'd0;
    assign pe_13_15_clk =
     1'b1 ? clk : 1'd0;
    assign pe_13_15_go =
     fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go ? 1'd1 : 1'd0;
    assign pe_13_15_left =
     fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go ? left_13_15_out : 32'd0;
    assign pe_13_15_top =
     fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go ? top_13_15_out : 32'd0;
    assign pe_13_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_13_2_go =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 1'd1 : 1'd0;
    assign pe_13_2_left =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? left_13_2_out : 32'd0;
    assign pe_13_2_top =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? top_13_2_out : 32'd0;
    assign pe_13_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_13_3_go =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? 1'd1 : 1'd0;
    assign pe_13_3_left =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? left_13_3_out : 32'd0;
    assign pe_13_3_top =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? top_13_3_out : 32'd0;
    assign pe_13_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_13_4_go =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? 1'd1 : 1'd0;
    assign pe_13_4_left =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? left_13_4_out : 32'd0;
    assign pe_13_4_top =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? top_13_4_out : 32'd0;
    assign pe_13_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_13_5_go =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? 1'd1 : 1'd0;
    assign pe_13_5_left =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? left_13_5_out : 32'd0;
    assign pe_13_5_top =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? top_13_5_out : 32'd0;
    assign pe_13_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_13_6_go =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? 1'd1 : 1'd0;
    assign pe_13_6_left =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? left_13_6_out : 32'd0;
    assign pe_13_6_top =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? top_13_6_out : 32'd0;
    assign pe_13_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_13_7_go =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? 1'd1 : 1'd0;
    assign pe_13_7_left =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? left_13_7_out : 32'd0;
    assign pe_13_7_top =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? top_13_7_out : 32'd0;
    assign pe_13_8_clk =
     1'b1 ? clk : 1'd0;
    assign pe_13_8_go =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? 1'd1 : 1'd0;
    assign pe_13_8_left =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? left_13_8_out : 32'd0;
    assign pe_13_8_top =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? top_13_8_out : 32'd0;
    assign pe_13_9_clk =
     1'b1 ? clk : 1'd0;
    assign pe_13_9_go =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? 1'd1 : 1'd0;
    assign pe_13_9_left =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? left_13_9_out : 32'd0;
    assign pe_13_9_top =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? top_13_9_out : 32'd0;
    assign pe_14_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_14_0_go =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign pe_14_0_left =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? left_14_0_out : 32'd0;
    assign pe_14_0_top =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? top_14_0_out : 32'd0;
    assign pe_14_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_14_1_go =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 1'd1 : 1'd0;
    assign pe_14_1_left =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? left_14_1_out : 32'd0;
    assign pe_14_1_top =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? top_14_1_out : 32'd0;
    assign pe_14_10_clk =
     1'b1 ? clk : 1'd0;
    assign pe_14_10_go =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? 1'd1 : 1'd0;
    assign pe_14_10_left =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? left_14_10_out : 32'd0;
    assign pe_14_10_top =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? top_14_10_out : 32'd0;
    assign pe_14_11_clk =
     1'b1 ? clk : 1'd0;
    assign pe_14_11_go =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? 1'd1 : 1'd0;
    assign pe_14_11_left =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? left_14_11_out : 32'd0;
    assign pe_14_11_top =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? top_14_11_out : 32'd0;
    assign pe_14_12_clk =
     1'b1 ? clk : 1'd0;
    assign pe_14_12_go =
     fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? 1'd1 : 1'd0;
    assign pe_14_12_left =
     fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? left_14_12_out : 32'd0;
    assign pe_14_12_top =
     fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? top_14_12_out : 32'd0;
    assign pe_14_13_clk =
     1'b1 ? clk : 1'd0;
    assign pe_14_13_go =
     fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go ? 1'd1 : 1'd0;
    assign pe_14_13_left =
     fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go ? left_14_13_out : 32'd0;
    assign pe_14_13_top =
     fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go ? top_14_13_out : 32'd0;
    assign pe_14_14_clk =
     1'b1 ? clk : 1'd0;
    assign pe_14_14_go =
     fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go ? 1'd1 : 1'd0;
    assign pe_14_14_left =
     fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go ? left_14_14_out : 32'd0;
    assign pe_14_14_top =
     fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go ? top_14_14_out : 32'd0;
    assign pe_14_15_clk =
     1'b1 ? clk : 1'd0;
    assign pe_14_15_go =
     fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go | fsm90_out < 3'd5 & fsm92_out >= 10'd267 & fsm92_out < 10'd272 & go ? 1'd1 : 1'd0;
    assign pe_14_15_left =
     fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go | fsm90_out < 3'd5 & fsm92_out >= 10'd267 & fsm92_out < 10'd272 & go ? left_14_15_out : 32'd0;
    assign pe_14_15_top =
     fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go | fsm90_out < 3'd5 & fsm92_out >= 10'd267 & fsm92_out < 10'd272 & go ? top_14_15_out : 32'd0;
    assign pe_14_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_14_2_go =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? 1'd1 : 1'd0;
    assign pe_14_2_left =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? left_14_2_out : 32'd0;
    assign pe_14_2_top =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? top_14_2_out : 32'd0;
    assign pe_14_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_14_3_go =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? 1'd1 : 1'd0;
    assign pe_14_3_left =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? left_14_3_out : 32'd0;
    assign pe_14_3_top =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? top_14_3_out : 32'd0;
    assign pe_14_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_14_4_go =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? 1'd1 : 1'd0;
    assign pe_14_4_left =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? left_14_4_out : 32'd0;
    assign pe_14_4_top =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? top_14_4_out : 32'd0;
    assign pe_14_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_14_5_go =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? 1'd1 : 1'd0;
    assign pe_14_5_left =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? left_14_5_out : 32'd0;
    assign pe_14_5_top =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? top_14_5_out : 32'd0;
    assign pe_14_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_14_6_go =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? 1'd1 : 1'd0;
    assign pe_14_6_left =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? left_14_6_out : 32'd0;
    assign pe_14_6_top =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? top_14_6_out : 32'd0;
    assign pe_14_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_14_7_go =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? 1'd1 : 1'd0;
    assign pe_14_7_left =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? left_14_7_out : 32'd0;
    assign pe_14_7_top =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? top_14_7_out : 32'd0;
    assign pe_14_8_clk =
     1'b1 ? clk : 1'd0;
    assign pe_14_8_go =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? 1'd1 : 1'd0;
    assign pe_14_8_left =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? left_14_8_out : 32'd0;
    assign pe_14_8_top =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? top_14_8_out : 32'd0;
    assign pe_14_9_clk =
     1'b1 ? clk : 1'd0;
    assign pe_14_9_go =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? 1'd1 : 1'd0;
    assign pe_14_9_left =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? left_14_9_out : 32'd0;
    assign pe_14_9_top =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? top_14_9_out : 32'd0;
    assign pe_15_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_15_0_go =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 1'd1 : 1'd0;
    assign pe_15_0_left =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? left_15_0_out : 32'd0;
    assign pe_15_0_top =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? top_15_0_out : 32'd0;
    assign pe_15_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_15_1_go =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? 1'd1 : 1'd0;
    assign pe_15_1_left =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? left_15_1_out : 32'd0;
    assign pe_15_1_top =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? top_15_1_out : 32'd0;
    assign pe_15_10_clk =
     1'b1 ? clk : 1'd0;
    assign pe_15_10_go =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? 1'd1 : 1'd0;
    assign pe_15_10_left =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? left_15_10_out : 32'd0;
    assign pe_15_10_top =
     fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go ? top_15_10_out : 32'd0;
    assign pe_15_11_clk =
     1'b1 ? clk : 1'd0;
    assign pe_15_11_go =
     fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? 1'd1 : 1'd0;
    assign pe_15_11_left =
     fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? left_15_11_out : 32'd0;
    assign pe_15_11_top =
     fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go ? top_15_11_out : 32'd0;
    assign pe_15_12_clk =
     1'b1 ? clk : 1'd0;
    assign pe_15_12_go =
     fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go ? 1'd1 : 1'd0;
    assign pe_15_12_left =
     fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go ? left_15_12_out : 32'd0;
    assign pe_15_12_top =
     fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go ? top_15_12_out : 32'd0;
    assign pe_15_13_clk =
     1'b1 ? clk : 1'd0;
    assign pe_15_13_go =
     fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go ? 1'd1 : 1'd0;
    assign pe_15_13_left =
     fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go ? left_15_13_out : 32'd0;
    assign pe_15_13_top =
     fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go ? top_15_13_out : 32'd0;
    assign pe_15_14_clk =
     1'b1 ? clk : 1'd0;
    assign pe_15_14_go =
     fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go | fsm90_out < 3'd5 & fsm92_out >= 10'd267 & fsm92_out < 10'd272 & go ? 1'd1 : 1'd0;
    assign pe_15_14_left =
     fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go | fsm90_out < 3'd5 & fsm92_out >= 10'd267 & fsm92_out < 10'd272 & go ? left_15_14_out : 32'd0;
    assign pe_15_14_top =
     fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go | fsm90_out < 3'd5 & fsm92_out >= 10'd267 & fsm92_out < 10'd272 & go ? top_15_14_out : 32'd0;
    assign pe_15_15_clk =
     1'b1 ? clk : 1'd0;
    assign pe_15_15_go =
     fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go | fsm90_out < 3'd5 & fsm92_out >= 10'd267 & fsm92_out < 10'd272 & go | fsm92_out >= 10'd273 & fsm92_out < 10'd278 & go ? 1'd1 : 1'd0;
    assign pe_15_15_left =
     fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go | fsm90_out < 3'd5 & fsm92_out >= 10'd267 & fsm92_out < 10'd272 & go | fsm92_out >= 10'd273 & fsm92_out < 10'd278 & go ? left_15_15_out : 32'd0;
    assign pe_15_15_top =
     fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go | fsm82_out < 3'd5 & fsm92_out >= 10'd243 & fsm92_out < 10'd248 & go | fsm84_out < 3'd5 & fsm92_out >= 10'd249 & fsm92_out < 10'd254 & go | fsm86_out < 3'd5 & fsm92_out >= 10'd255 & fsm92_out < 10'd260 & go | fsm88_out < 3'd5 & fsm92_out >= 10'd261 & fsm92_out < 10'd266 & go | fsm90_out < 3'd5 & fsm92_out >= 10'd267 & fsm92_out < 10'd272 & go | fsm92_out >= 10'd273 & fsm92_out < 10'd278 & go ? top_15_15_out : 32'd0;
    assign pe_15_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_15_2_go =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? 1'd1 : 1'd0;
    assign pe_15_2_left =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? left_15_2_out : 32'd0;
    assign pe_15_2_top =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? top_15_2_out : 32'd0;
    assign pe_15_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_15_3_go =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? 1'd1 : 1'd0;
    assign pe_15_3_left =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? left_15_3_out : 32'd0;
    assign pe_15_3_top =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? top_15_3_out : 32'd0;
    assign pe_15_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_15_4_go =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? 1'd1 : 1'd0;
    assign pe_15_4_left =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? left_15_4_out : 32'd0;
    assign pe_15_4_top =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? top_15_4_out : 32'd0;
    assign pe_15_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_15_5_go =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? 1'd1 : 1'd0;
    assign pe_15_5_left =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? left_15_5_out : 32'd0;
    assign pe_15_5_top =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? top_15_5_out : 32'd0;
    assign pe_15_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_15_6_go =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? 1'd1 : 1'd0;
    assign pe_15_6_left =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? left_15_6_out : 32'd0;
    assign pe_15_6_top =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? top_15_6_out : 32'd0;
    assign pe_15_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_15_7_go =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? 1'd1 : 1'd0;
    assign pe_15_7_left =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? left_15_7_out : 32'd0;
    assign pe_15_7_top =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? top_15_7_out : 32'd0;
    assign pe_15_8_clk =
     1'b1 ? clk : 1'd0;
    assign pe_15_8_go =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? 1'd1 : 1'd0;
    assign pe_15_8_left =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? left_15_8_out : 32'd0;
    assign pe_15_8_top =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? top_15_8_out : 32'd0;
    assign pe_15_9_clk =
     1'b1 ? clk : 1'd0;
    assign pe_15_9_go =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? 1'd1 : 1'd0;
    assign pe_15_9_left =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? left_15_9_out : 32'd0;
    assign pe_15_9_top =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? top_15_9_out : 32'd0;
    assign pe_1_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_0_go =
     fsm4_out < 3'd5 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? 1'd1 : 1'd0;
    assign pe_1_0_left =
     fsm4_out < 3'd5 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? left_1_0_out : 32'd0;
    assign pe_1_0_top =
     fsm4_out < 3'd5 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? top_1_0_out : 32'd0;
    assign pe_1_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_1_go =
     fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? 1'd1 : 1'd0;
    assign pe_1_1_left =
     fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? left_1_1_out : 32'd0;
    assign pe_1_1_top =
     fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? top_1_1_out : 32'd0;
    assign pe_1_10_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_10_go =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 1'd1 : 1'd0;
    assign pe_1_10_left =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? left_1_10_out : 32'd0;
    assign pe_1_10_top =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? top_1_10_out : 32'd0;
    assign pe_1_11_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_11_go =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 1'd1 : 1'd0;
    assign pe_1_11_left =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? left_1_11_out : 32'd0;
    assign pe_1_11_top =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? top_1_11_out : 32'd0;
    assign pe_1_12_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_12_go =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 1'd1 : 1'd0;
    assign pe_1_12_left =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? left_1_12_out : 32'd0;
    assign pe_1_12_top =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? top_1_12_out : 32'd0;
    assign pe_1_13_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_13_go =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign pe_1_13_left =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? left_1_13_out : 32'd0;
    assign pe_1_13_top =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? top_1_13_out : 32'd0;
    assign pe_1_14_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_14_go =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 1'd1 : 1'd0;
    assign pe_1_14_left =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? left_1_14_out : 32'd0;
    assign pe_1_14_top =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? top_1_14_out : 32'd0;
    assign pe_1_15_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_15_go =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? 1'd1 : 1'd0;
    assign pe_1_15_left =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? left_1_15_out : 32'd0;
    assign pe_1_15_top =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? top_1_15_out : 32'd0;
    assign pe_1_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_2_go =
     fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? 1'd1 : 1'd0;
    assign pe_1_2_left =
     fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? left_1_2_out : 32'd0;
    assign pe_1_2_top =
     fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? top_1_2_out : 32'd0;
    assign pe_1_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_3_go =
     fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? 1'd1 : 1'd0;
    assign pe_1_3_left =
     fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? left_1_3_out : 32'd0;
    assign pe_1_3_top =
     fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? top_1_3_out : 32'd0;
    assign pe_1_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_4_go =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? 1'd1 : 1'd0;
    assign pe_1_4_left =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? left_1_4_out : 32'd0;
    assign pe_1_4_top =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? top_1_4_out : 32'd0;
    assign pe_1_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_5_go =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? 1'd1 : 1'd0;
    assign pe_1_5_left =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? left_1_5_out : 32'd0;
    assign pe_1_5_top =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? top_1_5_out : 32'd0;
    assign pe_1_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_6_go =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? 1'd1 : 1'd0;
    assign pe_1_6_left =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? left_1_6_out : 32'd0;
    assign pe_1_6_top =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? top_1_6_out : 32'd0;
    assign pe_1_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_7_go =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? 1'd1 : 1'd0;
    assign pe_1_7_left =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? left_1_7_out : 32'd0;
    assign pe_1_7_top =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? top_1_7_out : 32'd0;
    assign pe_1_8_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_8_go =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? 1'd1 : 1'd0;
    assign pe_1_8_left =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? left_1_8_out : 32'd0;
    assign pe_1_8_top =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? top_1_8_out : 32'd0;
    assign pe_1_9_clk =
     1'b1 ? clk : 1'd0;
    assign pe_1_9_go =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? 1'd1 : 1'd0;
    assign pe_1_9_left =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? left_1_9_out : 32'd0;
    assign pe_1_9_top =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? top_1_9_out : 32'd0;
    assign pe_2_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_0_go =
     fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? 1'd1 : 1'd0;
    assign pe_2_0_left =
     fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? left_2_0_out : 32'd0;
    assign pe_2_0_top =
     fsm6_out < 3'd5 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? top_2_0_out : 32'd0;
    assign pe_2_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_1_go =
     fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? 1'd1 : 1'd0;
    assign pe_2_1_left =
     fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? left_2_1_out : 32'd0;
    assign pe_2_1_top =
     fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? top_2_1_out : 32'd0;
    assign pe_2_10_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_10_go =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 1'd1 : 1'd0;
    assign pe_2_10_left =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? left_2_10_out : 32'd0;
    assign pe_2_10_top =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? top_2_10_out : 32'd0;
    assign pe_2_11_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_11_go =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 1'd1 : 1'd0;
    assign pe_2_11_left =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? left_2_11_out : 32'd0;
    assign pe_2_11_top =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? top_2_11_out : 32'd0;
    assign pe_2_12_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_12_go =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign pe_2_12_left =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? left_2_12_out : 32'd0;
    assign pe_2_12_top =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? top_2_12_out : 32'd0;
    assign pe_2_13_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_13_go =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 1'd1 : 1'd0;
    assign pe_2_13_left =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? left_2_13_out : 32'd0;
    assign pe_2_13_top =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? top_2_13_out : 32'd0;
    assign pe_2_14_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_14_go =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? 1'd1 : 1'd0;
    assign pe_2_14_left =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? left_2_14_out : 32'd0;
    assign pe_2_14_top =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? top_2_14_out : 32'd0;
    assign pe_2_15_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_15_go =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? 1'd1 : 1'd0;
    assign pe_2_15_left =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? left_2_15_out : 32'd0;
    assign pe_2_15_top =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? top_2_15_out : 32'd0;
    assign pe_2_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_2_go =
     fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? 1'd1 : 1'd0;
    assign pe_2_2_left =
     fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? left_2_2_out : 32'd0;
    assign pe_2_2_top =
     fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? top_2_2_out : 32'd0;
    assign pe_2_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_3_go =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? 1'd1 : 1'd0;
    assign pe_2_3_left =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? left_2_3_out : 32'd0;
    assign pe_2_3_top =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? top_2_3_out : 32'd0;
    assign pe_2_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_4_go =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? 1'd1 : 1'd0;
    assign pe_2_4_left =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? left_2_4_out : 32'd0;
    assign pe_2_4_top =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? top_2_4_out : 32'd0;
    assign pe_2_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_5_go =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? 1'd1 : 1'd0;
    assign pe_2_5_left =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? left_2_5_out : 32'd0;
    assign pe_2_5_top =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? top_2_5_out : 32'd0;
    assign pe_2_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_6_go =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? 1'd1 : 1'd0;
    assign pe_2_6_left =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? left_2_6_out : 32'd0;
    assign pe_2_6_top =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? top_2_6_out : 32'd0;
    assign pe_2_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_7_go =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? 1'd1 : 1'd0;
    assign pe_2_7_left =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? left_2_7_out : 32'd0;
    assign pe_2_7_top =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? top_2_7_out : 32'd0;
    assign pe_2_8_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_8_go =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? 1'd1 : 1'd0;
    assign pe_2_8_left =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? left_2_8_out : 32'd0;
    assign pe_2_8_top =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? top_2_8_out : 32'd0;
    assign pe_2_9_clk =
     1'b1 ? clk : 1'd0;
    assign pe_2_9_go =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 1'd1 : 1'd0;
    assign pe_2_9_left =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? left_2_9_out : 32'd0;
    assign pe_2_9_top =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? top_2_9_out : 32'd0;
    assign pe_3_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_0_go =
     fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? 1'd1 : 1'd0;
    assign pe_3_0_left =
     fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? left_3_0_out : 32'd0;
    assign pe_3_0_top =
     fsm8_out < 3'd5 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? top_3_0_out : 32'd0;
    assign pe_3_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_1_go =
     fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? 1'd1 : 1'd0;
    assign pe_3_1_left =
     fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? left_3_1_out : 32'd0;
    assign pe_3_1_top =
     fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? top_3_1_out : 32'd0;
    assign pe_3_10_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_10_go =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 1'd1 : 1'd0;
    assign pe_3_10_left =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? left_3_10_out : 32'd0;
    assign pe_3_10_top =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? top_3_10_out : 32'd0;
    assign pe_3_11_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_11_go =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign pe_3_11_left =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? left_3_11_out : 32'd0;
    assign pe_3_11_top =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? top_3_11_out : 32'd0;
    assign pe_3_12_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_12_go =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 1'd1 : 1'd0;
    assign pe_3_12_left =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? left_3_12_out : 32'd0;
    assign pe_3_12_top =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? top_3_12_out : 32'd0;
    assign pe_3_13_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_13_go =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? 1'd1 : 1'd0;
    assign pe_3_13_left =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? left_3_13_out : 32'd0;
    assign pe_3_13_top =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? top_3_13_out : 32'd0;
    assign pe_3_14_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_14_go =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? 1'd1 : 1'd0;
    assign pe_3_14_left =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? left_3_14_out : 32'd0;
    assign pe_3_14_top =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? top_3_14_out : 32'd0;
    assign pe_3_15_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_15_go =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? 1'd1 : 1'd0;
    assign pe_3_15_left =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? left_3_15_out : 32'd0;
    assign pe_3_15_top =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? top_3_15_out : 32'd0;
    assign pe_3_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_2_go =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? 1'd1 : 1'd0;
    assign pe_3_2_left =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? left_3_2_out : 32'd0;
    assign pe_3_2_top =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? top_3_2_out : 32'd0;
    assign pe_3_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_3_go =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? 1'd1 : 1'd0;
    assign pe_3_3_left =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? left_3_3_out : 32'd0;
    assign pe_3_3_top =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? top_3_3_out : 32'd0;
    assign pe_3_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_4_go =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? 1'd1 : 1'd0;
    assign pe_3_4_left =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? left_3_4_out : 32'd0;
    assign pe_3_4_top =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? top_3_4_out : 32'd0;
    assign pe_3_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_5_go =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? 1'd1 : 1'd0;
    assign pe_3_5_left =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? left_3_5_out : 32'd0;
    assign pe_3_5_top =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? top_3_5_out : 32'd0;
    assign pe_3_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_6_go =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? 1'd1 : 1'd0;
    assign pe_3_6_left =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? left_3_6_out : 32'd0;
    assign pe_3_6_top =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? top_3_6_out : 32'd0;
    assign pe_3_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_7_go =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? 1'd1 : 1'd0;
    assign pe_3_7_left =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? left_3_7_out : 32'd0;
    assign pe_3_7_top =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? top_3_7_out : 32'd0;
    assign pe_3_8_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_8_go =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 1'd1 : 1'd0;
    assign pe_3_8_left =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? left_3_8_out : 32'd0;
    assign pe_3_8_top =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? top_3_8_out : 32'd0;
    assign pe_3_9_clk =
     1'b1 ? clk : 1'd0;
    assign pe_3_9_go =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 1'd1 : 1'd0;
    assign pe_3_9_left =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? left_3_9_out : 32'd0;
    assign pe_3_9_top =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? top_3_9_out : 32'd0;
    assign pe_4_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_0_go =
     fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? 1'd1 : 1'd0;
    assign pe_4_0_left =
     fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? left_4_0_out : 32'd0;
    assign pe_4_0_top =
     fsm10_out < 3'd5 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? top_4_0_out : 32'd0;
    assign pe_4_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_1_go =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? 1'd1 : 1'd0;
    assign pe_4_1_left =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? left_4_1_out : 32'd0;
    assign pe_4_1_top =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? top_4_1_out : 32'd0;
    assign pe_4_10_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_10_go =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign pe_4_10_left =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? left_4_10_out : 32'd0;
    assign pe_4_10_top =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? top_4_10_out : 32'd0;
    assign pe_4_11_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_11_go =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 1'd1 : 1'd0;
    assign pe_4_11_left =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? left_4_11_out : 32'd0;
    assign pe_4_11_top =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? top_4_11_out : 32'd0;
    assign pe_4_12_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_12_go =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? 1'd1 : 1'd0;
    assign pe_4_12_left =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? left_4_12_out : 32'd0;
    assign pe_4_12_top =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? top_4_12_out : 32'd0;
    assign pe_4_13_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_13_go =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? 1'd1 : 1'd0;
    assign pe_4_13_left =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? left_4_13_out : 32'd0;
    assign pe_4_13_top =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? top_4_13_out : 32'd0;
    assign pe_4_14_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_14_go =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? 1'd1 : 1'd0;
    assign pe_4_14_left =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? left_4_14_out : 32'd0;
    assign pe_4_14_top =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? top_4_14_out : 32'd0;
    assign pe_4_15_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_15_go =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? 1'd1 : 1'd0;
    assign pe_4_15_left =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? left_4_15_out : 32'd0;
    assign pe_4_15_top =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? top_4_15_out : 32'd0;
    assign pe_4_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_2_go =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? 1'd1 : 1'd0;
    assign pe_4_2_left =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? left_4_2_out : 32'd0;
    assign pe_4_2_top =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? top_4_2_out : 32'd0;
    assign pe_4_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_3_go =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? 1'd1 : 1'd0;
    assign pe_4_3_left =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? left_4_3_out : 32'd0;
    assign pe_4_3_top =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? top_4_3_out : 32'd0;
    assign pe_4_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_4_go =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? 1'd1 : 1'd0;
    assign pe_4_4_left =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? left_4_4_out : 32'd0;
    assign pe_4_4_top =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? top_4_4_out : 32'd0;
    assign pe_4_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_5_go =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? 1'd1 : 1'd0;
    assign pe_4_5_left =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? left_4_5_out : 32'd0;
    assign pe_4_5_top =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? top_4_5_out : 32'd0;
    assign pe_4_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_6_go =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? 1'd1 : 1'd0;
    assign pe_4_6_left =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? left_4_6_out : 32'd0;
    assign pe_4_6_top =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? top_4_6_out : 32'd0;
    assign pe_4_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_7_go =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 1'd1 : 1'd0;
    assign pe_4_7_left =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? left_4_7_out : 32'd0;
    assign pe_4_7_top =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? top_4_7_out : 32'd0;
    assign pe_4_8_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_8_go =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 1'd1 : 1'd0;
    assign pe_4_8_left =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? left_4_8_out : 32'd0;
    assign pe_4_8_top =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? top_4_8_out : 32'd0;
    assign pe_4_9_clk =
     1'b1 ? clk : 1'd0;
    assign pe_4_9_go =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 1'd1 : 1'd0;
    assign pe_4_9_left =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? left_4_9_out : 32'd0;
    assign pe_4_9_top =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? top_4_9_out : 32'd0;
    assign pe_5_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_0_go =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? 1'd1 : 1'd0;
    assign pe_5_0_left =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? left_5_0_out : 32'd0;
    assign pe_5_0_top =
     fsm12_out < 3'd5 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? top_5_0_out : 32'd0;
    assign pe_5_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_1_go =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? 1'd1 : 1'd0;
    assign pe_5_1_left =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? left_5_1_out : 32'd0;
    assign pe_5_1_top =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? top_5_1_out : 32'd0;
    assign pe_5_10_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_10_go =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 1'd1 : 1'd0;
    assign pe_5_10_left =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? left_5_10_out : 32'd0;
    assign pe_5_10_top =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? top_5_10_out : 32'd0;
    assign pe_5_11_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_11_go =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? 1'd1 : 1'd0;
    assign pe_5_11_left =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? left_5_11_out : 32'd0;
    assign pe_5_11_top =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? top_5_11_out : 32'd0;
    assign pe_5_12_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_12_go =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? 1'd1 : 1'd0;
    assign pe_5_12_left =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? left_5_12_out : 32'd0;
    assign pe_5_12_top =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? top_5_12_out : 32'd0;
    assign pe_5_13_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_13_go =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? 1'd1 : 1'd0;
    assign pe_5_13_left =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? left_5_13_out : 32'd0;
    assign pe_5_13_top =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? top_5_13_out : 32'd0;
    assign pe_5_14_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_14_go =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? 1'd1 : 1'd0;
    assign pe_5_14_left =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? left_5_14_out : 32'd0;
    assign pe_5_14_top =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? top_5_14_out : 32'd0;
    assign pe_5_15_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_15_go =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? 1'd1 : 1'd0;
    assign pe_5_15_left =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? left_5_15_out : 32'd0;
    assign pe_5_15_top =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? top_5_15_out : 32'd0;
    assign pe_5_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_2_go =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? 1'd1 : 1'd0;
    assign pe_5_2_left =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? left_5_2_out : 32'd0;
    assign pe_5_2_top =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? top_5_2_out : 32'd0;
    assign pe_5_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_3_go =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? 1'd1 : 1'd0;
    assign pe_5_3_left =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? left_5_3_out : 32'd0;
    assign pe_5_3_top =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? top_5_3_out : 32'd0;
    assign pe_5_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_4_go =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? 1'd1 : 1'd0;
    assign pe_5_4_left =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? left_5_4_out : 32'd0;
    assign pe_5_4_top =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? top_5_4_out : 32'd0;
    assign pe_5_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_5_go =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? 1'd1 : 1'd0;
    assign pe_5_5_left =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? left_5_5_out : 32'd0;
    assign pe_5_5_top =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? top_5_5_out : 32'd0;
    assign pe_5_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_6_go =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 1'd1 : 1'd0;
    assign pe_5_6_left =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? left_5_6_out : 32'd0;
    assign pe_5_6_top =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? top_5_6_out : 32'd0;
    assign pe_5_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_7_go =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 1'd1 : 1'd0;
    assign pe_5_7_left =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? left_5_7_out : 32'd0;
    assign pe_5_7_top =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? top_5_7_out : 32'd0;
    assign pe_5_8_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_8_go =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 1'd1 : 1'd0;
    assign pe_5_8_left =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? left_5_8_out : 32'd0;
    assign pe_5_8_top =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? top_5_8_out : 32'd0;
    assign pe_5_9_clk =
     1'b1 ? clk : 1'd0;
    assign pe_5_9_go =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign pe_5_9_left =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? left_5_9_out : 32'd0;
    assign pe_5_9_top =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? top_5_9_out : 32'd0;
    assign pe_6_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_0_go =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? 1'd1 : 1'd0;
    assign pe_6_0_left =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? left_6_0_out : 32'd0;
    assign pe_6_0_top =
     fsm14_out < 3'd5 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? top_6_0_out : 32'd0;
    assign pe_6_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_1_go =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? 1'd1 : 1'd0;
    assign pe_6_1_left =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? left_6_1_out : 32'd0;
    assign pe_6_1_top =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? top_6_1_out : 32'd0;
    assign pe_6_10_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_10_go =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? 1'd1 : 1'd0;
    assign pe_6_10_left =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? left_6_10_out : 32'd0;
    assign pe_6_10_top =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? top_6_10_out : 32'd0;
    assign pe_6_11_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_11_go =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? 1'd1 : 1'd0;
    assign pe_6_11_left =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? left_6_11_out : 32'd0;
    assign pe_6_11_top =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? top_6_11_out : 32'd0;
    assign pe_6_12_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_12_go =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? 1'd1 : 1'd0;
    assign pe_6_12_left =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? left_6_12_out : 32'd0;
    assign pe_6_12_top =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? top_6_12_out : 32'd0;
    assign pe_6_13_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_13_go =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? 1'd1 : 1'd0;
    assign pe_6_13_left =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? left_6_13_out : 32'd0;
    assign pe_6_13_top =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? top_6_13_out : 32'd0;
    assign pe_6_14_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_14_go =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? 1'd1 : 1'd0;
    assign pe_6_14_left =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? left_6_14_out : 32'd0;
    assign pe_6_14_top =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? top_6_14_out : 32'd0;
    assign pe_6_15_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_15_go =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? 1'd1 : 1'd0;
    assign pe_6_15_left =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? left_6_15_out : 32'd0;
    assign pe_6_15_top =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? top_6_15_out : 32'd0;
    assign pe_6_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_2_go =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? 1'd1 : 1'd0;
    assign pe_6_2_left =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? left_6_2_out : 32'd0;
    assign pe_6_2_top =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? top_6_2_out : 32'd0;
    assign pe_6_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_3_go =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? 1'd1 : 1'd0;
    assign pe_6_3_left =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? left_6_3_out : 32'd0;
    assign pe_6_3_top =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? top_6_3_out : 32'd0;
    assign pe_6_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_4_go =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? 1'd1 : 1'd0;
    assign pe_6_4_left =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? left_6_4_out : 32'd0;
    assign pe_6_4_top =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? top_6_4_out : 32'd0;
    assign pe_6_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_5_go =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 1'd1 : 1'd0;
    assign pe_6_5_left =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? left_6_5_out : 32'd0;
    assign pe_6_5_top =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? top_6_5_out : 32'd0;
    assign pe_6_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_6_go =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 1'd1 : 1'd0;
    assign pe_6_6_left =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? left_6_6_out : 32'd0;
    assign pe_6_6_top =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? top_6_6_out : 32'd0;
    assign pe_6_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_7_go =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 1'd1 : 1'd0;
    assign pe_6_7_left =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? left_6_7_out : 32'd0;
    assign pe_6_7_top =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? top_6_7_out : 32'd0;
    assign pe_6_8_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_8_go =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign pe_6_8_left =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? left_6_8_out : 32'd0;
    assign pe_6_8_top =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? top_6_8_out : 32'd0;
    assign pe_6_9_clk =
     1'b1 ? clk : 1'd0;
    assign pe_6_9_go =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 1'd1 : 1'd0;
    assign pe_6_9_left =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? left_6_9_out : 32'd0;
    assign pe_6_9_top =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? top_6_9_out : 32'd0;
    assign pe_7_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_0_go =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? 1'd1 : 1'd0;
    assign pe_7_0_left =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? left_7_0_out : 32'd0;
    assign pe_7_0_top =
     fsm16_out < 3'd5 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? top_7_0_out : 32'd0;
    assign pe_7_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_1_go =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? 1'd1 : 1'd0;
    assign pe_7_1_left =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? left_7_1_out : 32'd0;
    assign pe_7_1_top =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? top_7_1_out : 32'd0;
    assign pe_7_10_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_10_go =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? 1'd1 : 1'd0;
    assign pe_7_10_left =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? left_7_10_out : 32'd0;
    assign pe_7_10_top =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? top_7_10_out : 32'd0;
    assign pe_7_11_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_11_go =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? 1'd1 : 1'd0;
    assign pe_7_11_left =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? left_7_11_out : 32'd0;
    assign pe_7_11_top =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? top_7_11_out : 32'd0;
    assign pe_7_12_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_12_go =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? 1'd1 : 1'd0;
    assign pe_7_12_left =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? left_7_12_out : 32'd0;
    assign pe_7_12_top =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? top_7_12_out : 32'd0;
    assign pe_7_13_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_13_go =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? 1'd1 : 1'd0;
    assign pe_7_13_left =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? left_7_13_out : 32'd0;
    assign pe_7_13_top =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? top_7_13_out : 32'd0;
    assign pe_7_14_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_14_go =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? 1'd1 : 1'd0;
    assign pe_7_14_left =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? left_7_14_out : 32'd0;
    assign pe_7_14_top =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? top_7_14_out : 32'd0;
    assign pe_7_15_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_15_go =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? 1'd1 : 1'd0;
    assign pe_7_15_left =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? left_7_15_out : 32'd0;
    assign pe_7_15_top =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? top_7_15_out : 32'd0;
    assign pe_7_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_2_go =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? 1'd1 : 1'd0;
    assign pe_7_2_left =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? left_7_2_out : 32'd0;
    assign pe_7_2_top =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? top_7_2_out : 32'd0;
    assign pe_7_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_3_go =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? 1'd1 : 1'd0;
    assign pe_7_3_left =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? left_7_3_out : 32'd0;
    assign pe_7_3_top =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? top_7_3_out : 32'd0;
    assign pe_7_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_4_go =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 1'd1 : 1'd0;
    assign pe_7_4_left =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? left_7_4_out : 32'd0;
    assign pe_7_4_top =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? top_7_4_out : 32'd0;
    assign pe_7_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_5_go =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 1'd1 : 1'd0;
    assign pe_7_5_left =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? left_7_5_out : 32'd0;
    assign pe_7_5_top =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? top_7_5_out : 32'd0;
    assign pe_7_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_6_go =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 1'd1 : 1'd0;
    assign pe_7_6_left =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? left_7_6_out : 32'd0;
    assign pe_7_6_top =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? top_7_6_out : 32'd0;
    assign pe_7_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_7_go =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign pe_7_7_left =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? left_7_7_out : 32'd0;
    assign pe_7_7_top =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? top_7_7_out : 32'd0;
    assign pe_7_8_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_8_go =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 1'd1 : 1'd0;
    assign pe_7_8_left =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? left_7_8_out : 32'd0;
    assign pe_7_8_top =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? top_7_8_out : 32'd0;
    assign pe_7_9_clk =
     1'b1 ? clk : 1'd0;
    assign pe_7_9_go =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? 1'd1 : 1'd0;
    assign pe_7_9_left =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? left_7_9_out : 32'd0;
    assign pe_7_9_top =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? top_7_9_out : 32'd0;
    assign pe_8_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_8_0_go =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? 1'd1 : 1'd0;
    assign pe_8_0_left =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? left_8_0_out : 32'd0;
    assign pe_8_0_top =
     fsm18_out < 3'd5 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? top_8_0_out : 32'd0;
    assign pe_8_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_8_1_go =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? 1'd1 : 1'd0;
    assign pe_8_1_left =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? left_8_1_out : 32'd0;
    assign pe_8_1_top =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? top_8_1_out : 32'd0;
    assign pe_8_10_clk =
     1'b1 ? clk : 1'd0;
    assign pe_8_10_go =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? 1'd1 : 1'd0;
    assign pe_8_10_left =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? left_8_10_out : 32'd0;
    assign pe_8_10_top =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? top_8_10_out : 32'd0;
    assign pe_8_11_clk =
     1'b1 ? clk : 1'd0;
    assign pe_8_11_go =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? 1'd1 : 1'd0;
    assign pe_8_11_left =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? left_8_11_out : 32'd0;
    assign pe_8_11_top =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? top_8_11_out : 32'd0;
    assign pe_8_12_clk =
     1'b1 ? clk : 1'd0;
    assign pe_8_12_go =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? 1'd1 : 1'd0;
    assign pe_8_12_left =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? left_8_12_out : 32'd0;
    assign pe_8_12_top =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? top_8_12_out : 32'd0;
    assign pe_8_13_clk =
     1'b1 ? clk : 1'd0;
    assign pe_8_13_go =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? 1'd1 : 1'd0;
    assign pe_8_13_left =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? left_8_13_out : 32'd0;
    assign pe_8_13_top =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? top_8_13_out : 32'd0;
    assign pe_8_14_clk =
     1'b1 ? clk : 1'd0;
    assign pe_8_14_go =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? 1'd1 : 1'd0;
    assign pe_8_14_left =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? left_8_14_out : 32'd0;
    assign pe_8_14_top =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? top_8_14_out : 32'd0;
    assign pe_8_15_clk =
     1'b1 ? clk : 1'd0;
    assign pe_8_15_go =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? 1'd1 : 1'd0;
    assign pe_8_15_left =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? left_8_15_out : 32'd0;
    assign pe_8_15_top =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? top_8_15_out : 32'd0;
    assign pe_8_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_8_2_go =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? 1'd1 : 1'd0;
    assign pe_8_2_left =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? left_8_2_out : 32'd0;
    assign pe_8_2_top =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? top_8_2_out : 32'd0;
    assign pe_8_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_8_3_go =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 1'd1 : 1'd0;
    assign pe_8_3_left =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? left_8_3_out : 32'd0;
    assign pe_8_3_top =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? top_8_3_out : 32'd0;
    assign pe_8_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_8_4_go =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 1'd1 : 1'd0;
    assign pe_8_4_left =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? left_8_4_out : 32'd0;
    assign pe_8_4_top =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? top_8_4_out : 32'd0;
    assign pe_8_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_8_5_go =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 1'd1 : 1'd0;
    assign pe_8_5_left =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? left_8_5_out : 32'd0;
    assign pe_8_5_top =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? top_8_5_out : 32'd0;
    assign pe_8_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_8_6_go =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign pe_8_6_left =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? left_8_6_out : 32'd0;
    assign pe_8_6_top =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? top_8_6_out : 32'd0;
    assign pe_8_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_8_7_go =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 1'd1 : 1'd0;
    assign pe_8_7_left =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? left_8_7_out : 32'd0;
    assign pe_8_7_top =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? top_8_7_out : 32'd0;
    assign pe_8_8_clk =
     1'b1 ? clk : 1'd0;
    assign pe_8_8_go =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? 1'd1 : 1'd0;
    assign pe_8_8_left =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? left_8_8_out : 32'd0;
    assign pe_8_8_top =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? top_8_8_out : 32'd0;
    assign pe_8_9_clk =
     1'b1 ? clk : 1'd0;
    assign pe_8_9_go =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? 1'd1 : 1'd0;
    assign pe_8_9_left =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? left_8_9_out : 32'd0;
    assign pe_8_9_top =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? top_8_9_out : 32'd0;
    assign pe_9_0_clk =
     1'b1 ? clk : 1'd0;
    assign pe_9_0_go =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? 1'd1 : 1'd0;
    assign pe_9_0_left =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? left_9_0_out : 32'd0;
    assign pe_9_0_top =
     fsm20_out < 3'd5 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? top_9_0_out : 32'd0;
    assign pe_9_1_clk =
     1'b1 ? clk : 1'd0;
    assign pe_9_1_go =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? 1'd1 : 1'd0;
    assign pe_9_1_left =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? left_9_1_out : 32'd0;
    assign pe_9_1_top =
     fsm22_out < 3'd5 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? top_9_1_out : 32'd0;
    assign pe_9_10_clk =
     1'b1 ? clk : 1'd0;
    assign pe_9_10_go =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? 1'd1 : 1'd0;
    assign pe_9_10_left =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? left_9_10_out : 32'd0;
    assign pe_9_10_top =
     fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go ? top_9_10_out : 32'd0;
    assign pe_9_11_clk =
     1'b1 ? clk : 1'd0;
    assign pe_9_11_go =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? 1'd1 : 1'd0;
    assign pe_9_11_left =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? left_9_11_out : 32'd0;
    assign pe_9_11_top =
     fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go ? top_9_11_out : 32'd0;
    assign pe_9_12_clk =
     1'b1 ? clk : 1'd0;
    assign pe_9_12_go =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? 1'd1 : 1'd0;
    assign pe_9_12_left =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? left_9_12_out : 32'd0;
    assign pe_9_12_top =
     fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go ? top_9_12_out : 32'd0;
    assign pe_9_13_clk =
     1'b1 ? clk : 1'd0;
    assign pe_9_13_go =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? 1'd1 : 1'd0;
    assign pe_9_13_left =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? left_9_13_out : 32'd0;
    assign pe_9_13_top =
     fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go ? top_9_13_out : 32'd0;
    assign pe_9_14_clk =
     1'b1 ? clk : 1'd0;
    assign pe_9_14_go =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? 1'd1 : 1'd0;
    assign pe_9_14_left =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? left_9_14_out : 32'd0;
    assign pe_9_14_top =
     fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go ? top_9_14_out : 32'd0;
    assign pe_9_15_clk =
     1'b1 ? clk : 1'd0;
    assign pe_9_15_go =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? 1'd1 : 1'd0;
    assign pe_9_15_left =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? left_9_15_out : 32'd0;
    assign pe_9_15_top =
     fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go | fsm70_out < 3'd5 & fsm92_out >= 10'd207 & fsm92_out < 10'd212 & go | fsm72_out < 3'd5 & fsm92_out >= 10'd213 & fsm92_out < 10'd218 & go | fsm74_out < 3'd5 & fsm92_out >= 10'd219 & fsm92_out < 10'd224 & go | fsm76_out < 3'd5 & fsm92_out >= 10'd225 & fsm92_out < 10'd230 & go | fsm78_out < 3'd5 & fsm92_out >= 10'd231 & fsm92_out < 10'd236 & go | fsm80_out < 3'd5 & fsm92_out >= 10'd237 & fsm92_out < 10'd242 & go ? top_9_15_out : 32'd0;
    assign pe_9_2_clk =
     1'b1 ? clk : 1'd0;
    assign pe_9_2_go =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 1'd1 : 1'd0;
    assign pe_9_2_left =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? left_9_2_out : 32'd0;
    assign pe_9_2_top =
     fsm24_out < 3'd5 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? top_9_2_out : 32'd0;
    assign pe_9_3_clk =
     1'b1 ? clk : 1'd0;
    assign pe_9_3_go =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 1'd1 : 1'd0;
    assign pe_9_3_left =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? left_9_3_out : 32'd0;
    assign pe_9_3_top =
     fsm26_out < 3'd5 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? top_9_3_out : 32'd0;
    assign pe_9_4_clk =
     1'b1 ? clk : 1'd0;
    assign pe_9_4_go =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 1'd1 : 1'd0;
    assign pe_9_4_left =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? left_9_4_out : 32'd0;
    assign pe_9_4_top =
     fsm28_out < 3'd5 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? top_9_4_out : 32'd0;
    assign pe_9_5_clk =
     1'b1 ? clk : 1'd0;
    assign pe_9_5_go =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign pe_9_5_left =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? left_9_5_out : 32'd0;
    assign pe_9_5_top =
     fsm30_out < 3'd5 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? top_9_5_out : 32'd0;
    assign pe_9_6_clk =
     1'b1 ? clk : 1'd0;
    assign pe_9_6_go =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? 1'd1 : 1'd0;
    assign pe_9_6_left =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? left_9_6_out : 32'd0;
    assign pe_9_6_top =
     fsm32_out < 3'd5 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go ? top_9_6_out : 32'd0;
    assign pe_9_7_clk =
     1'b1 ? clk : 1'd0;
    assign pe_9_7_go =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? 1'd1 : 1'd0;
    assign pe_9_7_left =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? left_9_7_out : 32'd0;
    assign pe_9_7_top =
     fsm34_out < 3'd5 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go ? top_9_7_out : 32'd0;
    assign pe_9_8_clk =
     1'b1 ? clk : 1'd0;
    assign pe_9_8_go =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? 1'd1 : 1'd0;
    assign pe_9_8_left =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? left_9_8_out : 32'd0;
    assign pe_9_8_top =
     fsm36_out < 3'd5 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go ? top_9_8_out : 32'd0;
    assign pe_9_9_clk =
     1'b1 ? clk : 1'd0;
    assign pe_9_9_go =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? 1'd1 : 1'd0;
    assign pe_9_9_left =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? left_9_9_out : 32'd0;
    assign pe_9_9_top =
     fsm38_out < 3'd5 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd5 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd5 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd5 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd5 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd5 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd5 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd5 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd5 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd5 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd5 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd5 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go | fsm62_out < 3'd5 & fsm92_out >= 10'd183 & fsm92_out < 10'd188 & go | fsm64_out < 3'd5 & fsm92_out >= 10'd189 & fsm92_out < 10'd194 & go | fsm66_out < 3'd5 & fsm92_out >= 10'd195 & fsm92_out < 10'd200 & go | fsm68_out < 3'd5 & fsm92_out >= 10'd201 & fsm92_out < 10'd206 & go ? top_9_9_out : 32'd0;
    assign t0_add_left =
     fsm0_out < 1'd1 & fsm92_out == 10'd1 & go | fsm2_out < 3'd1 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go ? 5'd1 : 5'd0;
    assign t0_add_right =
     fsm0_out < 1'd1 & fsm92_out == 10'd1 & go | fsm2_out < 3'd1 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go ? t0_idx_out : 5'd0;
    assign t0_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t0_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm0_out < 1'd1 & fsm92_out == 10'd1 & go | fsm2_out < 3'd1 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go ? t0_add_out : 5'd0;
    assign t0_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm0_out < 1'd1 & fsm92_out == 10'd1 & go | fsm2_out < 3'd1 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go ? 1'd1 : 1'd0;
    assign t10_add_left =
     fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? 5'd1 : 5'd0;
    assign t10_add_right =
     fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? t10_idx_out : 5'd0;
    assign t10_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t10_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? t10_add_out : 5'd0;
    assign t10_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go ? 1'd1 : 1'd0;
    assign t11_add_left =
     fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? 5'd1 : 5'd0;
    assign t11_add_right =
     fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? t11_idx_out : 5'd0;
    assign t11_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t11_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? t11_add_out : 5'd0;
    assign t11_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go ? 1'd1 : 1'd0;
    assign t12_add_left =
     fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 5'd1 : 5'd0;
    assign t12_add_right =
     fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? t12_idx_out : 5'd0;
    assign t12_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t12_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? t12_add_out : 5'd0;
    assign t12_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go ? 1'd1 : 1'd0;
    assign t13_add_left =
     fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 5'd1 : 5'd0;
    assign t13_add_right =
     fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? t13_idx_out : 5'd0;
    assign t13_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t13_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? t13_add_out : 5'd0;
    assign t13_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go ? 1'd1 : 1'd0;
    assign t14_add_left =
     fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd1 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 5'd1 : 5'd0;
    assign t14_add_right =
     fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd1 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? t14_idx_out : 5'd0;
    assign t14_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t14_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd1 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? t14_add_out : 5'd0;
    assign t14_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd1 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go ? 1'd1 : 1'd0;
    assign t15_add_left =
     fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd1 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd1 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 5'd1 : 5'd0;
    assign t15_add_right =
     fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd1 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd1 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? t15_idx_out : 5'd0;
    assign t15_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t15_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd1 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd1 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? t15_add_out : 5'd0;
    assign t15_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go | fsm50_out < 3'd1 & fsm92_out >= 10'd147 & fsm92_out < 10'd152 & go | fsm52_out < 3'd1 & fsm92_out >= 10'd153 & fsm92_out < 10'd158 & go | fsm54_out < 3'd1 & fsm92_out >= 10'd159 & fsm92_out < 10'd164 & go | fsm56_out < 3'd1 & fsm92_out >= 10'd165 & fsm92_out < 10'd170 & go | fsm58_out < 3'd1 & fsm92_out >= 10'd171 & fsm92_out < 10'd176 & go | fsm60_out < 3'd1 & fsm92_out >= 10'd177 & fsm92_out < 10'd182 & go ? 1'd1 : 1'd0;
    assign t1_add_left =
     fsm2_out < 3'd1 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go ? 5'd1 : 5'd0;
    assign t1_add_right =
     fsm2_out < 3'd1 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go ? t1_idx_out : 5'd0;
    assign t1_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t1_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm2_out < 3'd1 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go ? t1_add_out : 5'd0;
    assign t1_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm2_out < 3'd1 & fsm92_out >= 10'd3 & fsm92_out < 10'd8 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go ? 1'd1 : 1'd0;
    assign t2_add_left =
     fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? 5'd1 : 5'd0;
    assign t2_add_right =
     fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? t2_idx_out : 5'd0;
    assign t2_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t2_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? t2_add_out : 5'd0;
    assign t2_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm4_out < 3'd1 & fsm92_out >= 10'd9 & fsm92_out < 10'd14 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go ? 1'd1 : 1'd0;
    assign t3_add_left =
     fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? 5'd1 : 5'd0;
    assign t3_add_right =
     fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? t3_idx_out : 5'd0;
    assign t3_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t3_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? t3_add_out : 5'd0;
    assign t3_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm6_out < 3'd1 & fsm92_out >= 10'd15 & fsm92_out < 10'd20 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go ? 1'd1 : 1'd0;
    assign t4_add_left =
     fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? 5'd1 : 5'd0;
    assign t4_add_right =
     fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? t4_idx_out : 5'd0;
    assign t4_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t4_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? t4_add_out : 5'd0;
    assign t4_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm8_out < 3'd1 & fsm92_out >= 10'd21 & fsm92_out < 10'd26 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go ? 1'd1 : 1'd0;
    assign t5_add_left =
     fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? 5'd1 : 5'd0;
    assign t5_add_right =
     fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? t5_idx_out : 5'd0;
    assign t5_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t5_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? t5_add_out : 5'd0;
    assign t5_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm10_out < 3'd1 & fsm92_out >= 10'd27 & fsm92_out < 10'd32 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go ? 1'd1 : 1'd0;
    assign t6_add_left =
     fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? 5'd1 : 5'd0;
    assign t6_add_right =
     fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? t6_idx_out : 5'd0;
    assign t6_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t6_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? t6_add_out : 5'd0;
    assign t6_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm12_out < 3'd1 & fsm92_out >= 10'd33 & fsm92_out < 10'd38 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go ? 1'd1 : 1'd0;
    assign t7_add_left =
     fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? 5'd1 : 5'd0;
    assign t7_add_right =
     fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? t7_idx_out : 5'd0;
    assign t7_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t7_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? t7_add_out : 5'd0;
    assign t7_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm14_out < 3'd1 & fsm92_out >= 10'd39 & fsm92_out < 10'd44 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go ? 1'd1 : 1'd0;
    assign t8_add_left =
     fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? 5'd1 : 5'd0;
    assign t8_add_right =
     fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? t8_idx_out : 5'd0;
    assign t8_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t8_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? t8_add_out : 5'd0;
    assign t8_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm16_out < 3'd1 & fsm92_out >= 10'd45 & fsm92_out < 10'd50 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go ? 1'd1 : 1'd0;
    assign t9_add_left =
     fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? 5'd1 : 5'd0;
    assign t9_add_right =
     fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? t9_idx_out : 5'd0;
    assign t9_idx_clk =
     1'b1 ? clk : 1'd0;
    assign t9_idx_in =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go ? 5'd31 :
     fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? t9_add_out : 5'd0;
    assign t9_idx_write_en =
     fsm_out < 1'd1 & fsm92_out == 10'd0 & go | fsm18_out < 3'd1 & fsm92_out >= 10'd51 & fsm92_out < 10'd56 & go | fsm20_out < 3'd1 & fsm92_out >= 10'd57 & fsm92_out < 10'd62 & go | fsm22_out < 3'd1 & fsm92_out >= 10'd63 & fsm92_out < 10'd68 & go | fsm24_out < 3'd1 & fsm92_out >= 10'd69 & fsm92_out < 10'd74 & go | fsm26_out < 3'd1 & fsm92_out >= 10'd75 & fsm92_out < 10'd80 & go | fsm28_out < 3'd1 & fsm92_out >= 10'd81 & fsm92_out < 10'd86 & go | fsm30_out < 3'd1 & fsm92_out >= 10'd87 & fsm92_out < 10'd92 & go | fsm32_out < 3'd1 & fsm92_out >= 10'd93 & fsm92_out < 10'd98 & go | fsm34_out < 3'd1 & fsm92_out >= 10'd99 & fsm92_out < 10'd104 & go | fsm36_out < 3'd1 & fsm92_out >= 10'd105 & fsm92_out < 10'd110 & go | fsm38_out < 3'd1 & fsm92_out >= 10'd111 & fsm92_out < 10'd116 & go | fsm40_out < 3'd1 & fsm92_out >= 10'd117 & fsm92_out < 10'd122 & go | fsm42_out < 3'd1 & fsm92_out >= 10'd123 & fsm92_out < 10'd128 & go | fsm44_out < 3'd1 & fsm92_out >= 10'd129 & fsm92_out < 10'd134 & go | fsm46_out < 3'd1 & fsm92_out >= 10'd135 & fsm92_out < 10'd140 & go | fsm48_out < 3'd1 & fsm92_out >= 10'd141 & fsm92_out < 10'd146 & go ? 1'd1 : 1'd0;
    assign top_0_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_0_in =
     fsm1_out < 1'd1 & fsm92_out == 10'd2 & go | fsm3_out < 1'd1 & fsm92_out == 10'd8 & go | fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go ? t0_read_data : 32'd0;
    assign top_0_0_write_en =
     fsm1_out < 1'd1 & fsm92_out == 10'd2 & go | fsm3_out < 1'd1 & fsm92_out == 10'd8 & go | fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go ? 1'd1 : 1'd0;
    assign top_0_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_1_in =
     fsm3_out < 1'd1 & fsm92_out == 10'd8 & go | fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go ? t1_read_data : 32'd0;
    assign top_0_1_write_en =
     fsm3_out < 1'd1 & fsm92_out == 10'd8 & go | fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go ? 1'd1 : 1'd0;
    assign top_0_10_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_10_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? t10_read_data : 32'd0;
    assign top_0_10_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign top_0_11_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_11_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? t11_read_data : 32'd0;
    assign top_0_11_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign top_0_12_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_12_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? t12_read_data : 32'd0;
    assign top_0_12_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign top_0_13_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_13_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? t13_read_data : 32'd0;
    assign top_0_13_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign top_0_14_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_14_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? t14_read_data : 32'd0;
    assign top_0_14_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign top_0_15_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_15_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? t15_read_data : 32'd0;
    assign top_0_15_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign top_0_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_2_in =
     fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go ? t2_read_data : 32'd0;
    assign top_0_2_write_en =
     fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go ? 1'd1 : 1'd0;
    assign top_0_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_3_in =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? t3_read_data : 32'd0;
    assign top_0_3_write_en =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? 1'd1 : 1'd0;
    assign top_0_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_4_in =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? t4_read_data : 32'd0;
    assign top_0_4_write_en =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? 1'd1 : 1'd0;
    assign top_0_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_5_in =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? t5_read_data : 32'd0;
    assign top_0_5_write_en =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? 1'd1 : 1'd0;
    assign top_0_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_6_in =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? t6_read_data : 32'd0;
    assign top_0_6_write_en =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? 1'd1 : 1'd0;
    assign top_0_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_7_in =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? t7_read_data : 32'd0;
    assign top_0_7_write_en =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign top_0_8_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_8_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? t8_read_data : 32'd0;
    assign top_0_8_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign top_0_9_clk =
     1'b1 ? clk : 1'd0;
    assign top_0_9_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? t9_read_data : 32'd0;
    assign top_0_9_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign top_10_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_10_0_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? top_9_0_out : 32'd0;
    assign top_10_0_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign top_10_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_10_1_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? top_9_1_out : 32'd0;
    assign top_10_1_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign top_10_10_clk =
     1'b1 ? clk : 1'd0;
    assign top_10_10_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? top_9_10_out : 32'd0;
    assign top_10_10_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign top_10_11_clk =
     1'b1 ? clk : 1'd0;
    assign top_10_11_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? top_9_11_out : 32'd0;
    assign top_10_11_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign top_10_12_clk =
     1'b1 ? clk : 1'd0;
    assign top_10_12_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? top_9_12_out : 32'd0;
    assign top_10_12_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign top_10_13_clk =
     1'b1 ? clk : 1'd0;
    assign top_10_13_in =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? top_9_13_out : 32'd0;
    assign top_10_13_write_en =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign top_10_14_clk =
     1'b1 ? clk : 1'd0;
    assign top_10_14_in =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? top_9_14_out : 32'd0;
    assign top_10_14_write_en =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? 1'd1 : 1'd0;
    assign top_10_15_clk =
     1'b1 ? clk : 1'd0;
    assign top_10_15_in =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? top_9_15_out : 32'd0;
    assign top_10_15_write_en =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? 1'd1 : 1'd0;
    assign top_10_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_10_2_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? top_9_2_out : 32'd0;
    assign top_10_2_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign top_10_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_10_3_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? top_9_3_out : 32'd0;
    assign top_10_3_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign top_10_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_10_4_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? top_9_4_out : 32'd0;
    assign top_10_4_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign top_10_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_10_5_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? top_9_5_out : 32'd0;
    assign top_10_5_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign top_10_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_10_6_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? top_9_6_out : 32'd0;
    assign top_10_6_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign top_10_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_10_7_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? top_9_7_out : 32'd0;
    assign top_10_7_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign top_10_8_clk =
     1'b1 ? clk : 1'd0;
    assign top_10_8_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? top_9_8_out : 32'd0;
    assign top_10_8_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign top_10_9_clk =
     1'b1 ? clk : 1'd0;
    assign top_10_9_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? top_9_9_out : 32'd0;
    assign top_10_9_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign top_11_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_11_0_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? top_10_0_out : 32'd0;
    assign top_11_0_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign top_11_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_11_1_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? top_10_1_out : 32'd0;
    assign top_11_1_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign top_11_10_clk =
     1'b1 ? clk : 1'd0;
    assign top_11_10_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? top_10_10_out : 32'd0;
    assign top_11_10_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign top_11_11_clk =
     1'b1 ? clk : 1'd0;
    assign top_11_11_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? top_10_11_out : 32'd0;
    assign top_11_11_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign top_11_12_clk =
     1'b1 ? clk : 1'd0;
    assign top_11_12_in =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? top_10_12_out : 32'd0;
    assign top_11_12_write_en =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign top_11_13_clk =
     1'b1 ? clk : 1'd0;
    assign top_11_13_in =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? top_10_13_out : 32'd0;
    assign top_11_13_write_en =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? 1'd1 : 1'd0;
    assign top_11_14_clk =
     1'b1 ? clk : 1'd0;
    assign top_11_14_in =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? top_10_14_out : 32'd0;
    assign top_11_14_write_en =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? 1'd1 : 1'd0;
    assign top_11_15_clk =
     1'b1 ? clk : 1'd0;
    assign top_11_15_in =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? top_10_15_out : 32'd0;
    assign top_11_15_write_en =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? 1'd1 : 1'd0;
    assign top_11_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_11_2_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? top_10_2_out : 32'd0;
    assign top_11_2_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign top_11_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_11_3_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? top_10_3_out : 32'd0;
    assign top_11_3_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign top_11_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_11_4_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? top_10_4_out : 32'd0;
    assign top_11_4_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign top_11_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_11_5_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? top_10_5_out : 32'd0;
    assign top_11_5_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign top_11_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_11_6_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? top_10_6_out : 32'd0;
    assign top_11_6_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign top_11_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_11_7_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? top_10_7_out : 32'd0;
    assign top_11_7_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign top_11_8_clk =
     1'b1 ? clk : 1'd0;
    assign top_11_8_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? top_10_8_out : 32'd0;
    assign top_11_8_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign top_11_9_clk =
     1'b1 ? clk : 1'd0;
    assign top_11_9_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? top_10_9_out : 32'd0;
    assign top_11_9_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign top_12_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_12_0_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? top_11_0_out : 32'd0;
    assign top_12_0_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign top_12_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_12_1_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? top_11_1_out : 32'd0;
    assign top_12_1_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign top_12_10_clk =
     1'b1 ? clk : 1'd0;
    assign top_12_10_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? top_11_10_out : 32'd0;
    assign top_12_10_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign top_12_11_clk =
     1'b1 ? clk : 1'd0;
    assign top_12_11_in =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? top_11_11_out : 32'd0;
    assign top_12_11_write_en =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign top_12_12_clk =
     1'b1 ? clk : 1'd0;
    assign top_12_12_in =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? top_11_12_out : 32'd0;
    assign top_12_12_write_en =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? 1'd1 : 1'd0;
    assign top_12_13_clk =
     1'b1 ? clk : 1'd0;
    assign top_12_13_in =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? top_11_13_out : 32'd0;
    assign top_12_13_write_en =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? 1'd1 : 1'd0;
    assign top_12_14_clk =
     1'b1 ? clk : 1'd0;
    assign top_12_14_in =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? top_11_14_out : 32'd0;
    assign top_12_14_write_en =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? 1'd1 : 1'd0;
    assign top_12_15_clk =
     1'b1 ? clk : 1'd0;
    assign top_12_15_in =
     fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go ? top_11_15_out : 32'd0;
    assign top_12_15_write_en =
     fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go ? 1'd1 : 1'd0;
    assign top_12_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_12_2_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? top_11_2_out : 32'd0;
    assign top_12_2_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign top_12_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_12_3_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? top_11_3_out : 32'd0;
    assign top_12_3_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign top_12_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_12_4_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? top_11_4_out : 32'd0;
    assign top_12_4_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign top_12_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_12_5_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? top_11_5_out : 32'd0;
    assign top_12_5_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign top_12_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_12_6_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? top_11_6_out : 32'd0;
    assign top_12_6_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign top_12_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_12_7_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? top_11_7_out : 32'd0;
    assign top_12_7_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign top_12_8_clk =
     1'b1 ? clk : 1'd0;
    assign top_12_8_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? top_11_8_out : 32'd0;
    assign top_12_8_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign top_12_9_clk =
     1'b1 ? clk : 1'd0;
    assign top_12_9_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? top_11_9_out : 32'd0;
    assign top_12_9_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign top_13_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_13_0_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? top_12_0_out : 32'd0;
    assign top_13_0_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign top_13_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_13_1_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? top_12_1_out : 32'd0;
    assign top_13_1_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign top_13_10_clk =
     1'b1 ? clk : 1'd0;
    assign top_13_10_in =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? top_12_10_out : 32'd0;
    assign top_13_10_write_en =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign top_13_11_clk =
     1'b1 ? clk : 1'd0;
    assign top_13_11_in =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? top_12_11_out : 32'd0;
    assign top_13_11_write_en =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? 1'd1 : 1'd0;
    assign top_13_12_clk =
     1'b1 ? clk : 1'd0;
    assign top_13_12_in =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? top_12_12_out : 32'd0;
    assign top_13_12_write_en =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? 1'd1 : 1'd0;
    assign top_13_13_clk =
     1'b1 ? clk : 1'd0;
    assign top_13_13_in =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? top_12_13_out : 32'd0;
    assign top_13_13_write_en =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? 1'd1 : 1'd0;
    assign top_13_14_clk =
     1'b1 ? clk : 1'd0;
    assign top_13_14_in =
     fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go ? top_12_14_out : 32'd0;
    assign top_13_14_write_en =
     fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go ? 1'd1 : 1'd0;
    assign top_13_15_clk =
     1'b1 ? clk : 1'd0;
    assign top_13_15_in =
     fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go ? top_12_15_out : 32'd0;
    assign top_13_15_write_en =
     fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go ? 1'd1 : 1'd0;
    assign top_13_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_13_2_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? top_12_2_out : 32'd0;
    assign top_13_2_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign top_13_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_13_3_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? top_12_3_out : 32'd0;
    assign top_13_3_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign top_13_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_13_4_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? top_12_4_out : 32'd0;
    assign top_13_4_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign top_13_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_13_5_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? top_12_5_out : 32'd0;
    assign top_13_5_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign top_13_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_13_6_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? top_12_6_out : 32'd0;
    assign top_13_6_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign top_13_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_13_7_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? top_12_7_out : 32'd0;
    assign top_13_7_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign top_13_8_clk =
     1'b1 ? clk : 1'd0;
    assign top_13_8_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? top_12_8_out : 32'd0;
    assign top_13_8_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign top_13_9_clk =
     1'b1 ? clk : 1'd0;
    assign top_13_9_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? top_12_9_out : 32'd0;
    assign top_13_9_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign top_14_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_14_0_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? top_13_0_out : 32'd0;
    assign top_14_0_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign top_14_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_14_1_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? top_13_1_out : 32'd0;
    assign top_14_1_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign top_14_10_clk =
     1'b1 ? clk : 1'd0;
    assign top_14_10_in =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? top_13_10_out : 32'd0;
    assign top_14_10_write_en =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? 1'd1 : 1'd0;
    assign top_14_11_clk =
     1'b1 ? clk : 1'd0;
    assign top_14_11_in =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? top_13_11_out : 32'd0;
    assign top_14_11_write_en =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? 1'd1 : 1'd0;
    assign top_14_12_clk =
     1'b1 ? clk : 1'd0;
    assign top_14_12_in =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? top_13_12_out : 32'd0;
    assign top_14_12_write_en =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? 1'd1 : 1'd0;
    assign top_14_13_clk =
     1'b1 ? clk : 1'd0;
    assign top_14_13_in =
     fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go ? top_13_13_out : 32'd0;
    assign top_14_13_write_en =
     fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go ? 1'd1 : 1'd0;
    assign top_14_14_clk =
     1'b1 ? clk : 1'd0;
    assign top_14_14_in =
     fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go ? top_13_14_out : 32'd0;
    assign top_14_14_write_en =
     fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go ? 1'd1 : 1'd0;
    assign top_14_15_clk =
     1'b1 ? clk : 1'd0;
    assign top_14_15_in =
     fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go | fsm89_out < 1'd1 & fsm92_out == 10'd266 & go ? top_13_15_out : 32'd0;
    assign top_14_15_write_en =
     fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go | fsm89_out < 1'd1 & fsm92_out == 10'd266 & go ? 1'd1 : 1'd0;
    assign top_14_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_14_2_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? top_13_2_out : 32'd0;
    assign top_14_2_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign top_14_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_14_3_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? top_13_3_out : 32'd0;
    assign top_14_3_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign top_14_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_14_4_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? top_13_4_out : 32'd0;
    assign top_14_4_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign top_14_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_14_5_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? top_13_5_out : 32'd0;
    assign top_14_5_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign top_14_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_14_6_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? top_13_6_out : 32'd0;
    assign top_14_6_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign top_14_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_14_7_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? top_13_7_out : 32'd0;
    assign top_14_7_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign top_14_8_clk =
     1'b1 ? clk : 1'd0;
    assign top_14_8_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? top_13_8_out : 32'd0;
    assign top_14_8_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign top_14_9_clk =
     1'b1 ? clk : 1'd0;
    assign top_14_9_in =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? top_13_9_out : 32'd0;
    assign top_14_9_write_en =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign top_15_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_15_0_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? top_14_0_out : 32'd0;
    assign top_15_0_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign top_15_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_15_1_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? top_14_1_out : 32'd0;
    assign top_15_1_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign top_15_10_clk =
     1'b1 ? clk : 1'd0;
    assign top_15_10_in =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? top_14_10_out : 32'd0;
    assign top_15_10_write_en =
     fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go ? 1'd1 : 1'd0;
    assign top_15_11_clk =
     1'b1 ? clk : 1'd0;
    assign top_15_11_in =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? top_14_11_out : 32'd0;
    assign top_15_11_write_en =
     fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go ? 1'd1 : 1'd0;
    assign top_15_12_clk =
     1'b1 ? clk : 1'd0;
    assign top_15_12_in =
     fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go ? top_14_12_out : 32'd0;
    assign top_15_12_write_en =
     fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go ? 1'd1 : 1'd0;
    assign top_15_13_clk =
     1'b1 ? clk : 1'd0;
    assign top_15_13_in =
     fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go ? top_14_13_out : 32'd0;
    assign top_15_13_write_en =
     fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go ? 1'd1 : 1'd0;
    assign top_15_14_clk =
     1'b1 ? clk : 1'd0;
    assign top_15_14_in =
     fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go | fsm89_out < 1'd1 & fsm92_out == 10'd266 & go ? top_14_14_out : 32'd0;
    assign top_15_14_write_en =
     fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go | fsm89_out < 1'd1 & fsm92_out == 10'd266 & go ? 1'd1 : 1'd0;
    assign top_15_15_clk =
     1'b1 ? clk : 1'd0;
    assign top_15_15_in =
     fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go | fsm89_out < 1'd1 & fsm92_out == 10'd266 & go | fsm91_out < 1'd1 & fsm92_out == 10'd272 & go ? top_14_15_out : 32'd0;
    assign top_15_15_write_en =
     fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go | fsm81_out < 1'd1 & fsm92_out == 10'd242 & go | fsm83_out < 1'd1 & fsm92_out == 10'd248 & go | fsm85_out < 1'd1 & fsm92_out == 10'd254 & go | fsm87_out < 1'd1 & fsm92_out == 10'd260 & go | fsm89_out < 1'd1 & fsm92_out == 10'd266 & go | fsm91_out < 1'd1 & fsm92_out == 10'd272 & go ? 1'd1 : 1'd0;
    assign top_15_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_15_2_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? top_14_2_out : 32'd0;
    assign top_15_2_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign top_15_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_15_3_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? top_14_3_out : 32'd0;
    assign top_15_3_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign top_15_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_15_4_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? top_14_4_out : 32'd0;
    assign top_15_4_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign top_15_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_15_5_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? top_14_5_out : 32'd0;
    assign top_15_5_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign top_15_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_15_6_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? top_14_6_out : 32'd0;
    assign top_15_6_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign top_15_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_15_7_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? top_14_7_out : 32'd0;
    assign top_15_7_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign top_15_8_clk =
     1'b1 ? clk : 1'd0;
    assign top_15_8_in =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? top_14_8_out : 32'd0;
    assign top_15_8_write_en =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign top_15_9_clk =
     1'b1 ? clk : 1'd0;
    assign top_15_9_in =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? top_14_9_out : 32'd0;
    assign top_15_9_write_en =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? 1'd1 : 1'd0;
    assign top_1_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_0_in =
     fsm3_out < 1'd1 & fsm92_out == 10'd8 & go | fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go ? top_0_0_out : 32'd0;
    assign top_1_0_write_en =
     fsm3_out < 1'd1 & fsm92_out == 10'd8 & go | fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go ? 1'd1 : 1'd0;
    assign top_1_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_1_in =
     fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go ? top_0_1_out : 32'd0;
    assign top_1_1_write_en =
     fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go ? 1'd1 : 1'd0;
    assign top_1_10_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_10_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? top_0_10_out : 32'd0;
    assign top_1_10_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign top_1_11_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_11_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? top_0_11_out : 32'd0;
    assign top_1_11_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign top_1_12_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_12_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? top_0_12_out : 32'd0;
    assign top_1_12_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign top_1_13_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_13_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? top_0_13_out : 32'd0;
    assign top_1_13_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign top_1_14_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_14_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? top_0_14_out : 32'd0;
    assign top_1_14_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign top_1_15_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_15_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? top_0_15_out : 32'd0;
    assign top_1_15_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign top_1_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_2_in =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? top_0_2_out : 32'd0;
    assign top_1_2_write_en =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? 1'd1 : 1'd0;
    assign top_1_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_3_in =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? top_0_3_out : 32'd0;
    assign top_1_3_write_en =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? 1'd1 : 1'd0;
    assign top_1_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_4_in =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? top_0_4_out : 32'd0;
    assign top_1_4_write_en =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? 1'd1 : 1'd0;
    assign top_1_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_5_in =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? top_0_5_out : 32'd0;
    assign top_1_5_write_en =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? 1'd1 : 1'd0;
    assign top_1_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_6_in =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? top_0_6_out : 32'd0;
    assign top_1_6_write_en =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign top_1_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_7_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? top_0_7_out : 32'd0;
    assign top_1_7_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign top_1_8_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_8_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? top_0_8_out : 32'd0;
    assign top_1_8_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign top_1_9_clk =
     1'b1 ? clk : 1'd0;
    assign top_1_9_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? top_0_9_out : 32'd0;
    assign top_1_9_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign top_2_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_0_in =
     fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go ? top_1_0_out : 32'd0;
    assign top_2_0_write_en =
     fsm5_out < 1'd1 & fsm92_out == 10'd14 & go | fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go ? 1'd1 : 1'd0;
    assign top_2_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_1_in =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? top_1_1_out : 32'd0;
    assign top_2_1_write_en =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? 1'd1 : 1'd0;
    assign top_2_10_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_10_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? top_1_10_out : 32'd0;
    assign top_2_10_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign top_2_11_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_11_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? top_1_11_out : 32'd0;
    assign top_2_11_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign top_2_12_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_12_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? top_1_12_out : 32'd0;
    assign top_2_12_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign top_2_13_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_13_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? top_1_13_out : 32'd0;
    assign top_2_13_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign top_2_14_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_14_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? top_1_14_out : 32'd0;
    assign top_2_14_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign top_2_15_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_15_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? top_1_15_out : 32'd0;
    assign top_2_15_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign top_2_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_2_in =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? top_1_2_out : 32'd0;
    assign top_2_2_write_en =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? 1'd1 : 1'd0;
    assign top_2_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_3_in =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? top_1_3_out : 32'd0;
    assign top_2_3_write_en =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? 1'd1 : 1'd0;
    assign top_2_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_4_in =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? top_1_4_out : 32'd0;
    assign top_2_4_write_en =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? 1'd1 : 1'd0;
    assign top_2_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_5_in =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? top_1_5_out : 32'd0;
    assign top_2_5_write_en =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign top_2_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_6_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? top_1_6_out : 32'd0;
    assign top_2_6_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign top_2_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_7_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? top_1_7_out : 32'd0;
    assign top_2_7_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign top_2_8_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_8_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? top_1_8_out : 32'd0;
    assign top_2_8_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign top_2_9_clk =
     1'b1 ? clk : 1'd0;
    assign top_2_9_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? top_1_9_out : 32'd0;
    assign top_2_9_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign top_3_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_0_in =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? top_2_0_out : 32'd0;
    assign top_3_0_write_en =
     fsm7_out < 1'd1 & fsm92_out == 10'd20 & go | fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go ? 1'd1 : 1'd0;
    assign top_3_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_1_in =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? top_2_1_out : 32'd0;
    assign top_3_1_write_en =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? 1'd1 : 1'd0;
    assign top_3_10_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_10_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? top_2_10_out : 32'd0;
    assign top_3_10_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign top_3_11_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_11_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? top_2_11_out : 32'd0;
    assign top_3_11_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign top_3_12_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_12_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? top_2_12_out : 32'd0;
    assign top_3_12_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign top_3_13_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_13_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? top_2_13_out : 32'd0;
    assign top_3_13_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign top_3_14_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_14_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? top_2_14_out : 32'd0;
    assign top_3_14_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign top_3_15_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_15_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? top_2_15_out : 32'd0;
    assign top_3_15_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign top_3_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_2_in =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? top_2_2_out : 32'd0;
    assign top_3_2_write_en =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? 1'd1 : 1'd0;
    assign top_3_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_3_in =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? top_2_3_out : 32'd0;
    assign top_3_3_write_en =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? 1'd1 : 1'd0;
    assign top_3_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_4_in =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? top_2_4_out : 32'd0;
    assign top_3_4_write_en =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign top_3_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_5_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? top_2_5_out : 32'd0;
    assign top_3_5_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign top_3_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_6_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? top_2_6_out : 32'd0;
    assign top_3_6_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign top_3_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_7_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? top_2_7_out : 32'd0;
    assign top_3_7_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign top_3_8_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_8_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? top_2_8_out : 32'd0;
    assign top_3_8_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign top_3_9_clk =
     1'b1 ? clk : 1'd0;
    assign top_3_9_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? top_2_9_out : 32'd0;
    assign top_3_9_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign top_4_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_0_in =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? top_3_0_out : 32'd0;
    assign top_4_0_write_en =
     fsm9_out < 1'd1 & fsm92_out == 10'd26 & go | fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go ? 1'd1 : 1'd0;
    assign top_4_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_1_in =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? top_3_1_out : 32'd0;
    assign top_4_1_write_en =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? 1'd1 : 1'd0;
    assign top_4_10_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_10_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? top_3_10_out : 32'd0;
    assign top_4_10_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign top_4_11_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_11_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? top_3_11_out : 32'd0;
    assign top_4_11_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign top_4_12_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_12_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? top_3_12_out : 32'd0;
    assign top_4_12_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign top_4_13_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_13_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? top_3_13_out : 32'd0;
    assign top_4_13_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign top_4_14_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_14_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? top_3_14_out : 32'd0;
    assign top_4_14_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign top_4_15_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_15_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? top_3_15_out : 32'd0;
    assign top_4_15_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign top_4_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_2_in =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? top_3_2_out : 32'd0;
    assign top_4_2_write_en =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? 1'd1 : 1'd0;
    assign top_4_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_3_in =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? top_3_3_out : 32'd0;
    assign top_4_3_write_en =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign top_4_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_4_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? top_3_4_out : 32'd0;
    assign top_4_4_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign top_4_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_5_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? top_3_5_out : 32'd0;
    assign top_4_5_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign top_4_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_6_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? top_3_6_out : 32'd0;
    assign top_4_6_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign top_4_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_7_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? top_3_7_out : 32'd0;
    assign top_4_7_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign top_4_8_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_8_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? top_3_8_out : 32'd0;
    assign top_4_8_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign top_4_9_clk =
     1'b1 ? clk : 1'd0;
    assign top_4_9_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? top_3_9_out : 32'd0;
    assign top_4_9_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign top_5_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_0_in =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? top_4_0_out : 32'd0;
    assign top_5_0_write_en =
     fsm11_out < 1'd1 & fsm92_out == 10'd32 & go | fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go ? 1'd1 : 1'd0;
    assign top_5_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_1_in =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? top_4_1_out : 32'd0;
    assign top_5_1_write_en =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? 1'd1 : 1'd0;
    assign top_5_10_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_10_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? top_4_10_out : 32'd0;
    assign top_5_10_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign top_5_11_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_11_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? top_4_11_out : 32'd0;
    assign top_5_11_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign top_5_12_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_12_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? top_4_12_out : 32'd0;
    assign top_5_12_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign top_5_13_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_13_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? top_4_13_out : 32'd0;
    assign top_5_13_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign top_5_14_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_14_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? top_4_14_out : 32'd0;
    assign top_5_14_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign top_5_15_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_15_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? top_4_15_out : 32'd0;
    assign top_5_15_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign top_5_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_2_in =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? top_4_2_out : 32'd0;
    assign top_5_2_write_en =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign top_5_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_3_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? top_4_3_out : 32'd0;
    assign top_5_3_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign top_5_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_4_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? top_4_4_out : 32'd0;
    assign top_5_4_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign top_5_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_5_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? top_4_5_out : 32'd0;
    assign top_5_5_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign top_5_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_6_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? top_4_6_out : 32'd0;
    assign top_5_6_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign top_5_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_7_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? top_4_7_out : 32'd0;
    assign top_5_7_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign top_5_8_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_8_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? top_4_8_out : 32'd0;
    assign top_5_8_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign top_5_9_clk =
     1'b1 ? clk : 1'd0;
    assign top_5_9_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? top_4_9_out : 32'd0;
    assign top_5_9_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign top_6_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_0_in =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? top_5_0_out : 32'd0;
    assign top_6_0_write_en =
     fsm13_out < 1'd1 & fsm92_out == 10'd38 & go | fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go ? 1'd1 : 1'd0;
    assign top_6_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_1_in =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? top_5_1_out : 32'd0;
    assign top_6_1_write_en =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign top_6_10_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_10_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? top_5_10_out : 32'd0;
    assign top_6_10_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign top_6_11_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_11_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? top_5_11_out : 32'd0;
    assign top_6_11_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign top_6_12_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_12_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? top_5_12_out : 32'd0;
    assign top_6_12_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign top_6_13_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_13_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? top_5_13_out : 32'd0;
    assign top_6_13_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign top_6_14_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_14_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? top_5_14_out : 32'd0;
    assign top_6_14_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign top_6_15_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_15_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? top_5_15_out : 32'd0;
    assign top_6_15_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign top_6_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_2_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? top_5_2_out : 32'd0;
    assign top_6_2_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign top_6_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_3_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? top_5_3_out : 32'd0;
    assign top_6_3_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign top_6_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_4_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? top_5_4_out : 32'd0;
    assign top_6_4_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign top_6_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_5_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? top_5_5_out : 32'd0;
    assign top_6_5_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign top_6_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_6_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? top_5_6_out : 32'd0;
    assign top_6_6_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign top_6_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_7_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? top_5_7_out : 32'd0;
    assign top_6_7_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign top_6_8_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_8_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? top_5_8_out : 32'd0;
    assign top_6_8_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign top_6_9_clk =
     1'b1 ? clk : 1'd0;
    assign top_6_9_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? top_5_9_out : 32'd0;
    assign top_6_9_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign top_7_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_0_in =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? top_6_0_out : 32'd0;
    assign top_7_0_write_en =
     fsm15_out < 1'd1 & fsm92_out == 10'd44 & go | fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go ? 1'd1 : 1'd0;
    assign top_7_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_1_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? top_6_1_out : 32'd0;
    assign top_7_1_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign top_7_10_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_10_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? top_6_10_out : 32'd0;
    assign top_7_10_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign top_7_11_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_11_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? top_6_11_out : 32'd0;
    assign top_7_11_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign top_7_12_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_12_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? top_6_12_out : 32'd0;
    assign top_7_12_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign top_7_13_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_13_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? top_6_13_out : 32'd0;
    assign top_7_13_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign top_7_14_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_14_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? top_6_14_out : 32'd0;
    assign top_7_14_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign top_7_15_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_15_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? top_6_15_out : 32'd0;
    assign top_7_15_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign top_7_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_2_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? top_6_2_out : 32'd0;
    assign top_7_2_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign top_7_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_3_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? top_6_3_out : 32'd0;
    assign top_7_3_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign top_7_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_4_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? top_6_4_out : 32'd0;
    assign top_7_4_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign top_7_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_5_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? top_6_5_out : 32'd0;
    assign top_7_5_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign top_7_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_6_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? top_6_6_out : 32'd0;
    assign top_7_6_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign top_7_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_7_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? top_6_7_out : 32'd0;
    assign top_7_7_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign top_7_8_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_8_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? top_6_8_out : 32'd0;
    assign top_7_8_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign top_7_9_clk =
     1'b1 ? clk : 1'd0;
    assign top_7_9_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? top_6_9_out : 32'd0;
    assign top_7_9_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign top_8_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_8_0_in =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? top_7_0_out : 32'd0;
    assign top_8_0_write_en =
     fsm17_out < 1'd1 & fsm92_out == 10'd50 & go | fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go ? 1'd1 : 1'd0;
    assign top_8_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_8_1_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? top_7_1_out : 32'd0;
    assign top_8_1_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign top_8_10_clk =
     1'b1 ? clk : 1'd0;
    assign top_8_10_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? top_7_10_out : 32'd0;
    assign top_8_10_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
    assign top_8_11_clk =
     1'b1 ? clk : 1'd0;
    assign top_8_11_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? top_7_11_out : 32'd0;
    assign top_8_11_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign top_8_12_clk =
     1'b1 ? clk : 1'd0;
    assign top_8_12_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? top_7_12_out : 32'd0;
    assign top_8_12_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign top_8_13_clk =
     1'b1 ? clk : 1'd0;
    assign top_8_13_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? top_7_13_out : 32'd0;
    assign top_8_13_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign top_8_14_clk =
     1'b1 ? clk : 1'd0;
    assign top_8_14_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? top_7_14_out : 32'd0;
    assign top_8_14_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign top_8_15_clk =
     1'b1 ? clk : 1'd0;
    assign top_8_15_in =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? top_7_15_out : 32'd0;
    assign top_8_15_write_en =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign top_8_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_8_2_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? top_7_2_out : 32'd0;
    assign top_8_2_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign top_8_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_8_3_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? top_7_3_out : 32'd0;
    assign top_8_3_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign top_8_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_8_4_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? top_7_4_out : 32'd0;
    assign top_8_4_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign top_8_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_8_5_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? top_7_5_out : 32'd0;
    assign top_8_5_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign top_8_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_8_6_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? top_7_6_out : 32'd0;
    assign top_8_6_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign top_8_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_8_7_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? top_7_7_out : 32'd0;
    assign top_8_7_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign top_8_8_clk =
     1'b1 ? clk : 1'd0;
    assign top_8_8_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? top_7_8_out : 32'd0;
    assign top_8_8_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign top_8_9_clk =
     1'b1 ? clk : 1'd0;
    assign top_8_9_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? top_7_9_out : 32'd0;
    assign top_8_9_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign top_9_0_clk =
     1'b1 ? clk : 1'd0;
    assign top_9_0_in =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? top_8_0_out : 32'd0;
    assign top_9_0_write_en =
     fsm19_out < 1'd1 & fsm92_out == 10'd56 & go | fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go ? 1'd1 : 1'd0;
    assign top_9_1_clk =
     1'b1 ? clk : 1'd0;
    assign top_9_1_in =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? top_8_1_out : 32'd0;
    assign top_9_1_write_en =
     fsm21_out < 1'd1 & fsm92_out == 10'd62 & go | fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go ? 1'd1 : 1'd0;
    assign top_9_10_clk =
     1'b1 ? clk : 1'd0;
    assign top_9_10_in =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? top_8_10_out : 32'd0;
    assign top_9_10_write_en =
     fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go ? 1'd1 : 1'd0;
    assign top_9_11_clk =
     1'b1 ? clk : 1'd0;
    assign top_9_11_in =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? top_8_11_out : 32'd0;
    assign top_9_11_write_en =
     fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go ? 1'd1 : 1'd0;
    assign top_9_12_clk =
     1'b1 ? clk : 1'd0;
    assign top_9_12_in =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? top_8_12_out : 32'd0;
    assign top_9_12_write_en =
     fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go ? 1'd1 : 1'd0;
    assign top_9_13_clk =
     1'b1 ? clk : 1'd0;
    assign top_9_13_in =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? top_8_13_out : 32'd0;
    assign top_9_13_write_en =
     fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go ? 1'd1 : 1'd0;
    assign top_9_14_clk =
     1'b1 ? clk : 1'd0;
    assign top_9_14_in =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? top_8_14_out : 32'd0;
    assign top_9_14_write_en =
     fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go ? 1'd1 : 1'd0;
    assign top_9_15_clk =
     1'b1 ? clk : 1'd0;
    assign top_9_15_in =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? top_8_15_out : 32'd0;
    assign top_9_15_write_en =
     fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go | fsm69_out < 1'd1 & fsm92_out == 10'd206 & go | fsm71_out < 1'd1 & fsm92_out == 10'd212 & go | fsm73_out < 1'd1 & fsm92_out == 10'd218 & go | fsm75_out < 1'd1 & fsm92_out == 10'd224 & go | fsm77_out < 1'd1 & fsm92_out == 10'd230 & go | fsm79_out < 1'd1 & fsm92_out == 10'd236 & go ? 1'd1 : 1'd0;
    assign top_9_2_clk =
     1'b1 ? clk : 1'd0;
    assign top_9_2_in =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? top_8_2_out : 32'd0;
    assign top_9_2_write_en =
     fsm23_out < 1'd1 & fsm92_out == 10'd68 & go | fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go ? 1'd1 : 1'd0;
    assign top_9_3_clk =
     1'b1 ? clk : 1'd0;
    assign top_9_3_in =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? top_8_3_out : 32'd0;
    assign top_9_3_write_en =
     fsm25_out < 1'd1 & fsm92_out == 10'd74 & go | fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go ? 1'd1 : 1'd0;
    assign top_9_4_clk =
     1'b1 ? clk : 1'd0;
    assign top_9_4_in =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? top_8_4_out : 32'd0;
    assign top_9_4_write_en =
     fsm27_out < 1'd1 & fsm92_out == 10'd80 & go | fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go ? 1'd1 : 1'd0;
    assign top_9_5_clk =
     1'b1 ? clk : 1'd0;
    assign top_9_5_in =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? top_8_5_out : 32'd0;
    assign top_9_5_write_en =
     fsm29_out < 1'd1 & fsm92_out == 10'd86 & go | fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go ? 1'd1 : 1'd0;
    assign top_9_6_clk =
     1'b1 ? clk : 1'd0;
    assign top_9_6_in =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? top_8_6_out : 32'd0;
    assign top_9_6_write_en =
     fsm31_out < 1'd1 & fsm92_out == 10'd92 & go | fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go ? 1'd1 : 1'd0;
    assign top_9_7_clk =
     1'b1 ? clk : 1'd0;
    assign top_9_7_in =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? top_8_7_out : 32'd0;
    assign top_9_7_write_en =
     fsm33_out < 1'd1 & fsm92_out == 10'd98 & go | fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go ? 1'd1 : 1'd0;
    assign top_9_8_clk =
     1'b1 ? clk : 1'd0;
    assign top_9_8_in =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? top_8_8_out : 32'd0;
    assign top_9_8_write_en =
     fsm35_out < 1'd1 & fsm92_out == 10'd104 & go | fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go ? 1'd1 : 1'd0;
    assign top_9_9_clk =
     1'b1 ? clk : 1'd0;
    assign top_9_9_in =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? top_8_9_out : 32'd0;
    assign top_9_9_write_en =
     fsm37_out < 1'd1 & fsm92_out == 10'd110 & go | fsm39_out < 1'd1 & fsm92_out == 10'd116 & go | fsm41_out < 1'd1 & fsm92_out == 10'd122 & go | fsm43_out < 1'd1 & fsm92_out == 10'd128 & go | fsm45_out < 1'd1 & fsm92_out == 10'd134 & go | fsm47_out < 1'd1 & fsm92_out == 10'd140 & go | fsm49_out < 1'd1 & fsm92_out == 10'd146 & go | fsm51_out < 1'd1 & fsm92_out == 10'd152 & go | fsm53_out < 1'd1 & fsm92_out == 10'd158 & go | fsm55_out < 1'd1 & fsm92_out == 10'd164 & go | fsm57_out < 1'd1 & fsm92_out == 10'd170 & go | fsm59_out < 1'd1 & fsm92_out == 10'd176 & go | fsm61_out < 1'd1 & fsm92_out == 10'd182 & go | fsm63_out < 1'd1 & fsm92_out == 10'd188 & go | fsm65_out < 1'd1 & fsm92_out == 10'd194 & go | fsm67_out < 1'd1 & fsm92_out == 10'd200 & go ? 1'd1 : 1'd0;
endmodule

module mac_pe (
    input logic [31:0] top,
    input logic [31:0] left,
    output logic [31:0] out,
    input logic go,
    input logic clk,
    output logic done
);
    logic [31:0] acc_in;
    logic acc_write_en;
    logic acc_clk;
    logic [31:0] acc_out;
    logic acc_done;
    logic [31:0] mul_reg_in;
    logic mul_reg_write_en;
    logic mul_reg_clk;
    logic [31:0] mul_reg_out;
    logic mul_reg_done;
    logic [31:0] add_left;
    logic [31:0] add_right;
    logic [31:0] add_out;
    logic mul_clk;
    logic mul_go;
    logic [31:0] mul_left;
    logic [31:0] mul_right;
    logic [31:0] mul_out;
    logic mul_done;
    logic [2:0] fsm_in;
    logic fsm_write_en;
    logic fsm_clk;
    logic [2:0] fsm_out;
    logic fsm_done;
    logic [2:0] incr_left;
    logic [2:0] incr_right;
    logic [2:0] incr_out;
    initial begin
        acc_in = 32'd0;
        acc_write_en = 1'd0;
        acc_clk = 1'd0;
        mul_reg_in = 32'd0;
        mul_reg_write_en = 1'd0;
        mul_reg_clk = 1'd0;
        add_left = 32'd0;
        add_right = 32'd0;
        mul_clk = 1'd0;
        mul_go = 1'd0;
        mul_left = 32'd0;
        mul_right = 32'd0;
        fsm_in = 3'd0;
        fsm_write_en = 1'd0;
        fsm_clk = 1'd0;
        incr_left = 3'd0;
        incr_right = 3'd0;
    end
    std_reg # (
        .width(32)
    ) acc (
        .clk(acc_clk),
        .done(acc_done),
        .in(acc_in),
        .out(acc_out),
        .write_en(acc_write_en)
    );
    std_reg # (
        .width(32)
    ) mul_reg (
        .clk(mul_reg_clk),
        .done(mul_reg_done),
        .in(mul_reg_in),
        .out(mul_reg_out),
        .write_en(mul_reg_write_en)
    );
    std_add # (
        .width(32)
    ) add (
        .left(add_left),
        .out(add_out),
        .right(add_right)
    );
    std_mult_pipe # (
        .width(32)
    ) mul (
        .clk(mul_clk),
        .done(mul_done),
        .go(mul_go),
        .left(mul_left),
        .out(mul_out),
        .right(mul_right)
    );
    std_reg # (
        .width(3)
    ) fsm (
        .clk(fsm_clk),
        .done(fsm_done),
        .in(fsm_in),
        .out(fsm_out),
        .write_en(fsm_write_en)
    );
    std_add # (
        .width(3)
    ) incr (
        .left(incr_left),
        .out(incr_out),
        .right(incr_right)
    );
    assign done =
     fsm_out == 3'd5 ? 1'd1 : 1'd0;
    assign out =
     1'b1 ? acc_out : 32'd0;
    assign acc_clk =
     1'b1 ? clk : 1'd0;
    assign acc_in =
     fsm_out == 3'd4 & go ? add_out : 32'd0;
    assign acc_write_en =
     fsm_out == 3'd4 & go ? 1'd1 : 1'd0;
    assign add_left =
     fsm_out == 3'd4 & go ? acc_out : 32'd0;
    assign add_right =
     fsm_out == 3'd4 & go ? mul_reg_out : 32'd0;
    assign fsm_clk =
     1'b1 ? clk : 1'd0;
    assign fsm_in =
     fsm_out == 3'd5 ? 3'd0 :
     fsm_out != 3'd5 & go ? incr_out : 3'd0;
    assign fsm_write_en =
     fsm_out != 3'd5 & go | fsm_out == 3'd5 ? 1'd1 : 1'd0;
    assign incr_left =
     go ? 3'd1 : 3'd0;
    assign incr_right =
     go ? fsm_out : 3'd0;
    assign mul_clk =
     1'b1 ? clk : 1'd0;
    assign mul_go =
     ~mul_done & fsm_out < 3'd4 & go ? 1'd1 : 1'd0;
    assign mul_left =
     fsm_out < 3'd4 & go ? top : 32'd0;
    assign mul_right =
     fsm_out < 3'd4 & go ? left : 32'd0;
    assign mul_reg_clk =
     1'b1 ? clk : 1'd0;
    assign mul_reg_in =
     mul_done & fsm_out < 3'd4 & go ? mul_out : 32'd0;
    assign mul_reg_write_en =
     mul_done & fsm_out < 3'd4 & go ? 1'd1 : 1'd0;
endmodule
