
/// This is mostly used for testing the static guarantees currently.
/// A realistic implementation would probably take four cycles.
module pipelined_mult (
    input wire clk,
    input wire reset,
    // inputs
    input wire [31:0] left,
    input wire [31:0] right,
    // The input has been committed
    output wire [31:0] out
);

logic [31:0] lt, rt, buff0, buff1, buff2, tmp_prod;

assign out = buff2;
assign tmp_prod = lt * rt;

always_ff @(posedge clk) begin
    if (reset) begin
        lt <= 0;
        rt <= 0;
        buff0 <= 0;
        buff1 <= 0;
        buff2 <= 0;
    end else begin
        lt <= left;
        rt <= right;
        buff0 <= tmp_prod;
        buff1 <= buff0;
        buff2 <= buff1;
    end
end

endmodule

module bb_pipelined_mult(
	               input wire [31:0] left,
	               input wire [31:0] right,
	               output wire [31:0] out,
	               input wire clk
	               );
`ifdef __ICARUS__
   reg [31:0] reg0;
   reg [31:0] reg1;
   reg [31:0] reg2;
   reg [31:0] reg3;
   always @( posedge clk ) begin
      reg0 <= left * right;
      reg1 <= reg0;
      reg2 <= reg1;
      reg3 <= reg2;
   end
   assign out = reg3;
`elsif VERILATOR
   reg [31:0] reg0;
   reg [31:0] reg1;
   reg [31:0] reg2;
   reg [31:0] reg3;
   always @( posedge clk ) begin
      reg0 <= left * right;
      reg1 <= reg0;
      reg2 <= reg1;
      reg3 <= reg2;
   end
   assign out = reg3;
`else
   // mul_uint32 is a black box module generated by Xilinx's IP Core generator.
   // Generation commands are in the synth.tcl file.
   mul_uint32 mul_uint32 (
                   .A(left),
                   .B(right),
                   .P(out),
                   .CLK(clk)
                   );
`endif
endmodule
/* verilator lint_off MULTITOP */
/// =================== Unsigned, Fixed Point =========================
module std_fp_add #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  assign out = left + right;
endmodule

module std_fp_sub #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module std_fp_mult_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16,
    parameter SIGNED = 0
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    input  logic             go,
    input  logic             clk,
    input  logic             reset,
    output logic [WIDTH-1:0] out,
    output logic             done
);
  logic [WIDTH-1:0]          rtmp;
  logic [WIDTH-1:0]          ltmp;
  logic [(WIDTH << 1) - 1:0] out_tmp;
  // Buffer used to walk through the 3 cycles of the pipeline.
  logic done_buf[1:0];

  assign done = done_buf[1];

  assign out = out_tmp[(WIDTH << 1) - INT_WIDTH - 1 : WIDTH - INT_WIDTH];

  // If the done buffer is completely empty and go is high then execution
  // just started.
  logic start;
  assign start = go;

  // Start sending the done signal.
  always_ff @(posedge clk) begin
    if (start)
      done_buf[0] <= 1;
    else
      done_buf[0] <= 0;
  end

  // Push the done signal through the pipeline.
  always_ff @(posedge clk) begin
    if (go) begin
      done_buf[1] <= done_buf[0];
    end else begin
      done_buf[1] <= 0;
    end
  end

  // Register the inputs
  always_ff @(posedge clk) begin
    if (reset) begin
      rtmp <= 0;
      ltmp <= 0;
    end else if (go) begin
      if (SIGNED) begin
        rtmp <= $signed(right);
        ltmp <= $signed(left);
      end else begin
        rtmp <= right;
        ltmp <= left;
      end
    end else begin
      rtmp <= 0;
      ltmp <= 0;
    end

  end

  // Compute the output and save it into out_tmp
  always_ff @(posedge clk) begin
    if (reset) begin
      out_tmp <= 0;
    end else if (go) begin
      if (SIGNED) begin
        // In the first cycle, this performs an invalid computation because
        // ltmp and rtmp only get their actual values in cycle 1
        out_tmp <= $signed(
          { {WIDTH{ltmp[WIDTH-1]}}, ltmp} *
          { {WIDTH{rtmp[WIDTH-1]}}, rtmp}
        );
      end else begin
        out_tmp <= ltmp * rtmp;
      end
    end else begin
      out_tmp <= out_tmp;
    end
  end
endmodule

/* verilator lint_off WIDTH */
module std_fp_div_pipe #(
  parameter WIDTH = 32,
  parameter INT_WIDTH = 16,
  parameter FRAC_WIDTH = 16
) (
    input  logic             go,
    input  logic             clk,
    input  logic             reset,
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out_remainder,
    output logic [WIDTH-1:0] out_quotient,
    output logic             done
);
    localparam ITERATIONS = WIDTH + FRAC_WIDTH;

    logic [WIDTH-1:0] quotient, quotient_next;
    logic [WIDTH:0] acc, acc_next;
    logic [$clog2(ITERATIONS)-1:0] idx;
    logic start, running, finished, dividend_is_zero;

    assign start = go && !running;
    assign dividend_is_zero = start && left == 0;
    assign finished = idx == ITERATIONS - 1 && running;

    always_ff @(posedge clk) begin
      if (reset || finished || dividend_is_zero)
        running <= 0;
      else if (start)
        running <= 1;
      else
        running <= running;
    end

    always_comb begin
      if (acc >= {1'b0, right}) begin
        acc_next = acc - right;
        {acc_next, quotient_next} = {acc_next[WIDTH-1:0], quotient, 1'b1};
      end else begin
        {acc_next, quotient_next} = {acc, quotient} << 1;
      end
    end

    // `done` signaling
    always_ff @(posedge clk) begin
      if (dividend_is_zero || finished)
        done <= 1;
      else
        done <= 0;
    end

    always_ff @(posedge clk) begin
      if (running)
        idx <= idx + 1;
      else
        idx <= 0;
    end

    always_ff @(posedge clk) begin
      if (reset) begin
        out_quotient <= 0;
        out_remainder <= 0;
      end else if (start) begin
        out_quotient <= 0;
        out_remainder <= left;
      end else if (go == 0) begin
        out_quotient <= out_quotient;
        out_remainder <= out_remainder;
      end else if (dividend_is_zero) begin
        out_quotient <= 0;
        out_remainder <= 0;
      end else if (finished) begin
        out_quotient <= quotient_next;
        out_remainder <= out_remainder;
      end else begin
        out_quotient <= out_quotient;
        if (right <= out_remainder)
          out_remainder <= out_remainder - right;
        else
          out_remainder <= out_remainder;
      end
    end

    always_ff @(posedge clk) begin
      if (reset) begin
        acc <= 0;
        quotient <= 0;
      end else if (start) begin
        {acc, quotient} <= {{WIDTH{1'b0}}, left, 1'b0};
      end else begin
        acc <= acc_next;
        quotient <= quotient_next;
      end
    end
endmodule

module std_fp_gt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic             out
);
  assign out = left > right;
endmodule

/// =================== Signed, Fixed Point =========================
module std_fp_sadd #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left + right);
endmodule

module std_fp_ssub #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);

  assign out = $signed(left - right);
endmodule

module std_fp_smult_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  [WIDTH-1:0]              left,
    input  [WIDTH-1:0]              right,
    input  logic                    reset,
    input  logic                    go,
    input  logic                    clk,
    output logic [WIDTH-1:0]        out,
    output logic                    done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(INT_WIDTH),
    .FRAC_WIDTH(FRAC_WIDTH),
    .SIGNED(1)
  ) comp (
    .clk(clk),
    .done(done),
    .reset(reset),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

module std_fp_sdiv_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input                     clk,
    input                     go,
    input                     reset,
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out_quotient,
    output signed [WIDTH-1:0] out_remainder,
    output logic              done
);

  logic signed [WIDTH-1:0] left_abs, right_abs, comp_out_q, comp_out_r, right_save, out_rem_intermediate;

  // Registers to figure out how to transform outputs.
  logic different_signs, left_sign, right_sign;

  // Latch the value of control registers so that their available after
  // go signal becomes low.
  always_ff @(posedge clk) begin
    if (go) begin
      right_save <= right_abs;
      left_sign <= left[WIDTH-1];
      right_sign <= right[WIDTH-1];
    end else begin
      left_sign <= left_sign;
      right_save <= right_save;
      right_sign <= right_sign;
    end
  end

  assign right_abs = right[WIDTH-1] ? -right : right;
  assign left_abs = left[WIDTH-1] ? -left : left;

  assign different_signs = left_sign ^ right_sign;
  assign out_quotient = different_signs ? -comp_out_q : comp_out_q;

  // Remainder is computed as:
  //  t0 = |left| % |right|
  //  t1 = if left * right < 0 and t0 != 0 then |right| - t0 else t0
  //  rem = if right < 0 then -t1 else t1
  assign out_rem_intermediate = different_signs & |comp_out_r ? $signed(right_save - comp_out_r) : comp_out_r;
  assign out_remainder = right_sign ? -out_rem_intermediate : out_rem_intermediate;

  std_fp_div_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(INT_WIDTH),
    .FRAC_WIDTH(FRAC_WIDTH)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left_abs),
    .right(right_abs),
    .out_quotient(comp_out_q),
    .out_remainder(comp_out_r)
  );
endmodule

module std_fp_sgt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic signed [WIDTH-1:0] left,
    input  logic signed [WIDTH-1:0] right,
    output logic signed             out
);
  assign out = $signed(left > right);
endmodule

module std_fp_slt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
   input logic signed [WIDTH-1:0] left,
   input logic signed [WIDTH-1:0] right,
   output logic signed            out
);
  assign out = $signed(left < right);
endmodule

/// =================== Unsigned, Bitnum =========================
module std_mult_pipe #(
    parameter WIDTH = 32
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    input  logic             reset,
    input  logic             go,
    input  logic             clk,
    output logic [WIDTH-1:0] out,
    output logic             done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(WIDTH),
    .FRAC_WIDTH(0),
    .SIGNED(0)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

module std_div_pipe #(
    parameter WIDTH = 32
) (
    input                    reset,
    input                    clk,
    input                    go,
    input        [WIDTH-1:0] left,
    input        [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out_remainder,
    output logic [WIDTH-1:0] out_quotient,
    output logic             done
);

  logic [WIDTH-1:0] dividend;
  logic [(WIDTH-1)*2:0] divisor;
  logic [WIDTH-1:0] quotient;
  logic [WIDTH-1:0] quotient_msk;
  logic start, running, finished, dividend_is_zero;

  assign start = go && !running;
  assign finished = quotient_msk == 0 && running;
  assign dividend_is_zero = start && left == 0;

  always_ff @(posedge clk) begin
    // Early return if the divisor is zero.
    if (finished || dividend_is_zero)
      done <= 1;
    else
      done <= 0;
  end

  always_ff @(posedge clk) begin
    if (reset || finished || dividend_is_zero)
      running <= 0;
    else if (start)
      running <= 1;
    else
      running <= running;
  end

  // Outputs
  always_ff @(posedge clk) begin
    if (dividend_is_zero || start) begin
      out_quotient <= 0;
      out_remainder <= 0;
    end else if (finished) begin
      out_quotient <= quotient;
      out_remainder <= dividend;
    end else begin
      // Otherwise, explicitly latch the values.
      out_quotient <= out_quotient;
      out_remainder <= out_remainder;
    end
  end

  // Calculate the quotient mask.
  always_ff @(posedge clk) begin
    if (start)
      quotient_msk <= 1 << WIDTH - 1;
    else if (running)
      quotient_msk <= quotient_msk >> 1;
    else
      quotient_msk <= quotient_msk;
  end

  // Calculate the quotient.
  always_ff @(posedge clk) begin
    if (start)
      quotient <= 0;
    else if (divisor <= dividend)
      quotient <= quotient | quotient_msk;
    else
      quotient <= quotient;
  end

  // Calculate the dividend.
  always_ff @(posedge clk) begin
    if (start)
      dividend <= left;
    else if (divisor <= dividend)
      dividend <= dividend - divisor;
    else
      dividend <= dividend;
  end

  always_ff @(posedge clk) begin
    if (start) begin
      divisor <= right << WIDTH - 1;
    end else if (finished) begin
      divisor <= 0;
    end else begin
      divisor <= divisor >> 1;
    end
  end

  // Simulation self test against unsynthesizable implementation.
  `ifdef VERILATOR
    logic [WIDTH-1:0] l, r;
    always_ff @(posedge clk) begin
      if (go) begin
        l <= left;
        r <= right;
      end else begin
        l <= l;
        r <= r;
      end
    end

    always @(posedge clk) begin
      if (done && $unsigned(out_remainder) != $unsigned(l % r))
        $error(
          "\nstd_div_pipe (Remainder): Computed and golden outputs do not match!\n",
          "left: %0d", $unsigned(l),
          "  right: %0d\n", $unsigned(r),
          "expected: %0d", $unsigned(l % r),
          "  computed: %0d", $unsigned(out_remainder)
        );

      if (done && $unsigned(out_quotient) != $unsigned(l / r))
        $error(
          "\nstd_div_pipe (Quotient): Computed and golden outputs do not match!\n",
          "left: %0d", $unsigned(l),
          "  right: %0d\n", $unsigned(r),
          "expected: %0d", $unsigned(l / r),
          "  computed: %0d", $unsigned(out_quotient)
        );
    end
  `endif
endmodule

/// =================== Signed, Bitnum =========================
module std_sadd #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left + right);
endmodule

module std_ssub #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left - right);
endmodule

module std_smult_pipe #(
    parameter WIDTH = 32
) (
    input  logic                    reset,
    input  logic                    go,
    input  logic                    clk,
    input  signed       [WIDTH-1:0] left,
    input  signed       [WIDTH-1:0] right,
    output logic signed [WIDTH-1:0] out,
    output logic                    done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(WIDTH),
    .FRAC_WIDTH(0),
    .SIGNED(1)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

/* verilator lint_off WIDTH */
module std_sdiv_pipe #(
    parameter WIDTH = 32
) (
    input                           reset,
    input                           clk,
    input                           go,
    input  logic signed [WIDTH-1:0] left,
    input  logic signed [WIDTH-1:0] right,
    output logic signed [WIDTH-1:0] out_quotient,
    output logic signed [WIDTH-1:0] out_remainder,
    output logic                    done
);

  logic signed [WIDTH-1:0] left_abs, right_abs, comp_out_q, comp_out_r, right_save, out_rem_intermediate;

  // Registers to figure out how to transform outputs.
  logic different_signs, left_sign, right_sign;

  // Latch the value of control registers so that their available after
  // go signal becomes low.
  always_ff @(posedge clk) begin
    if (go) begin
      right_save <= right_abs;
      left_sign <= left[WIDTH-1];
      right_sign <= right[WIDTH-1];
    end else begin
      left_sign <= left_sign;
      right_save <= right_save;
      right_sign <= right_sign;
    end
  end

  assign right_abs = right[WIDTH-1] ? -right : right;
  assign left_abs = left[WIDTH-1] ? -left : left;

  assign different_signs = left_sign ^ right_sign;
  assign out_quotient = different_signs ? -comp_out_q : comp_out_q;

  // Remainder is computed as:
  //  t0 = |left| % |right|
  //  t1 = if left * right < 0 and t0 != 0 then |right| - t0 else t0
  //  rem = if right < 0 then -t1 else t1
  assign out_rem_intermediate = different_signs & |comp_out_r ? $signed(right_save - comp_out_r) : comp_out_r;
  assign out_remainder = right_sign ? -out_rem_intermediate : out_rem_intermediate;

  std_div_pipe #(
    .WIDTH(WIDTH)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left_abs),
    .right(right_abs),
    .out_quotient(comp_out_q),
    .out_remainder(comp_out_r)
  );

  // Simulation self test against unsynthesizable implementation.
  `ifdef VERILATOR
    logic signed [WIDTH-1:0] l, r;
    always_ff @(posedge clk) begin
      if (go) begin
        l <= left;
        r <= right;
      end else begin
        l <= l;
        r <= r;
      end
    end

    always @(posedge clk) begin
      if (done && out_quotient != $signed(l / r))
        $error(
          "\nstd_sdiv_pipe (Quotient): Computed and golden outputs do not match!\n",
          "left: %0d", l,
          "  right: %0d\n", r,
          "expected: %0d", $signed(l / r),
          "  computed: %0d", $signed(out_quotient),
        );
      if (done && out_remainder != $signed(((l % r) + r) % r))
        $error(
          "\nstd_sdiv_pipe (Remainder): Computed and golden outputs do not match!\n",
          "left: %0d", l,
          "  right: %0d\n", r,
          "expected: %0d", $signed(((l % r) + r) % r),
          "  computed: %0d", $signed(out_remainder),
        );
    end
  `endif
endmodule

module std_sgt #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left > right);
endmodule

module std_slt #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left < right);
endmodule

module std_seq #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left == right);
endmodule

module std_sneq #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left != right);
endmodule

module std_sge #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left >= right);
endmodule

module std_sle #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left <= right);
endmodule

module std_slsh #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = left <<< right;
endmodule

module std_srsh #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = left >>> right;
endmodule

/**
 * Core primitives for Calyx.
 * Implements core primitives used by the compiler.
 *
 * Conventions:
 * - All parameter names must be SNAKE_CASE and all caps.
 * - Port names must be snake_case, no caps.
 */
`default_nettype none

module std_slice #(
    parameter IN_WIDTH  = 32,
    parameter OUT_WIDTH = 32
) (
   input wire                   logic [ IN_WIDTH-1:0] in,
   output logic [OUT_WIDTH-1:0] out
);
  assign out = in[OUT_WIDTH-1:0];

  `ifdef VERILATOR
    always_comb begin
      if (IN_WIDTH < OUT_WIDTH)
        $error(
          "std_slice: Input width less than output width\n",
          "IN_WIDTH: %0d", IN_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_pad #(
    parameter IN_WIDTH  = 32,
    parameter OUT_WIDTH = 32
) (
   input wire logic [IN_WIDTH-1:0]  in,
   output logic     [OUT_WIDTH-1:0] out
);
  localparam EXTEND = OUT_WIDTH - IN_WIDTH;
  assign out = { {EXTEND {1'b0}}, in};

  `ifdef VERILATOR
    always_comb begin
      if (IN_WIDTH > OUT_WIDTH)
        $error(
          "std_pad: Output width less than input width\n",
          "IN_WIDTH: %0d", IN_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_cat #(
  parameter LEFT_WIDTH  = 32,
  parameter RIGHT_WIDTH = 32,
  parameter OUT_WIDTH = 64
) (
  input wire logic [LEFT_WIDTH-1:0] left,
  input wire logic [RIGHT_WIDTH-1:0] right,
  output logic [OUT_WIDTH-1:0] out
);
  assign out = {left, right};

  `ifdef VERILATOR
    always_comb begin
      if (LEFT_WIDTH + RIGHT_WIDTH != OUT_WIDTH)
        $error(
          "std_cat: Output width must equal sum of input widths\n",
          "LEFT_WIDTH: %0d", LEFT_WIDTH,
          "RIGHT_WIDTH: %0d", RIGHT_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_not #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] in,
   output logic [WIDTH-1:0] out
);
  assign out = ~in;
endmodule

module std_and #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left & right;
endmodule

module std_or #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left | right;
endmodule

module std_xor #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left ^ right;
endmodule

module std_sub #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module std_gt #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left > right;
endmodule

module std_lt #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left < right;
endmodule

module std_eq #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left == right;
endmodule

module std_neq #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left != right;
endmodule

module std_ge #(
    parameter WIDTH = 32
) (
    input wire   logic [WIDTH-1:0] left,
    input wire   logic [WIDTH-1:0] right,
    output logic out
);
  assign out = left >= right;
endmodule

module std_le #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left <= right;
endmodule

module std_lsh #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left << right;
endmodule

module std_rsh #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left >> right;
endmodule

/// this primitive is intended to be used
/// for lowering purposes (not in source programs)
module std_mux #(
    parameter WIDTH = 32
) (
   input wire               logic cond,
   input wire               logic [WIDTH-1:0] tru,
   input wire               logic [WIDTH-1:0] fal,
   output logic [WIDTH-1:0] out
);
  assign out = cond ? tru : fal;
endmodule

module std_mem_d1 #(
    parameter WIDTH = 32,
    parameter SIZE = 16,
    parameter IDX_SIZE = 4
) (
   input wire                logic [IDX_SIZE-1:0] addr0,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  logic [WIDTH-1:0] mem[SIZE-1:0];

  /* verilator lint_off WIDTH */
  assign read_data = mem[addr0];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= SIZE)
        $error(
          "std_mem_d1: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "SIZE: %0d", SIZE
        );
    end
  `endif
endmodule

module std_mem_d2 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0];

  assign read_data = mem[addr0][addr1];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d2: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d2: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
    end
  `endif
endmodule

module std_mem_d3 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D2_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4,
    parameter D2_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [D2_IDX_SIZE-1:0] addr2,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0][D2_SIZE-1:0];

  assign read_data = mem[addr0][addr1][addr2];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1][addr2] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
      if (addr2 >= D2_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr2: %0d\n", addr2,
          "D2_SIZE: %0d", D2_SIZE
        );
    end
  `endif
endmodule

module std_mem_d4 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D2_SIZE = 16,
    parameter D3_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4,
    parameter D2_IDX_SIZE = 4,
    parameter D3_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [D2_IDX_SIZE-1:0] addr2,
   input wire                logic [D3_IDX_SIZE-1:0] addr3,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0][D2_SIZE-1:0][D3_SIZE-1:0];

  assign read_data = mem[addr0][addr1][addr2][addr3];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1][addr2][addr3] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
      if (addr2 >= D2_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr2: %0d\n", addr2,
          "D2_SIZE: %0d", D2_SIZE
        );
      if (addr3 >= D3_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr3: %0d\n", addr3,
          "D3_SIZE: %0d", D3_SIZE
        );
    end
  `endif
endmodule

`default_nettype wire

module undef #(
    parameter WIDTH = 32
) (
   output logic [WIDTH-1:0] out
);
assign out = 'x;
endmodule

module std_const #(
    parameter WIDTH = 32,
    parameter VALUE = 32
) (
   output logic [WIDTH-1:0] out
);
assign out = VALUE;
endmodule

module std_wire #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] in,
   output logic [WIDTH-1:0] out
);
assign out = in;
endmodule

module std_add #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] left,
   input logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
assign out = left + right;
endmodule

module std_reg #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] in,
   input logic write_en,
   input logic clk,
   input logic reset,
   output logic [WIDTH-1:0] out,
   output logic done
);
always_ff @(posedge clk) begin
    if (reset) begin
       out <= 0;
       done <= 0;
    end else if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module mac_pe(
  input logic [31:0] top,
  input logic [31:0] left,
  input logic mul_ready,
  output logic [31:0] out,
  input logic go,
  input logic clk,
  input logic reset,
  output logic done
);
// COMPONENT START: mac_pe
logic [31:0] acc_in;
logic acc_write_en;
logic acc_clk;
logic acc_reset;
logic [31:0] acc_out;
logic acc_done;
logic [31:0] add_left;
logic [31:0] add_right;
logic [31:0] add_out;
logic mul_clk;
logic [31:0] mul_left;
logic [31:0] mul_right;
logic [31:0] mul_out;
logic fsm_in;
logic fsm_write_en;
logic fsm_clk;
logic fsm_reset;
logic fsm_out;
logic fsm_done;
logic ud_out;
logic adder_left;
logic adder_right;
logic adder_out;
logic signal_reg_in;
logic signal_reg_write_en;
logic signal_reg_clk;
logic signal_reg_reset;
logic signal_reg_out;
logic signal_reg_done;
logic early_reset_static_par_go_in;
logic early_reset_static_par_go_out;
logic early_reset_static_par_done_in;
logic early_reset_static_par_done_out;
logic wrapper_early_reset_static_par_go_in;
logic wrapper_early_reset_static_par_go_out;
logic wrapper_early_reset_static_par_done_in;
logic wrapper_early_reset_static_par_done_out;
std_reg # (
    .WIDTH(32)
) acc (
    .clk(acc_clk),
    .done(acc_done),
    .in(acc_in),
    .out(acc_out),
    .reset(acc_reset),
    .write_en(acc_write_en)
);
std_add # (
    .WIDTH(32)
) add (
    .left(add_left),
    .out(add_out),
    .right(add_right)
);
bb_pipelined_mult mul (
    .clk(mul_clk),
    .left(mul_left),
    .out(mul_out),
    .right(mul_right)
);
std_reg # (
    .WIDTH(1)
) fsm (
    .clk(fsm_clk),
    .done(fsm_done),
    .in(fsm_in),
    .out(fsm_out),
    .reset(fsm_reset),
    .write_en(fsm_write_en)
);
undef # (
    .WIDTH(1)
) ud (
    .out(ud_out)
);
std_add # (
    .WIDTH(1)
) adder (
    .left(adder_left),
    .out(adder_out),
    .right(adder_right)
);
std_reg # (
    .WIDTH(1)
) signal_reg (
    .clk(signal_reg_clk),
    .done(signal_reg_done),
    .in(signal_reg_in),
    .out(signal_reg_out),
    .reset(signal_reg_reset),
    .write_en(signal_reg_write_en)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_go (
    .in(early_reset_static_par_go_in),
    .out(early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_done (
    .in(early_reset_static_par_done_in),
    .out(early_reset_static_par_done_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_go (
    .in(wrapper_early_reset_static_par_go_in),
    .out(wrapper_early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_done (
    .in(wrapper_early_reset_static_par_done_in),
    .out(wrapper_early_reset_static_par_done_out)
);
wire _guard0 = 1;
wire _guard1 = early_reset_static_par_go_out;
wire _guard2 = early_reset_static_par_go_out;
wire _guard3 = wrapper_early_reset_static_par_done_out;
wire _guard4 = early_reset_static_par_go_out;
wire _guard5 = fsm_out != 1'd0;
wire _guard6 = early_reset_static_par_go_out;
wire _guard7 = _guard5 & _guard6;
wire _guard8 = fsm_out == 1'd0;
wire _guard9 = early_reset_static_par_go_out;
wire _guard10 = _guard8 & _guard9;
wire _guard11 = early_reset_static_par_go_out;
wire _guard12 = early_reset_static_par_go_out;
wire _guard13 = fsm_out == 1'd0;
wire _guard14 = signal_reg_out;
wire _guard15 = _guard13 & _guard14;
wire _guard16 = fsm_out == 1'd0;
wire _guard17 = signal_reg_out;
wire _guard18 = _guard16 & _guard17;
wire _guard19 = fsm_out == 1'd0;
wire _guard20 = signal_reg_out;
wire _guard21 = ~_guard20;
wire _guard22 = _guard19 & _guard21;
wire _guard23 = wrapper_early_reset_static_par_go_out;
wire _guard24 = _guard22 & _guard23;
wire _guard25 = _guard18 | _guard24;
wire _guard26 = fsm_out == 1'd0;
wire _guard27 = signal_reg_out;
wire _guard28 = ~_guard27;
wire _guard29 = _guard26 & _guard28;
wire _guard30 = wrapper_early_reset_static_par_go_out;
wire _guard31 = _guard29 & _guard30;
wire _guard32 = fsm_out == 1'd0;
wire _guard33 = signal_reg_out;
wire _guard34 = _guard32 & _guard33;
wire _guard35 = early_reset_static_par_go_out;
wire _guard36 = early_reset_static_par_go_out;
wire _guard37 = early_reset_static_par_go_out;
wire _guard38 = early_reset_static_par_go_out;
wire _guard39 = wrapper_early_reset_static_par_go_out;
assign acc_write_en =
  _guard1 ? mul_ready :
  1'd0;
assign acc_clk = clk;
assign acc_reset = reset;
assign acc_in = add_out;
assign done = _guard3;
assign out = acc_out;
assign fsm_write_en = _guard4;
assign fsm_clk = clk;
assign fsm_reset = reset;
assign fsm_in =
  _guard7 ? adder_out :
  _guard10 ? 1'd0 :
  1'd0;
assign adder_left =
  _guard11 ? fsm_out :
  1'd0;
assign adder_right = _guard12;
assign wrapper_early_reset_static_par_go_in = go;
assign wrapper_early_reset_static_par_done_in = _guard15;
assign early_reset_static_par_done_in = ud_out;
assign signal_reg_write_en = _guard25;
assign signal_reg_clk = clk;
assign signal_reg_reset = reset;
assign signal_reg_in =
  _guard31 ? 1'd1 :
  _guard34 ? 1'd0 :
  1'd0;
assign add_left = acc_out;
assign add_right = mul_out;
assign mul_clk = clk;
assign mul_left =
  _guard37 ? top :
  32'd0;
assign mul_right =
  _guard38 ? left :
  32'd0;
assign early_reset_static_par_go_in = _guard39;
// COMPONENT END: mac_pe
endmodule
module main(
  input logic go,
  input logic clk,
  input logic reset,
  output logic done,
  output logic [4:0] t0_addr0,
  output logic [31:0] t0_write_data,
  output logic t0_write_en,
  output logic t0_clk,
  output logic t0_reset,
  input logic [31:0] t0_read_data,
  input logic t0_done,
  output logic [4:0] t1_addr0,
  output logic [31:0] t1_write_data,
  output logic t1_write_en,
  output logic t1_clk,
  output logic t1_reset,
  input logic [31:0] t1_read_data,
  input logic t1_done,
  output logic [4:0] t2_addr0,
  output logic [31:0] t2_write_data,
  output logic t2_write_en,
  output logic t2_clk,
  output logic t2_reset,
  input logic [31:0] t2_read_data,
  input logic t2_done,
  output logic [4:0] t3_addr0,
  output logic [31:0] t3_write_data,
  output logic t3_write_en,
  output logic t3_clk,
  output logic t3_reset,
  input logic [31:0] t3_read_data,
  input logic t3_done,
  output logic [4:0] t4_addr0,
  output logic [31:0] t4_write_data,
  output logic t4_write_en,
  output logic t4_clk,
  output logic t4_reset,
  input logic [31:0] t4_read_data,
  input logic t4_done,
  output logic [4:0] t5_addr0,
  output logic [31:0] t5_write_data,
  output logic t5_write_en,
  output logic t5_clk,
  output logic t5_reset,
  input logic [31:0] t5_read_data,
  input logic t5_done,
  output logic [4:0] t6_addr0,
  output logic [31:0] t6_write_data,
  output logic t6_write_en,
  output logic t6_clk,
  output logic t6_reset,
  input logic [31:0] t6_read_data,
  input logic t6_done,
  output logic [4:0] t7_addr0,
  output logic [31:0] t7_write_data,
  output logic t7_write_en,
  output logic t7_clk,
  output logic t7_reset,
  input logic [31:0] t7_read_data,
  input logic t7_done,
  output logic [4:0] t8_addr0,
  output logic [31:0] t8_write_data,
  output logic t8_write_en,
  output logic t8_clk,
  output logic t8_reset,
  input logic [31:0] t8_read_data,
  input logic t8_done,
  output logic [4:0] t9_addr0,
  output logic [31:0] t9_write_data,
  output logic t9_write_en,
  output logic t9_clk,
  output logic t9_reset,
  input logic [31:0] t9_read_data,
  input logic t9_done,
  output logic [4:0] t10_addr0,
  output logic [31:0] t10_write_data,
  output logic t10_write_en,
  output logic t10_clk,
  output logic t10_reset,
  input logic [31:0] t10_read_data,
  input logic t10_done,
  output logic [4:0] t11_addr0,
  output logic [31:0] t11_write_data,
  output logic t11_write_en,
  output logic t11_clk,
  output logic t11_reset,
  input logic [31:0] t11_read_data,
  input logic t11_done,
  output logic [4:0] t12_addr0,
  output logic [31:0] t12_write_data,
  output logic t12_write_en,
  output logic t12_clk,
  output logic t12_reset,
  input logic [31:0] t12_read_data,
  input logic t12_done,
  output logic [4:0] t13_addr0,
  output logic [31:0] t13_write_data,
  output logic t13_write_en,
  output logic t13_clk,
  output logic t13_reset,
  input logic [31:0] t13_read_data,
  input logic t13_done,
  output logic [4:0] t14_addr0,
  output logic [31:0] t14_write_data,
  output logic t14_write_en,
  output logic t14_clk,
  output logic t14_reset,
  input logic [31:0] t14_read_data,
  input logic t14_done,
  output logic [4:0] t15_addr0,
  output logic [31:0] t15_write_data,
  output logic t15_write_en,
  output logic t15_clk,
  output logic t15_reset,
  input logic [31:0] t15_read_data,
  input logic t15_done,
  output logic [4:0] l0_addr0,
  output logic [31:0] l0_write_data,
  output logic l0_write_en,
  output logic l0_clk,
  output logic l0_reset,
  input logic [31:0] l0_read_data,
  input logic l0_done,
  output logic [4:0] l1_addr0,
  output logic [31:0] l1_write_data,
  output logic l1_write_en,
  output logic l1_clk,
  output logic l1_reset,
  input logic [31:0] l1_read_data,
  input logic l1_done,
  output logic [4:0] l2_addr0,
  output logic [31:0] l2_write_data,
  output logic l2_write_en,
  output logic l2_clk,
  output logic l2_reset,
  input logic [31:0] l2_read_data,
  input logic l2_done,
  output logic [4:0] l3_addr0,
  output logic [31:0] l3_write_data,
  output logic l3_write_en,
  output logic l3_clk,
  output logic l3_reset,
  input logic [31:0] l3_read_data,
  input logic l3_done,
  output logic [4:0] l4_addr0,
  output logic [31:0] l4_write_data,
  output logic l4_write_en,
  output logic l4_clk,
  output logic l4_reset,
  input logic [31:0] l4_read_data,
  input logic l4_done,
  output logic [4:0] l5_addr0,
  output logic [31:0] l5_write_data,
  output logic l5_write_en,
  output logic l5_clk,
  output logic l5_reset,
  input logic [31:0] l5_read_data,
  input logic l5_done,
  output logic [4:0] l6_addr0,
  output logic [31:0] l6_write_data,
  output logic l6_write_en,
  output logic l6_clk,
  output logic l6_reset,
  input logic [31:0] l6_read_data,
  input logic l6_done,
  output logic [4:0] l7_addr0,
  output logic [31:0] l7_write_data,
  output logic l7_write_en,
  output logic l7_clk,
  output logic l7_reset,
  input logic [31:0] l7_read_data,
  input logic l7_done,
  output logic [4:0] l8_addr0,
  output logic [31:0] l8_write_data,
  output logic l8_write_en,
  output logic l8_clk,
  output logic l8_reset,
  input logic [31:0] l8_read_data,
  input logic l8_done,
  output logic [4:0] l9_addr0,
  output logic [31:0] l9_write_data,
  output logic l9_write_en,
  output logic l9_clk,
  output logic l9_reset,
  input logic [31:0] l9_read_data,
  input logic l9_done,
  output logic [4:0] l10_addr0,
  output logic [31:0] l10_write_data,
  output logic l10_write_en,
  output logic l10_clk,
  output logic l10_reset,
  input logic [31:0] l10_read_data,
  input logic l10_done,
  output logic [4:0] l11_addr0,
  output logic [31:0] l11_write_data,
  output logic l11_write_en,
  output logic l11_clk,
  output logic l11_reset,
  input logic [31:0] l11_read_data,
  input logic l11_done,
  output logic [4:0] l12_addr0,
  output logic [31:0] l12_write_data,
  output logic l12_write_en,
  output logic l12_clk,
  output logic l12_reset,
  input logic [31:0] l12_read_data,
  input logic l12_done,
  output logic [4:0] l13_addr0,
  output logic [31:0] l13_write_data,
  output logic l13_write_en,
  output logic l13_clk,
  output logic l13_reset,
  input logic [31:0] l13_read_data,
  input logic l13_done,
  output logic [4:0] l14_addr0,
  output logic [31:0] l14_write_data,
  output logic l14_write_en,
  output logic l14_clk,
  output logic l14_reset,
  input logic [31:0] l14_read_data,
  input logic l14_done,
  output logic [4:0] l15_addr0,
  output logic [31:0] l15_write_data,
  output logic l15_write_en,
  output logic l15_clk,
  output logic l15_reset,
  input logic [31:0] l15_read_data,
  input logic l15_done,
  output logic [4:0] out_mem_0_addr0,
  output logic [31:0] out_mem_0_write_data,
  output logic out_mem_0_write_en,
  output logic out_mem_0_clk,
  output logic out_mem_0_reset,
  input logic [31:0] out_mem_0_read_data,
  input logic out_mem_0_done,
  output logic [4:0] out_mem_1_addr0,
  output logic [31:0] out_mem_1_write_data,
  output logic out_mem_1_write_en,
  output logic out_mem_1_clk,
  output logic out_mem_1_reset,
  input logic [31:0] out_mem_1_read_data,
  input logic out_mem_1_done,
  output logic [4:0] out_mem_2_addr0,
  output logic [31:0] out_mem_2_write_data,
  output logic out_mem_2_write_en,
  output logic out_mem_2_clk,
  output logic out_mem_2_reset,
  input logic [31:0] out_mem_2_read_data,
  input logic out_mem_2_done,
  output logic [4:0] out_mem_3_addr0,
  output logic [31:0] out_mem_3_write_data,
  output logic out_mem_3_write_en,
  output logic out_mem_3_clk,
  output logic out_mem_3_reset,
  input logic [31:0] out_mem_3_read_data,
  input logic out_mem_3_done,
  output logic [4:0] out_mem_4_addr0,
  output logic [31:0] out_mem_4_write_data,
  output logic out_mem_4_write_en,
  output logic out_mem_4_clk,
  output logic out_mem_4_reset,
  input logic [31:0] out_mem_4_read_data,
  input logic out_mem_4_done,
  output logic [4:0] out_mem_5_addr0,
  output logic [31:0] out_mem_5_write_data,
  output logic out_mem_5_write_en,
  output logic out_mem_5_clk,
  output logic out_mem_5_reset,
  input logic [31:0] out_mem_5_read_data,
  input logic out_mem_5_done,
  output logic [4:0] out_mem_6_addr0,
  output logic [31:0] out_mem_6_write_data,
  output logic out_mem_6_write_en,
  output logic out_mem_6_clk,
  output logic out_mem_6_reset,
  input logic [31:0] out_mem_6_read_data,
  input logic out_mem_6_done,
  output logic [4:0] out_mem_7_addr0,
  output logic [31:0] out_mem_7_write_data,
  output logic out_mem_7_write_en,
  output logic out_mem_7_clk,
  output logic out_mem_7_reset,
  input logic [31:0] out_mem_7_read_data,
  input logic out_mem_7_done,
  output logic [4:0] out_mem_8_addr0,
  output logic [31:0] out_mem_8_write_data,
  output logic out_mem_8_write_en,
  output logic out_mem_8_clk,
  output logic out_mem_8_reset,
  input logic [31:0] out_mem_8_read_data,
  input logic out_mem_8_done,
  output logic [4:0] out_mem_9_addr0,
  output logic [31:0] out_mem_9_write_data,
  output logic out_mem_9_write_en,
  output logic out_mem_9_clk,
  output logic out_mem_9_reset,
  input logic [31:0] out_mem_9_read_data,
  input logic out_mem_9_done,
  output logic [4:0] out_mem_10_addr0,
  output logic [31:0] out_mem_10_write_data,
  output logic out_mem_10_write_en,
  output logic out_mem_10_clk,
  output logic out_mem_10_reset,
  input logic [31:0] out_mem_10_read_data,
  input logic out_mem_10_done,
  output logic [4:0] out_mem_11_addr0,
  output logic [31:0] out_mem_11_write_data,
  output logic out_mem_11_write_en,
  output logic out_mem_11_clk,
  output logic out_mem_11_reset,
  input logic [31:0] out_mem_11_read_data,
  input logic out_mem_11_done,
  output logic [4:0] out_mem_12_addr0,
  output logic [31:0] out_mem_12_write_data,
  output logic out_mem_12_write_en,
  output logic out_mem_12_clk,
  output logic out_mem_12_reset,
  input logic [31:0] out_mem_12_read_data,
  input logic out_mem_12_done,
  output logic [4:0] out_mem_13_addr0,
  output logic [31:0] out_mem_13_write_data,
  output logic out_mem_13_write_en,
  output logic out_mem_13_clk,
  output logic out_mem_13_reset,
  input logic [31:0] out_mem_13_read_data,
  input logic out_mem_13_done,
  output logic [4:0] out_mem_14_addr0,
  output logic [31:0] out_mem_14_write_data,
  output logic out_mem_14_write_en,
  output logic out_mem_14_clk,
  output logic out_mem_14_reset,
  input logic [31:0] out_mem_14_read_data,
  input logic out_mem_14_done,
  output logic [4:0] out_mem_15_addr0,
  output logic [31:0] out_mem_15_write_data,
  output logic out_mem_15_write_en,
  output logic out_mem_15_clk,
  output logic out_mem_15_reset,
  input logic [31:0] out_mem_15_read_data,
  input logic out_mem_15_done
);
// COMPONENT START: main
logic [31:0] pe_0_0_top;
logic [31:0] pe_0_0_left;
logic pe_0_0_mul_ready;
logic [31:0] pe_0_0_out;
logic pe_0_0_go;
logic pe_0_0_clk;
logic pe_0_0_reset;
logic pe_0_0_done;
logic [31:0] top_0_0_in;
logic top_0_0_write_en;
logic top_0_0_clk;
logic top_0_0_reset;
logic [31:0] top_0_0_out;
logic top_0_0_done;
logic [31:0] left_0_0_in;
logic left_0_0_write_en;
logic left_0_0_clk;
logic left_0_0_reset;
logic [31:0] left_0_0_out;
logic left_0_0_done;
logic [31:0] pe_0_1_top;
logic [31:0] pe_0_1_left;
logic pe_0_1_mul_ready;
logic [31:0] pe_0_1_out;
logic pe_0_1_go;
logic pe_0_1_clk;
logic pe_0_1_reset;
logic pe_0_1_done;
logic [31:0] top_0_1_in;
logic top_0_1_write_en;
logic top_0_1_clk;
logic top_0_1_reset;
logic [31:0] top_0_1_out;
logic top_0_1_done;
logic [31:0] left_0_1_in;
logic left_0_1_write_en;
logic left_0_1_clk;
logic left_0_1_reset;
logic [31:0] left_0_1_out;
logic left_0_1_done;
logic [31:0] pe_0_2_top;
logic [31:0] pe_0_2_left;
logic pe_0_2_mul_ready;
logic [31:0] pe_0_2_out;
logic pe_0_2_go;
logic pe_0_2_clk;
logic pe_0_2_reset;
logic pe_0_2_done;
logic [31:0] top_0_2_in;
logic top_0_2_write_en;
logic top_0_2_clk;
logic top_0_2_reset;
logic [31:0] top_0_2_out;
logic top_0_2_done;
logic [31:0] left_0_2_in;
logic left_0_2_write_en;
logic left_0_2_clk;
logic left_0_2_reset;
logic [31:0] left_0_2_out;
logic left_0_2_done;
logic [31:0] pe_0_3_top;
logic [31:0] pe_0_3_left;
logic pe_0_3_mul_ready;
logic [31:0] pe_0_3_out;
logic pe_0_3_go;
logic pe_0_3_clk;
logic pe_0_3_reset;
logic pe_0_3_done;
logic [31:0] top_0_3_in;
logic top_0_3_write_en;
logic top_0_3_clk;
logic top_0_3_reset;
logic [31:0] top_0_3_out;
logic top_0_3_done;
logic [31:0] left_0_3_in;
logic left_0_3_write_en;
logic left_0_3_clk;
logic left_0_3_reset;
logic [31:0] left_0_3_out;
logic left_0_3_done;
logic [31:0] pe_0_4_top;
logic [31:0] pe_0_4_left;
logic pe_0_4_mul_ready;
logic [31:0] pe_0_4_out;
logic pe_0_4_go;
logic pe_0_4_clk;
logic pe_0_4_reset;
logic pe_0_4_done;
logic [31:0] top_0_4_in;
logic top_0_4_write_en;
logic top_0_4_clk;
logic top_0_4_reset;
logic [31:0] top_0_4_out;
logic top_0_4_done;
logic [31:0] left_0_4_in;
logic left_0_4_write_en;
logic left_0_4_clk;
logic left_0_4_reset;
logic [31:0] left_0_4_out;
logic left_0_4_done;
logic [31:0] pe_0_5_top;
logic [31:0] pe_0_5_left;
logic pe_0_5_mul_ready;
logic [31:0] pe_0_5_out;
logic pe_0_5_go;
logic pe_0_5_clk;
logic pe_0_5_reset;
logic pe_0_5_done;
logic [31:0] top_0_5_in;
logic top_0_5_write_en;
logic top_0_5_clk;
logic top_0_5_reset;
logic [31:0] top_0_5_out;
logic top_0_5_done;
logic [31:0] left_0_5_in;
logic left_0_5_write_en;
logic left_0_5_clk;
logic left_0_5_reset;
logic [31:0] left_0_5_out;
logic left_0_5_done;
logic [31:0] pe_0_6_top;
logic [31:0] pe_0_6_left;
logic pe_0_6_mul_ready;
logic [31:0] pe_0_6_out;
logic pe_0_6_go;
logic pe_0_6_clk;
logic pe_0_6_reset;
logic pe_0_6_done;
logic [31:0] top_0_6_in;
logic top_0_6_write_en;
logic top_0_6_clk;
logic top_0_6_reset;
logic [31:0] top_0_6_out;
logic top_0_6_done;
logic [31:0] left_0_6_in;
logic left_0_6_write_en;
logic left_0_6_clk;
logic left_0_6_reset;
logic [31:0] left_0_6_out;
logic left_0_6_done;
logic [31:0] pe_0_7_top;
logic [31:0] pe_0_7_left;
logic pe_0_7_mul_ready;
logic [31:0] pe_0_7_out;
logic pe_0_7_go;
logic pe_0_7_clk;
logic pe_0_7_reset;
logic pe_0_7_done;
logic [31:0] top_0_7_in;
logic top_0_7_write_en;
logic top_0_7_clk;
logic top_0_7_reset;
logic [31:0] top_0_7_out;
logic top_0_7_done;
logic [31:0] left_0_7_in;
logic left_0_7_write_en;
logic left_0_7_clk;
logic left_0_7_reset;
logic [31:0] left_0_7_out;
logic left_0_7_done;
logic [31:0] pe_0_8_top;
logic [31:0] pe_0_8_left;
logic pe_0_8_mul_ready;
logic [31:0] pe_0_8_out;
logic pe_0_8_go;
logic pe_0_8_clk;
logic pe_0_8_reset;
logic pe_0_8_done;
logic [31:0] top_0_8_in;
logic top_0_8_write_en;
logic top_0_8_clk;
logic top_0_8_reset;
logic [31:0] top_0_8_out;
logic top_0_8_done;
logic [31:0] left_0_8_in;
logic left_0_8_write_en;
logic left_0_8_clk;
logic left_0_8_reset;
logic [31:0] left_0_8_out;
logic left_0_8_done;
logic [31:0] pe_0_9_top;
logic [31:0] pe_0_9_left;
logic pe_0_9_mul_ready;
logic [31:0] pe_0_9_out;
logic pe_0_9_go;
logic pe_0_9_clk;
logic pe_0_9_reset;
logic pe_0_9_done;
logic [31:0] top_0_9_in;
logic top_0_9_write_en;
logic top_0_9_clk;
logic top_0_9_reset;
logic [31:0] top_0_9_out;
logic top_0_9_done;
logic [31:0] left_0_9_in;
logic left_0_9_write_en;
logic left_0_9_clk;
logic left_0_9_reset;
logic [31:0] left_0_9_out;
logic left_0_9_done;
logic [31:0] pe_0_10_top;
logic [31:0] pe_0_10_left;
logic pe_0_10_mul_ready;
logic [31:0] pe_0_10_out;
logic pe_0_10_go;
logic pe_0_10_clk;
logic pe_0_10_reset;
logic pe_0_10_done;
logic [31:0] top_0_10_in;
logic top_0_10_write_en;
logic top_0_10_clk;
logic top_0_10_reset;
logic [31:0] top_0_10_out;
logic top_0_10_done;
logic [31:0] left_0_10_in;
logic left_0_10_write_en;
logic left_0_10_clk;
logic left_0_10_reset;
logic [31:0] left_0_10_out;
logic left_0_10_done;
logic [31:0] pe_0_11_top;
logic [31:0] pe_0_11_left;
logic pe_0_11_mul_ready;
logic [31:0] pe_0_11_out;
logic pe_0_11_go;
logic pe_0_11_clk;
logic pe_0_11_reset;
logic pe_0_11_done;
logic [31:0] top_0_11_in;
logic top_0_11_write_en;
logic top_0_11_clk;
logic top_0_11_reset;
logic [31:0] top_0_11_out;
logic top_0_11_done;
logic [31:0] left_0_11_in;
logic left_0_11_write_en;
logic left_0_11_clk;
logic left_0_11_reset;
logic [31:0] left_0_11_out;
logic left_0_11_done;
logic [31:0] pe_0_12_top;
logic [31:0] pe_0_12_left;
logic pe_0_12_mul_ready;
logic [31:0] pe_0_12_out;
logic pe_0_12_go;
logic pe_0_12_clk;
logic pe_0_12_reset;
logic pe_0_12_done;
logic [31:0] top_0_12_in;
logic top_0_12_write_en;
logic top_0_12_clk;
logic top_0_12_reset;
logic [31:0] top_0_12_out;
logic top_0_12_done;
logic [31:0] left_0_12_in;
logic left_0_12_write_en;
logic left_0_12_clk;
logic left_0_12_reset;
logic [31:0] left_0_12_out;
logic left_0_12_done;
logic [31:0] pe_0_13_top;
logic [31:0] pe_0_13_left;
logic pe_0_13_mul_ready;
logic [31:0] pe_0_13_out;
logic pe_0_13_go;
logic pe_0_13_clk;
logic pe_0_13_reset;
logic pe_0_13_done;
logic [31:0] top_0_13_in;
logic top_0_13_write_en;
logic top_0_13_clk;
logic top_0_13_reset;
logic [31:0] top_0_13_out;
logic top_0_13_done;
logic [31:0] left_0_13_in;
logic left_0_13_write_en;
logic left_0_13_clk;
logic left_0_13_reset;
logic [31:0] left_0_13_out;
logic left_0_13_done;
logic [31:0] pe_0_14_top;
logic [31:0] pe_0_14_left;
logic pe_0_14_mul_ready;
logic [31:0] pe_0_14_out;
logic pe_0_14_go;
logic pe_0_14_clk;
logic pe_0_14_reset;
logic pe_0_14_done;
logic [31:0] top_0_14_in;
logic top_0_14_write_en;
logic top_0_14_clk;
logic top_0_14_reset;
logic [31:0] top_0_14_out;
logic top_0_14_done;
logic [31:0] left_0_14_in;
logic left_0_14_write_en;
logic left_0_14_clk;
logic left_0_14_reset;
logic [31:0] left_0_14_out;
logic left_0_14_done;
logic [31:0] pe_0_15_top;
logic [31:0] pe_0_15_left;
logic pe_0_15_mul_ready;
logic [31:0] pe_0_15_out;
logic pe_0_15_go;
logic pe_0_15_clk;
logic pe_0_15_reset;
logic pe_0_15_done;
logic [31:0] top_0_15_in;
logic top_0_15_write_en;
logic top_0_15_clk;
logic top_0_15_reset;
logic [31:0] top_0_15_out;
logic top_0_15_done;
logic [31:0] left_0_15_in;
logic left_0_15_write_en;
logic left_0_15_clk;
logic left_0_15_reset;
logic [31:0] left_0_15_out;
logic left_0_15_done;
logic [31:0] pe_1_0_top;
logic [31:0] pe_1_0_left;
logic pe_1_0_mul_ready;
logic [31:0] pe_1_0_out;
logic pe_1_0_go;
logic pe_1_0_clk;
logic pe_1_0_reset;
logic pe_1_0_done;
logic [31:0] top_1_0_in;
logic top_1_0_write_en;
logic top_1_0_clk;
logic top_1_0_reset;
logic [31:0] top_1_0_out;
logic top_1_0_done;
logic [31:0] left_1_0_in;
logic left_1_0_write_en;
logic left_1_0_clk;
logic left_1_0_reset;
logic [31:0] left_1_0_out;
logic left_1_0_done;
logic [31:0] pe_1_1_top;
logic [31:0] pe_1_1_left;
logic pe_1_1_mul_ready;
logic [31:0] pe_1_1_out;
logic pe_1_1_go;
logic pe_1_1_clk;
logic pe_1_1_reset;
logic pe_1_1_done;
logic [31:0] top_1_1_in;
logic top_1_1_write_en;
logic top_1_1_clk;
logic top_1_1_reset;
logic [31:0] top_1_1_out;
logic top_1_1_done;
logic [31:0] left_1_1_in;
logic left_1_1_write_en;
logic left_1_1_clk;
logic left_1_1_reset;
logic [31:0] left_1_1_out;
logic left_1_1_done;
logic [31:0] pe_1_2_top;
logic [31:0] pe_1_2_left;
logic pe_1_2_mul_ready;
logic [31:0] pe_1_2_out;
logic pe_1_2_go;
logic pe_1_2_clk;
logic pe_1_2_reset;
logic pe_1_2_done;
logic [31:0] top_1_2_in;
logic top_1_2_write_en;
logic top_1_2_clk;
logic top_1_2_reset;
logic [31:0] top_1_2_out;
logic top_1_2_done;
logic [31:0] left_1_2_in;
logic left_1_2_write_en;
logic left_1_2_clk;
logic left_1_2_reset;
logic [31:0] left_1_2_out;
logic left_1_2_done;
logic [31:0] pe_1_3_top;
logic [31:0] pe_1_3_left;
logic pe_1_3_mul_ready;
logic [31:0] pe_1_3_out;
logic pe_1_3_go;
logic pe_1_3_clk;
logic pe_1_3_reset;
logic pe_1_3_done;
logic [31:0] top_1_3_in;
logic top_1_3_write_en;
logic top_1_3_clk;
logic top_1_3_reset;
logic [31:0] top_1_3_out;
logic top_1_3_done;
logic [31:0] left_1_3_in;
logic left_1_3_write_en;
logic left_1_3_clk;
logic left_1_3_reset;
logic [31:0] left_1_3_out;
logic left_1_3_done;
logic [31:0] pe_1_4_top;
logic [31:0] pe_1_4_left;
logic pe_1_4_mul_ready;
logic [31:0] pe_1_4_out;
logic pe_1_4_go;
logic pe_1_4_clk;
logic pe_1_4_reset;
logic pe_1_4_done;
logic [31:0] top_1_4_in;
logic top_1_4_write_en;
logic top_1_4_clk;
logic top_1_4_reset;
logic [31:0] top_1_4_out;
logic top_1_4_done;
logic [31:0] left_1_4_in;
logic left_1_4_write_en;
logic left_1_4_clk;
logic left_1_4_reset;
logic [31:0] left_1_4_out;
logic left_1_4_done;
logic [31:0] pe_1_5_top;
logic [31:0] pe_1_5_left;
logic pe_1_5_mul_ready;
logic [31:0] pe_1_5_out;
logic pe_1_5_go;
logic pe_1_5_clk;
logic pe_1_5_reset;
logic pe_1_5_done;
logic [31:0] top_1_5_in;
logic top_1_5_write_en;
logic top_1_5_clk;
logic top_1_5_reset;
logic [31:0] top_1_5_out;
logic top_1_5_done;
logic [31:0] left_1_5_in;
logic left_1_5_write_en;
logic left_1_5_clk;
logic left_1_5_reset;
logic [31:0] left_1_5_out;
logic left_1_5_done;
logic [31:0] pe_1_6_top;
logic [31:0] pe_1_6_left;
logic pe_1_6_mul_ready;
logic [31:0] pe_1_6_out;
logic pe_1_6_go;
logic pe_1_6_clk;
logic pe_1_6_reset;
logic pe_1_6_done;
logic [31:0] top_1_6_in;
logic top_1_6_write_en;
logic top_1_6_clk;
logic top_1_6_reset;
logic [31:0] top_1_6_out;
logic top_1_6_done;
logic [31:0] left_1_6_in;
logic left_1_6_write_en;
logic left_1_6_clk;
logic left_1_6_reset;
logic [31:0] left_1_6_out;
logic left_1_6_done;
logic [31:0] pe_1_7_top;
logic [31:0] pe_1_7_left;
logic pe_1_7_mul_ready;
logic [31:0] pe_1_7_out;
logic pe_1_7_go;
logic pe_1_7_clk;
logic pe_1_7_reset;
logic pe_1_7_done;
logic [31:0] top_1_7_in;
logic top_1_7_write_en;
logic top_1_7_clk;
logic top_1_7_reset;
logic [31:0] top_1_7_out;
logic top_1_7_done;
logic [31:0] left_1_7_in;
logic left_1_7_write_en;
logic left_1_7_clk;
logic left_1_7_reset;
logic [31:0] left_1_7_out;
logic left_1_7_done;
logic [31:0] pe_1_8_top;
logic [31:0] pe_1_8_left;
logic pe_1_8_mul_ready;
logic [31:0] pe_1_8_out;
logic pe_1_8_go;
logic pe_1_8_clk;
logic pe_1_8_reset;
logic pe_1_8_done;
logic [31:0] top_1_8_in;
logic top_1_8_write_en;
logic top_1_8_clk;
logic top_1_8_reset;
logic [31:0] top_1_8_out;
logic top_1_8_done;
logic [31:0] left_1_8_in;
logic left_1_8_write_en;
logic left_1_8_clk;
logic left_1_8_reset;
logic [31:0] left_1_8_out;
logic left_1_8_done;
logic [31:0] pe_1_9_top;
logic [31:0] pe_1_9_left;
logic pe_1_9_mul_ready;
logic [31:0] pe_1_9_out;
logic pe_1_9_go;
logic pe_1_9_clk;
logic pe_1_9_reset;
logic pe_1_9_done;
logic [31:0] top_1_9_in;
logic top_1_9_write_en;
logic top_1_9_clk;
logic top_1_9_reset;
logic [31:0] top_1_9_out;
logic top_1_9_done;
logic [31:0] left_1_9_in;
logic left_1_9_write_en;
logic left_1_9_clk;
logic left_1_9_reset;
logic [31:0] left_1_9_out;
logic left_1_9_done;
logic [31:0] pe_1_10_top;
logic [31:0] pe_1_10_left;
logic pe_1_10_mul_ready;
logic [31:0] pe_1_10_out;
logic pe_1_10_go;
logic pe_1_10_clk;
logic pe_1_10_reset;
logic pe_1_10_done;
logic [31:0] top_1_10_in;
logic top_1_10_write_en;
logic top_1_10_clk;
logic top_1_10_reset;
logic [31:0] top_1_10_out;
logic top_1_10_done;
logic [31:0] left_1_10_in;
logic left_1_10_write_en;
logic left_1_10_clk;
logic left_1_10_reset;
logic [31:0] left_1_10_out;
logic left_1_10_done;
logic [31:0] pe_1_11_top;
logic [31:0] pe_1_11_left;
logic pe_1_11_mul_ready;
logic [31:0] pe_1_11_out;
logic pe_1_11_go;
logic pe_1_11_clk;
logic pe_1_11_reset;
logic pe_1_11_done;
logic [31:0] top_1_11_in;
logic top_1_11_write_en;
logic top_1_11_clk;
logic top_1_11_reset;
logic [31:0] top_1_11_out;
logic top_1_11_done;
logic [31:0] left_1_11_in;
logic left_1_11_write_en;
logic left_1_11_clk;
logic left_1_11_reset;
logic [31:0] left_1_11_out;
logic left_1_11_done;
logic [31:0] pe_1_12_top;
logic [31:0] pe_1_12_left;
logic pe_1_12_mul_ready;
logic [31:0] pe_1_12_out;
logic pe_1_12_go;
logic pe_1_12_clk;
logic pe_1_12_reset;
logic pe_1_12_done;
logic [31:0] top_1_12_in;
logic top_1_12_write_en;
logic top_1_12_clk;
logic top_1_12_reset;
logic [31:0] top_1_12_out;
logic top_1_12_done;
logic [31:0] left_1_12_in;
logic left_1_12_write_en;
logic left_1_12_clk;
logic left_1_12_reset;
logic [31:0] left_1_12_out;
logic left_1_12_done;
logic [31:0] pe_1_13_top;
logic [31:0] pe_1_13_left;
logic pe_1_13_mul_ready;
logic [31:0] pe_1_13_out;
logic pe_1_13_go;
logic pe_1_13_clk;
logic pe_1_13_reset;
logic pe_1_13_done;
logic [31:0] top_1_13_in;
logic top_1_13_write_en;
logic top_1_13_clk;
logic top_1_13_reset;
logic [31:0] top_1_13_out;
logic top_1_13_done;
logic [31:0] left_1_13_in;
logic left_1_13_write_en;
logic left_1_13_clk;
logic left_1_13_reset;
logic [31:0] left_1_13_out;
logic left_1_13_done;
logic [31:0] pe_1_14_top;
logic [31:0] pe_1_14_left;
logic pe_1_14_mul_ready;
logic [31:0] pe_1_14_out;
logic pe_1_14_go;
logic pe_1_14_clk;
logic pe_1_14_reset;
logic pe_1_14_done;
logic [31:0] top_1_14_in;
logic top_1_14_write_en;
logic top_1_14_clk;
logic top_1_14_reset;
logic [31:0] top_1_14_out;
logic top_1_14_done;
logic [31:0] left_1_14_in;
logic left_1_14_write_en;
logic left_1_14_clk;
logic left_1_14_reset;
logic [31:0] left_1_14_out;
logic left_1_14_done;
logic [31:0] pe_1_15_top;
logic [31:0] pe_1_15_left;
logic pe_1_15_mul_ready;
logic [31:0] pe_1_15_out;
logic pe_1_15_go;
logic pe_1_15_clk;
logic pe_1_15_reset;
logic pe_1_15_done;
logic [31:0] top_1_15_in;
logic top_1_15_write_en;
logic top_1_15_clk;
logic top_1_15_reset;
logic [31:0] top_1_15_out;
logic top_1_15_done;
logic [31:0] left_1_15_in;
logic left_1_15_write_en;
logic left_1_15_clk;
logic left_1_15_reset;
logic [31:0] left_1_15_out;
logic left_1_15_done;
logic [31:0] pe_2_0_top;
logic [31:0] pe_2_0_left;
logic pe_2_0_mul_ready;
logic [31:0] pe_2_0_out;
logic pe_2_0_go;
logic pe_2_0_clk;
logic pe_2_0_reset;
logic pe_2_0_done;
logic [31:0] top_2_0_in;
logic top_2_0_write_en;
logic top_2_0_clk;
logic top_2_0_reset;
logic [31:0] top_2_0_out;
logic top_2_0_done;
logic [31:0] left_2_0_in;
logic left_2_0_write_en;
logic left_2_0_clk;
logic left_2_0_reset;
logic [31:0] left_2_0_out;
logic left_2_0_done;
logic [31:0] pe_2_1_top;
logic [31:0] pe_2_1_left;
logic pe_2_1_mul_ready;
logic [31:0] pe_2_1_out;
logic pe_2_1_go;
logic pe_2_1_clk;
logic pe_2_1_reset;
logic pe_2_1_done;
logic [31:0] top_2_1_in;
logic top_2_1_write_en;
logic top_2_1_clk;
logic top_2_1_reset;
logic [31:0] top_2_1_out;
logic top_2_1_done;
logic [31:0] left_2_1_in;
logic left_2_1_write_en;
logic left_2_1_clk;
logic left_2_1_reset;
logic [31:0] left_2_1_out;
logic left_2_1_done;
logic [31:0] pe_2_2_top;
logic [31:0] pe_2_2_left;
logic pe_2_2_mul_ready;
logic [31:0] pe_2_2_out;
logic pe_2_2_go;
logic pe_2_2_clk;
logic pe_2_2_reset;
logic pe_2_2_done;
logic [31:0] top_2_2_in;
logic top_2_2_write_en;
logic top_2_2_clk;
logic top_2_2_reset;
logic [31:0] top_2_2_out;
logic top_2_2_done;
logic [31:0] left_2_2_in;
logic left_2_2_write_en;
logic left_2_2_clk;
logic left_2_2_reset;
logic [31:0] left_2_2_out;
logic left_2_2_done;
logic [31:0] pe_2_3_top;
logic [31:0] pe_2_3_left;
logic pe_2_3_mul_ready;
logic [31:0] pe_2_3_out;
logic pe_2_3_go;
logic pe_2_3_clk;
logic pe_2_3_reset;
logic pe_2_3_done;
logic [31:0] top_2_3_in;
logic top_2_3_write_en;
logic top_2_3_clk;
logic top_2_3_reset;
logic [31:0] top_2_3_out;
logic top_2_3_done;
logic [31:0] left_2_3_in;
logic left_2_3_write_en;
logic left_2_3_clk;
logic left_2_3_reset;
logic [31:0] left_2_3_out;
logic left_2_3_done;
logic [31:0] pe_2_4_top;
logic [31:0] pe_2_4_left;
logic pe_2_4_mul_ready;
logic [31:0] pe_2_4_out;
logic pe_2_4_go;
logic pe_2_4_clk;
logic pe_2_4_reset;
logic pe_2_4_done;
logic [31:0] top_2_4_in;
logic top_2_4_write_en;
logic top_2_4_clk;
logic top_2_4_reset;
logic [31:0] top_2_4_out;
logic top_2_4_done;
logic [31:0] left_2_4_in;
logic left_2_4_write_en;
logic left_2_4_clk;
logic left_2_4_reset;
logic [31:0] left_2_4_out;
logic left_2_4_done;
logic [31:0] pe_2_5_top;
logic [31:0] pe_2_5_left;
logic pe_2_5_mul_ready;
logic [31:0] pe_2_5_out;
logic pe_2_5_go;
logic pe_2_5_clk;
logic pe_2_5_reset;
logic pe_2_5_done;
logic [31:0] top_2_5_in;
logic top_2_5_write_en;
logic top_2_5_clk;
logic top_2_5_reset;
logic [31:0] top_2_5_out;
logic top_2_5_done;
logic [31:0] left_2_5_in;
logic left_2_5_write_en;
logic left_2_5_clk;
logic left_2_5_reset;
logic [31:0] left_2_5_out;
logic left_2_5_done;
logic [31:0] pe_2_6_top;
logic [31:0] pe_2_6_left;
logic pe_2_6_mul_ready;
logic [31:0] pe_2_6_out;
logic pe_2_6_go;
logic pe_2_6_clk;
logic pe_2_6_reset;
logic pe_2_6_done;
logic [31:0] top_2_6_in;
logic top_2_6_write_en;
logic top_2_6_clk;
logic top_2_6_reset;
logic [31:0] top_2_6_out;
logic top_2_6_done;
logic [31:0] left_2_6_in;
logic left_2_6_write_en;
logic left_2_6_clk;
logic left_2_6_reset;
logic [31:0] left_2_6_out;
logic left_2_6_done;
logic [31:0] pe_2_7_top;
logic [31:0] pe_2_7_left;
logic pe_2_7_mul_ready;
logic [31:0] pe_2_7_out;
logic pe_2_7_go;
logic pe_2_7_clk;
logic pe_2_7_reset;
logic pe_2_7_done;
logic [31:0] top_2_7_in;
logic top_2_7_write_en;
logic top_2_7_clk;
logic top_2_7_reset;
logic [31:0] top_2_7_out;
logic top_2_7_done;
logic [31:0] left_2_7_in;
logic left_2_7_write_en;
logic left_2_7_clk;
logic left_2_7_reset;
logic [31:0] left_2_7_out;
logic left_2_7_done;
logic [31:0] pe_2_8_top;
logic [31:0] pe_2_8_left;
logic pe_2_8_mul_ready;
logic [31:0] pe_2_8_out;
logic pe_2_8_go;
logic pe_2_8_clk;
logic pe_2_8_reset;
logic pe_2_8_done;
logic [31:0] top_2_8_in;
logic top_2_8_write_en;
logic top_2_8_clk;
logic top_2_8_reset;
logic [31:0] top_2_8_out;
logic top_2_8_done;
logic [31:0] left_2_8_in;
logic left_2_8_write_en;
logic left_2_8_clk;
logic left_2_8_reset;
logic [31:0] left_2_8_out;
logic left_2_8_done;
logic [31:0] pe_2_9_top;
logic [31:0] pe_2_9_left;
logic pe_2_9_mul_ready;
logic [31:0] pe_2_9_out;
logic pe_2_9_go;
logic pe_2_9_clk;
logic pe_2_9_reset;
logic pe_2_9_done;
logic [31:0] top_2_9_in;
logic top_2_9_write_en;
logic top_2_9_clk;
logic top_2_9_reset;
logic [31:0] top_2_9_out;
logic top_2_9_done;
logic [31:0] left_2_9_in;
logic left_2_9_write_en;
logic left_2_9_clk;
logic left_2_9_reset;
logic [31:0] left_2_9_out;
logic left_2_9_done;
logic [31:0] pe_2_10_top;
logic [31:0] pe_2_10_left;
logic pe_2_10_mul_ready;
logic [31:0] pe_2_10_out;
logic pe_2_10_go;
logic pe_2_10_clk;
logic pe_2_10_reset;
logic pe_2_10_done;
logic [31:0] top_2_10_in;
logic top_2_10_write_en;
logic top_2_10_clk;
logic top_2_10_reset;
logic [31:0] top_2_10_out;
logic top_2_10_done;
logic [31:0] left_2_10_in;
logic left_2_10_write_en;
logic left_2_10_clk;
logic left_2_10_reset;
logic [31:0] left_2_10_out;
logic left_2_10_done;
logic [31:0] pe_2_11_top;
logic [31:0] pe_2_11_left;
logic pe_2_11_mul_ready;
logic [31:0] pe_2_11_out;
logic pe_2_11_go;
logic pe_2_11_clk;
logic pe_2_11_reset;
logic pe_2_11_done;
logic [31:0] top_2_11_in;
logic top_2_11_write_en;
logic top_2_11_clk;
logic top_2_11_reset;
logic [31:0] top_2_11_out;
logic top_2_11_done;
logic [31:0] left_2_11_in;
logic left_2_11_write_en;
logic left_2_11_clk;
logic left_2_11_reset;
logic [31:0] left_2_11_out;
logic left_2_11_done;
logic [31:0] pe_2_12_top;
logic [31:0] pe_2_12_left;
logic pe_2_12_mul_ready;
logic [31:0] pe_2_12_out;
logic pe_2_12_go;
logic pe_2_12_clk;
logic pe_2_12_reset;
logic pe_2_12_done;
logic [31:0] top_2_12_in;
logic top_2_12_write_en;
logic top_2_12_clk;
logic top_2_12_reset;
logic [31:0] top_2_12_out;
logic top_2_12_done;
logic [31:0] left_2_12_in;
logic left_2_12_write_en;
logic left_2_12_clk;
logic left_2_12_reset;
logic [31:0] left_2_12_out;
logic left_2_12_done;
logic [31:0] pe_2_13_top;
logic [31:0] pe_2_13_left;
logic pe_2_13_mul_ready;
logic [31:0] pe_2_13_out;
logic pe_2_13_go;
logic pe_2_13_clk;
logic pe_2_13_reset;
logic pe_2_13_done;
logic [31:0] top_2_13_in;
logic top_2_13_write_en;
logic top_2_13_clk;
logic top_2_13_reset;
logic [31:0] top_2_13_out;
logic top_2_13_done;
logic [31:0] left_2_13_in;
logic left_2_13_write_en;
logic left_2_13_clk;
logic left_2_13_reset;
logic [31:0] left_2_13_out;
logic left_2_13_done;
logic [31:0] pe_2_14_top;
logic [31:0] pe_2_14_left;
logic pe_2_14_mul_ready;
logic [31:0] pe_2_14_out;
logic pe_2_14_go;
logic pe_2_14_clk;
logic pe_2_14_reset;
logic pe_2_14_done;
logic [31:0] top_2_14_in;
logic top_2_14_write_en;
logic top_2_14_clk;
logic top_2_14_reset;
logic [31:0] top_2_14_out;
logic top_2_14_done;
logic [31:0] left_2_14_in;
logic left_2_14_write_en;
logic left_2_14_clk;
logic left_2_14_reset;
logic [31:0] left_2_14_out;
logic left_2_14_done;
logic [31:0] pe_2_15_top;
logic [31:0] pe_2_15_left;
logic pe_2_15_mul_ready;
logic [31:0] pe_2_15_out;
logic pe_2_15_go;
logic pe_2_15_clk;
logic pe_2_15_reset;
logic pe_2_15_done;
logic [31:0] top_2_15_in;
logic top_2_15_write_en;
logic top_2_15_clk;
logic top_2_15_reset;
logic [31:0] top_2_15_out;
logic top_2_15_done;
logic [31:0] left_2_15_in;
logic left_2_15_write_en;
logic left_2_15_clk;
logic left_2_15_reset;
logic [31:0] left_2_15_out;
logic left_2_15_done;
logic [31:0] pe_3_0_top;
logic [31:0] pe_3_0_left;
logic pe_3_0_mul_ready;
logic [31:0] pe_3_0_out;
logic pe_3_0_go;
logic pe_3_0_clk;
logic pe_3_0_reset;
logic pe_3_0_done;
logic [31:0] top_3_0_in;
logic top_3_0_write_en;
logic top_3_0_clk;
logic top_3_0_reset;
logic [31:0] top_3_0_out;
logic top_3_0_done;
logic [31:0] left_3_0_in;
logic left_3_0_write_en;
logic left_3_0_clk;
logic left_3_0_reset;
logic [31:0] left_3_0_out;
logic left_3_0_done;
logic [31:0] pe_3_1_top;
logic [31:0] pe_3_1_left;
logic pe_3_1_mul_ready;
logic [31:0] pe_3_1_out;
logic pe_3_1_go;
logic pe_3_1_clk;
logic pe_3_1_reset;
logic pe_3_1_done;
logic [31:0] top_3_1_in;
logic top_3_1_write_en;
logic top_3_1_clk;
logic top_3_1_reset;
logic [31:0] top_3_1_out;
logic top_3_1_done;
logic [31:0] left_3_1_in;
logic left_3_1_write_en;
logic left_3_1_clk;
logic left_3_1_reset;
logic [31:0] left_3_1_out;
logic left_3_1_done;
logic [31:0] pe_3_2_top;
logic [31:0] pe_3_2_left;
logic pe_3_2_mul_ready;
logic [31:0] pe_3_2_out;
logic pe_3_2_go;
logic pe_3_2_clk;
logic pe_3_2_reset;
logic pe_3_2_done;
logic [31:0] top_3_2_in;
logic top_3_2_write_en;
logic top_3_2_clk;
logic top_3_2_reset;
logic [31:0] top_3_2_out;
logic top_3_2_done;
logic [31:0] left_3_2_in;
logic left_3_2_write_en;
logic left_3_2_clk;
logic left_3_2_reset;
logic [31:0] left_3_2_out;
logic left_3_2_done;
logic [31:0] pe_3_3_top;
logic [31:0] pe_3_3_left;
logic pe_3_3_mul_ready;
logic [31:0] pe_3_3_out;
logic pe_3_3_go;
logic pe_3_3_clk;
logic pe_3_3_reset;
logic pe_3_3_done;
logic [31:0] top_3_3_in;
logic top_3_3_write_en;
logic top_3_3_clk;
logic top_3_3_reset;
logic [31:0] top_3_3_out;
logic top_3_3_done;
logic [31:0] left_3_3_in;
logic left_3_3_write_en;
logic left_3_3_clk;
logic left_3_3_reset;
logic [31:0] left_3_3_out;
logic left_3_3_done;
logic [31:0] pe_3_4_top;
logic [31:0] pe_3_4_left;
logic pe_3_4_mul_ready;
logic [31:0] pe_3_4_out;
logic pe_3_4_go;
logic pe_3_4_clk;
logic pe_3_4_reset;
logic pe_3_4_done;
logic [31:0] top_3_4_in;
logic top_3_4_write_en;
logic top_3_4_clk;
logic top_3_4_reset;
logic [31:0] top_3_4_out;
logic top_3_4_done;
logic [31:0] left_3_4_in;
logic left_3_4_write_en;
logic left_3_4_clk;
logic left_3_4_reset;
logic [31:0] left_3_4_out;
logic left_3_4_done;
logic [31:0] pe_3_5_top;
logic [31:0] pe_3_5_left;
logic pe_3_5_mul_ready;
logic [31:0] pe_3_5_out;
logic pe_3_5_go;
logic pe_3_5_clk;
logic pe_3_5_reset;
logic pe_3_5_done;
logic [31:0] top_3_5_in;
logic top_3_5_write_en;
logic top_3_5_clk;
logic top_3_5_reset;
logic [31:0] top_3_5_out;
logic top_3_5_done;
logic [31:0] left_3_5_in;
logic left_3_5_write_en;
logic left_3_5_clk;
logic left_3_5_reset;
logic [31:0] left_3_5_out;
logic left_3_5_done;
logic [31:0] pe_3_6_top;
logic [31:0] pe_3_6_left;
logic pe_3_6_mul_ready;
logic [31:0] pe_3_6_out;
logic pe_3_6_go;
logic pe_3_6_clk;
logic pe_3_6_reset;
logic pe_3_6_done;
logic [31:0] top_3_6_in;
logic top_3_6_write_en;
logic top_3_6_clk;
logic top_3_6_reset;
logic [31:0] top_3_6_out;
logic top_3_6_done;
logic [31:0] left_3_6_in;
logic left_3_6_write_en;
logic left_3_6_clk;
logic left_3_6_reset;
logic [31:0] left_3_6_out;
logic left_3_6_done;
logic [31:0] pe_3_7_top;
logic [31:0] pe_3_7_left;
logic pe_3_7_mul_ready;
logic [31:0] pe_3_7_out;
logic pe_3_7_go;
logic pe_3_7_clk;
logic pe_3_7_reset;
logic pe_3_7_done;
logic [31:0] top_3_7_in;
logic top_3_7_write_en;
logic top_3_7_clk;
logic top_3_7_reset;
logic [31:0] top_3_7_out;
logic top_3_7_done;
logic [31:0] left_3_7_in;
logic left_3_7_write_en;
logic left_3_7_clk;
logic left_3_7_reset;
logic [31:0] left_3_7_out;
logic left_3_7_done;
logic [31:0] pe_3_8_top;
logic [31:0] pe_3_8_left;
logic pe_3_8_mul_ready;
logic [31:0] pe_3_8_out;
logic pe_3_8_go;
logic pe_3_8_clk;
logic pe_3_8_reset;
logic pe_3_8_done;
logic [31:0] top_3_8_in;
logic top_3_8_write_en;
logic top_3_8_clk;
logic top_3_8_reset;
logic [31:0] top_3_8_out;
logic top_3_8_done;
logic [31:0] left_3_8_in;
logic left_3_8_write_en;
logic left_3_8_clk;
logic left_3_8_reset;
logic [31:0] left_3_8_out;
logic left_3_8_done;
logic [31:0] pe_3_9_top;
logic [31:0] pe_3_9_left;
logic pe_3_9_mul_ready;
logic [31:0] pe_3_9_out;
logic pe_3_9_go;
logic pe_3_9_clk;
logic pe_3_9_reset;
logic pe_3_9_done;
logic [31:0] top_3_9_in;
logic top_3_9_write_en;
logic top_3_9_clk;
logic top_3_9_reset;
logic [31:0] top_3_9_out;
logic top_3_9_done;
logic [31:0] left_3_9_in;
logic left_3_9_write_en;
logic left_3_9_clk;
logic left_3_9_reset;
logic [31:0] left_3_9_out;
logic left_3_9_done;
logic [31:0] pe_3_10_top;
logic [31:0] pe_3_10_left;
logic pe_3_10_mul_ready;
logic [31:0] pe_3_10_out;
logic pe_3_10_go;
logic pe_3_10_clk;
logic pe_3_10_reset;
logic pe_3_10_done;
logic [31:0] top_3_10_in;
logic top_3_10_write_en;
logic top_3_10_clk;
logic top_3_10_reset;
logic [31:0] top_3_10_out;
logic top_3_10_done;
logic [31:0] left_3_10_in;
logic left_3_10_write_en;
logic left_3_10_clk;
logic left_3_10_reset;
logic [31:0] left_3_10_out;
logic left_3_10_done;
logic [31:0] pe_3_11_top;
logic [31:0] pe_3_11_left;
logic pe_3_11_mul_ready;
logic [31:0] pe_3_11_out;
logic pe_3_11_go;
logic pe_3_11_clk;
logic pe_3_11_reset;
logic pe_3_11_done;
logic [31:0] top_3_11_in;
logic top_3_11_write_en;
logic top_3_11_clk;
logic top_3_11_reset;
logic [31:0] top_3_11_out;
logic top_3_11_done;
logic [31:0] left_3_11_in;
logic left_3_11_write_en;
logic left_3_11_clk;
logic left_3_11_reset;
logic [31:0] left_3_11_out;
logic left_3_11_done;
logic [31:0] pe_3_12_top;
logic [31:0] pe_3_12_left;
logic pe_3_12_mul_ready;
logic [31:0] pe_3_12_out;
logic pe_3_12_go;
logic pe_3_12_clk;
logic pe_3_12_reset;
logic pe_3_12_done;
logic [31:0] top_3_12_in;
logic top_3_12_write_en;
logic top_3_12_clk;
logic top_3_12_reset;
logic [31:0] top_3_12_out;
logic top_3_12_done;
logic [31:0] left_3_12_in;
logic left_3_12_write_en;
logic left_3_12_clk;
logic left_3_12_reset;
logic [31:0] left_3_12_out;
logic left_3_12_done;
logic [31:0] pe_3_13_top;
logic [31:0] pe_3_13_left;
logic pe_3_13_mul_ready;
logic [31:0] pe_3_13_out;
logic pe_3_13_go;
logic pe_3_13_clk;
logic pe_3_13_reset;
logic pe_3_13_done;
logic [31:0] top_3_13_in;
logic top_3_13_write_en;
logic top_3_13_clk;
logic top_3_13_reset;
logic [31:0] top_3_13_out;
logic top_3_13_done;
logic [31:0] left_3_13_in;
logic left_3_13_write_en;
logic left_3_13_clk;
logic left_3_13_reset;
logic [31:0] left_3_13_out;
logic left_3_13_done;
logic [31:0] pe_3_14_top;
logic [31:0] pe_3_14_left;
logic pe_3_14_mul_ready;
logic [31:0] pe_3_14_out;
logic pe_3_14_go;
logic pe_3_14_clk;
logic pe_3_14_reset;
logic pe_3_14_done;
logic [31:0] top_3_14_in;
logic top_3_14_write_en;
logic top_3_14_clk;
logic top_3_14_reset;
logic [31:0] top_3_14_out;
logic top_3_14_done;
logic [31:0] left_3_14_in;
logic left_3_14_write_en;
logic left_3_14_clk;
logic left_3_14_reset;
logic [31:0] left_3_14_out;
logic left_3_14_done;
logic [31:0] pe_3_15_top;
logic [31:0] pe_3_15_left;
logic pe_3_15_mul_ready;
logic [31:0] pe_3_15_out;
logic pe_3_15_go;
logic pe_3_15_clk;
logic pe_3_15_reset;
logic pe_3_15_done;
logic [31:0] top_3_15_in;
logic top_3_15_write_en;
logic top_3_15_clk;
logic top_3_15_reset;
logic [31:0] top_3_15_out;
logic top_3_15_done;
logic [31:0] left_3_15_in;
logic left_3_15_write_en;
logic left_3_15_clk;
logic left_3_15_reset;
logic [31:0] left_3_15_out;
logic left_3_15_done;
logic [31:0] pe_4_0_top;
logic [31:0] pe_4_0_left;
logic pe_4_0_mul_ready;
logic [31:0] pe_4_0_out;
logic pe_4_0_go;
logic pe_4_0_clk;
logic pe_4_0_reset;
logic pe_4_0_done;
logic [31:0] top_4_0_in;
logic top_4_0_write_en;
logic top_4_0_clk;
logic top_4_0_reset;
logic [31:0] top_4_0_out;
logic top_4_0_done;
logic [31:0] left_4_0_in;
logic left_4_0_write_en;
logic left_4_0_clk;
logic left_4_0_reset;
logic [31:0] left_4_0_out;
logic left_4_0_done;
logic [31:0] pe_4_1_top;
logic [31:0] pe_4_1_left;
logic pe_4_1_mul_ready;
logic [31:0] pe_4_1_out;
logic pe_4_1_go;
logic pe_4_1_clk;
logic pe_4_1_reset;
logic pe_4_1_done;
logic [31:0] top_4_1_in;
logic top_4_1_write_en;
logic top_4_1_clk;
logic top_4_1_reset;
logic [31:0] top_4_1_out;
logic top_4_1_done;
logic [31:0] left_4_1_in;
logic left_4_1_write_en;
logic left_4_1_clk;
logic left_4_1_reset;
logic [31:0] left_4_1_out;
logic left_4_1_done;
logic [31:0] pe_4_2_top;
logic [31:0] pe_4_2_left;
logic pe_4_2_mul_ready;
logic [31:0] pe_4_2_out;
logic pe_4_2_go;
logic pe_4_2_clk;
logic pe_4_2_reset;
logic pe_4_2_done;
logic [31:0] top_4_2_in;
logic top_4_2_write_en;
logic top_4_2_clk;
logic top_4_2_reset;
logic [31:0] top_4_2_out;
logic top_4_2_done;
logic [31:0] left_4_2_in;
logic left_4_2_write_en;
logic left_4_2_clk;
logic left_4_2_reset;
logic [31:0] left_4_2_out;
logic left_4_2_done;
logic [31:0] pe_4_3_top;
logic [31:0] pe_4_3_left;
logic pe_4_3_mul_ready;
logic [31:0] pe_4_3_out;
logic pe_4_3_go;
logic pe_4_3_clk;
logic pe_4_3_reset;
logic pe_4_3_done;
logic [31:0] top_4_3_in;
logic top_4_3_write_en;
logic top_4_3_clk;
logic top_4_3_reset;
logic [31:0] top_4_3_out;
logic top_4_3_done;
logic [31:0] left_4_3_in;
logic left_4_3_write_en;
logic left_4_3_clk;
logic left_4_3_reset;
logic [31:0] left_4_3_out;
logic left_4_3_done;
logic [31:0] pe_4_4_top;
logic [31:0] pe_4_4_left;
logic pe_4_4_mul_ready;
logic [31:0] pe_4_4_out;
logic pe_4_4_go;
logic pe_4_4_clk;
logic pe_4_4_reset;
logic pe_4_4_done;
logic [31:0] top_4_4_in;
logic top_4_4_write_en;
logic top_4_4_clk;
logic top_4_4_reset;
logic [31:0] top_4_4_out;
logic top_4_4_done;
logic [31:0] left_4_4_in;
logic left_4_4_write_en;
logic left_4_4_clk;
logic left_4_4_reset;
logic [31:0] left_4_4_out;
logic left_4_4_done;
logic [31:0] pe_4_5_top;
logic [31:0] pe_4_5_left;
logic pe_4_5_mul_ready;
logic [31:0] pe_4_5_out;
logic pe_4_5_go;
logic pe_4_5_clk;
logic pe_4_5_reset;
logic pe_4_5_done;
logic [31:0] top_4_5_in;
logic top_4_5_write_en;
logic top_4_5_clk;
logic top_4_5_reset;
logic [31:0] top_4_5_out;
logic top_4_5_done;
logic [31:0] left_4_5_in;
logic left_4_5_write_en;
logic left_4_5_clk;
logic left_4_5_reset;
logic [31:0] left_4_5_out;
logic left_4_5_done;
logic [31:0] pe_4_6_top;
logic [31:0] pe_4_6_left;
logic pe_4_6_mul_ready;
logic [31:0] pe_4_6_out;
logic pe_4_6_go;
logic pe_4_6_clk;
logic pe_4_6_reset;
logic pe_4_6_done;
logic [31:0] top_4_6_in;
logic top_4_6_write_en;
logic top_4_6_clk;
logic top_4_6_reset;
logic [31:0] top_4_6_out;
logic top_4_6_done;
logic [31:0] left_4_6_in;
logic left_4_6_write_en;
logic left_4_6_clk;
logic left_4_6_reset;
logic [31:0] left_4_6_out;
logic left_4_6_done;
logic [31:0] pe_4_7_top;
logic [31:0] pe_4_7_left;
logic pe_4_7_mul_ready;
logic [31:0] pe_4_7_out;
logic pe_4_7_go;
logic pe_4_7_clk;
logic pe_4_7_reset;
logic pe_4_7_done;
logic [31:0] top_4_7_in;
logic top_4_7_write_en;
logic top_4_7_clk;
logic top_4_7_reset;
logic [31:0] top_4_7_out;
logic top_4_7_done;
logic [31:0] left_4_7_in;
logic left_4_7_write_en;
logic left_4_7_clk;
logic left_4_7_reset;
logic [31:0] left_4_7_out;
logic left_4_7_done;
logic [31:0] pe_4_8_top;
logic [31:0] pe_4_8_left;
logic pe_4_8_mul_ready;
logic [31:0] pe_4_8_out;
logic pe_4_8_go;
logic pe_4_8_clk;
logic pe_4_8_reset;
logic pe_4_8_done;
logic [31:0] top_4_8_in;
logic top_4_8_write_en;
logic top_4_8_clk;
logic top_4_8_reset;
logic [31:0] top_4_8_out;
logic top_4_8_done;
logic [31:0] left_4_8_in;
logic left_4_8_write_en;
logic left_4_8_clk;
logic left_4_8_reset;
logic [31:0] left_4_8_out;
logic left_4_8_done;
logic [31:0] pe_4_9_top;
logic [31:0] pe_4_9_left;
logic pe_4_9_mul_ready;
logic [31:0] pe_4_9_out;
logic pe_4_9_go;
logic pe_4_9_clk;
logic pe_4_9_reset;
logic pe_4_9_done;
logic [31:0] top_4_9_in;
logic top_4_9_write_en;
logic top_4_9_clk;
logic top_4_9_reset;
logic [31:0] top_4_9_out;
logic top_4_9_done;
logic [31:0] left_4_9_in;
logic left_4_9_write_en;
logic left_4_9_clk;
logic left_4_9_reset;
logic [31:0] left_4_9_out;
logic left_4_9_done;
logic [31:0] pe_4_10_top;
logic [31:0] pe_4_10_left;
logic pe_4_10_mul_ready;
logic [31:0] pe_4_10_out;
logic pe_4_10_go;
logic pe_4_10_clk;
logic pe_4_10_reset;
logic pe_4_10_done;
logic [31:0] top_4_10_in;
logic top_4_10_write_en;
logic top_4_10_clk;
logic top_4_10_reset;
logic [31:0] top_4_10_out;
logic top_4_10_done;
logic [31:0] left_4_10_in;
logic left_4_10_write_en;
logic left_4_10_clk;
logic left_4_10_reset;
logic [31:0] left_4_10_out;
logic left_4_10_done;
logic [31:0] pe_4_11_top;
logic [31:0] pe_4_11_left;
logic pe_4_11_mul_ready;
logic [31:0] pe_4_11_out;
logic pe_4_11_go;
logic pe_4_11_clk;
logic pe_4_11_reset;
logic pe_4_11_done;
logic [31:0] top_4_11_in;
logic top_4_11_write_en;
logic top_4_11_clk;
logic top_4_11_reset;
logic [31:0] top_4_11_out;
logic top_4_11_done;
logic [31:0] left_4_11_in;
logic left_4_11_write_en;
logic left_4_11_clk;
logic left_4_11_reset;
logic [31:0] left_4_11_out;
logic left_4_11_done;
logic [31:0] pe_4_12_top;
logic [31:0] pe_4_12_left;
logic pe_4_12_mul_ready;
logic [31:0] pe_4_12_out;
logic pe_4_12_go;
logic pe_4_12_clk;
logic pe_4_12_reset;
logic pe_4_12_done;
logic [31:0] top_4_12_in;
logic top_4_12_write_en;
logic top_4_12_clk;
logic top_4_12_reset;
logic [31:0] top_4_12_out;
logic top_4_12_done;
logic [31:0] left_4_12_in;
logic left_4_12_write_en;
logic left_4_12_clk;
logic left_4_12_reset;
logic [31:0] left_4_12_out;
logic left_4_12_done;
logic [31:0] pe_4_13_top;
logic [31:0] pe_4_13_left;
logic pe_4_13_mul_ready;
logic [31:0] pe_4_13_out;
logic pe_4_13_go;
logic pe_4_13_clk;
logic pe_4_13_reset;
logic pe_4_13_done;
logic [31:0] top_4_13_in;
logic top_4_13_write_en;
logic top_4_13_clk;
logic top_4_13_reset;
logic [31:0] top_4_13_out;
logic top_4_13_done;
logic [31:0] left_4_13_in;
logic left_4_13_write_en;
logic left_4_13_clk;
logic left_4_13_reset;
logic [31:0] left_4_13_out;
logic left_4_13_done;
logic [31:0] pe_4_14_top;
logic [31:0] pe_4_14_left;
logic pe_4_14_mul_ready;
logic [31:0] pe_4_14_out;
logic pe_4_14_go;
logic pe_4_14_clk;
logic pe_4_14_reset;
logic pe_4_14_done;
logic [31:0] top_4_14_in;
logic top_4_14_write_en;
logic top_4_14_clk;
logic top_4_14_reset;
logic [31:0] top_4_14_out;
logic top_4_14_done;
logic [31:0] left_4_14_in;
logic left_4_14_write_en;
logic left_4_14_clk;
logic left_4_14_reset;
logic [31:0] left_4_14_out;
logic left_4_14_done;
logic [31:0] pe_4_15_top;
logic [31:0] pe_4_15_left;
logic pe_4_15_mul_ready;
logic [31:0] pe_4_15_out;
logic pe_4_15_go;
logic pe_4_15_clk;
logic pe_4_15_reset;
logic pe_4_15_done;
logic [31:0] top_4_15_in;
logic top_4_15_write_en;
logic top_4_15_clk;
logic top_4_15_reset;
logic [31:0] top_4_15_out;
logic top_4_15_done;
logic [31:0] left_4_15_in;
logic left_4_15_write_en;
logic left_4_15_clk;
logic left_4_15_reset;
logic [31:0] left_4_15_out;
logic left_4_15_done;
logic [31:0] pe_5_0_top;
logic [31:0] pe_5_0_left;
logic pe_5_0_mul_ready;
logic [31:0] pe_5_0_out;
logic pe_5_0_go;
logic pe_5_0_clk;
logic pe_5_0_reset;
logic pe_5_0_done;
logic [31:0] top_5_0_in;
logic top_5_0_write_en;
logic top_5_0_clk;
logic top_5_0_reset;
logic [31:0] top_5_0_out;
logic top_5_0_done;
logic [31:0] left_5_0_in;
logic left_5_0_write_en;
logic left_5_0_clk;
logic left_5_0_reset;
logic [31:0] left_5_0_out;
logic left_5_0_done;
logic [31:0] pe_5_1_top;
logic [31:0] pe_5_1_left;
logic pe_5_1_mul_ready;
logic [31:0] pe_5_1_out;
logic pe_5_1_go;
logic pe_5_1_clk;
logic pe_5_1_reset;
logic pe_5_1_done;
logic [31:0] top_5_1_in;
logic top_5_1_write_en;
logic top_5_1_clk;
logic top_5_1_reset;
logic [31:0] top_5_1_out;
logic top_5_1_done;
logic [31:0] left_5_1_in;
logic left_5_1_write_en;
logic left_5_1_clk;
logic left_5_1_reset;
logic [31:0] left_5_1_out;
logic left_5_1_done;
logic [31:0] pe_5_2_top;
logic [31:0] pe_5_2_left;
logic pe_5_2_mul_ready;
logic [31:0] pe_5_2_out;
logic pe_5_2_go;
logic pe_5_2_clk;
logic pe_5_2_reset;
logic pe_5_2_done;
logic [31:0] top_5_2_in;
logic top_5_2_write_en;
logic top_5_2_clk;
logic top_5_2_reset;
logic [31:0] top_5_2_out;
logic top_5_2_done;
logic [31:0] left_5_2_in;
logic left_5_2_write_en;
logic left_5_2_clk;
logic left_5_2_reset;
logic [31:0] left_5_2_out;
logic left_5_2_done;
logic [31:0] pe_5_3_top;
logic [31:0] pe_5_3_left;
logic pe_5_3_mul_ready;
logic [31:0] pe_5_3_out;
logic pe_5_3_go;
logic pe_5_3_clk;
logic pe_5_3_reset;
logic pe_5_3_done;
logic [31:0] top_5_3_in;
logic top_5_3_write_en;
logic top_5_3_clk;
logic top_5_3_reset;
logic [31:0] top_5_3_out;
logic top_5_3_done;
logic [31:0] left_5_3_in;
logic left_5_3_write_en;
logic left_5_3_clk;
logic left_5_3_reset;
logic [31:0] left_5_3_out;
logic left_5_3_done;
logic [31:0] pe_5_4_top;
logic [31:0] pe_5_4_left;
logic pe_5_4_mul_ready;
logic [31:0] pe_5_4_out;
logic pe_5_4_go;
logic pe_5_4_clk;
logic pe_5_4_reset;
logic pe_5_4_done;
logic [31:0] top_5_4_in;
logic top_5_4_write_en;
logic top_5_4_clk;
logic top_5_4_reset;
logic [31:0] top_5_4_out;
logic top_5_4_done;
logic [31:0] left_5_4_in;
logic left_5_4_write_en;
logic left_5_4_clk;
logic left_5_4_reset;
logic [31:0] left_5_4_out;
logic left_5_4_done;
logic [31:0] pe_5_5_top;
logic [31:0] pe_5_5_left;
logic pe_5_5_mul_ready;
logic [31:0] pe_5_5_out;
logic pe_5_5_go;
logic pe_5_5_clk;
logic pe_5_5_reset;
logic pe_5_5_done;
logic [31:0] top_5_5_in;
logic top_5_5_write_en;
logic top_5_5_clk;
logic top_5_5_reset;
logic [31:0] top_5_5_out;
logic top_5_5_done;
logic [31:0] left_5_5_in;
logic left_5_5_write_en;
logic left_5_5_clk;
logic left_5_5_reset;
logic [31:0] left_5_5_out;
logic left_5_5_done;
logic [31:0] pe_5_6_top;
logic [31:0] pe_5_6_left;
logic pe_5_6_mul_ready;
logic [31:0] pe_5_6_out;
logic pe_5_6_go;
logic pe_5_6_clk;
logic pe_5_6_reset;
logic pe_5_6_done;
logic [31:0] top_5_6_in;
logic top_5_6_write_en;
logic top_5_6_clk;
logic top_5_6_reset;
logic [31:0] top_5_6_out;
logic top_5_6_done;
logic [31:0] left_5_6_in;
logic left_5_6_write_en;
logic left_5_6_clk;
logic left_5_6_reset;
logic [31:0] left_5_6_out;
logic left_5_6_done;
logic [31:0] pe_5_7_top;
logic [31:0] pe_5_7_left;
logic pe_5_7_mul_ready;
logic [31:0] pe_5_7_out;
logic pe_5_7_go;
logic pe_5_7_clk;
logic pe_5_7_reset;
logic pe_5_7_done;
logic [31:0] top_5_7_in;
logic top_5_7_write_en;
logic top_5_7_clk;
logic top_5_7_reset;
logic [31:0] top_5_7_out;
logic top_5_7_done;
logic [31:0] left_5_7_in;
logic left_5_7_write_en;
logic left_5_7_clk;
logic left_5_7_reset;
logic [31:0] left_5_7_out;
logic left_5_7_done;
logic [31:0] pe_5_8_top;
logic [31:0] pe_5_8_left;
logic pe_5_8_mul_ready;
logic [31:0] pe_5_8_out;
logic pe_5_8_go;
logic pe_5_8_clk;
logic pe_5_8_reset;
logic pe_5_8_done;
logic [31:0] top_5_8_in;
logic top_5_8_write_en;
logic top_5_8_clk;
logic top_5_8_reset;
logic [31:0] top_5_8_out;
logic top_5_8_done;
logic [31:0] left_5_8_in;
logic left_5_8_write_en;
logic left_5_8_clk;
logic left_5_8_reset;
logic [31:0] left_5_8_out;
logic left_5_8_done;
logic [31:0] pe_5_9_top;
logic [31:0] pe_5_9_left;
logic pe_5_9_mul_ready;
logic [31:0] pe_5_9_out;
logic pe_5_9_go;
logic pe_5_9_clk;
logic pe_5_9_reset;
logic pe_5_9_done;
logic [31:0] top_5_9_in;
logic top_5_9_write_en;
logic top_5_9_clk;
logic top_5_9_reset;
logic [31:0] top_5_9_out;
logic top_5_9_done;
logic [31:0] left_5_9_in;
logic left_5_9_write_en;
logic left_5_9_clk;
logic left_5_9_reset;
logic [31:0] left_5_9_out;
logic left_5_9_done;
logic [31:0] pe_5_10_top;
logic [31:0] pe_5_10_left;
logic pe_5_10_mul_ready;
logic [31:0] pe_5_10_out;
logic pe_5_10_go;
logic pe_5_10_clk;
logic pe_5_10_reset;
logic pe_5_10_done;
logic [31:0] top_5_10_in;
logic top_5_10_write_en;
logic top_5_10_clk;
logic top_5_10_reset;
logic [31:0] top_5_10_out;
logic top_5_10_done;
logic [31:0] left_5_10_in;
logic left_5_10_write_en;
logic left_5_10_clk;
logic left_5_10_reset;
logic [31:0] left_5_10_out;
logic left_5_10_done;
logic [31:0] pe_5_11_top;
logic [31:0] pe_5_11_left;
logic pe_5_11_mul_ready;
logic [31:0] pe_5_11_out;
logic pe_5_11_go;
logic pe_5_11_clk;
logic pe_5_11_reset;
logic pe_5_11_done;
logic [31:0] top_5_11_in;
logic top_5_11_write_en;
logic top_5_11_clk;
logic top_5_11_reset;
logic [31:0] top_5_11_out;
logic top_5_11_done;
logic [31:0] left_5_11_in;
logic left_5_11_write_en;
logic left_5_11_clk;
logic left_5_11_reset;
logic [31:0] left_5_11_out;
logic left_5_11_done;
logic [31:0] pe_5_12_top;
logic [31:0] pe_5_12_left;
logic pe_5_12_mul_ready;
logic [31:0] pe_5_12_out;
logic pe_5_12_go;
logic pe_5_12_clk;
logic pe_5_12_reset;
logic pe_5_12_done;
logic [31:0] top_5_12_in;
logic top_5_12_write_en;
logic top_5_12_clk;
logic top_5_12_reset;
logic [31:0] top_5_12_out;
logic top_5_12_done;
logic [31:0] left_5_12_in;
logic left_5_12_write_en;
logic left_5_12_clk;
logic left_5_12_reset;
logic [31:0] left_5_12_out;
logic left_5_12_done;
logic [31:0] pe_5_13_top;
logic [31:0] pe_5_13_left;
logic pe_5_13_mul_ready;
logic [31:0] pe_5_13_out;
logic pe_5_13_go;
logic pe_5_13_clk;
logic pe_5_13_reset;
logic pe_5_13_done;
logic [31:0] top_5_13_in;
logic top_5_13_write_en;
logic top_5_13_clk;
logic top_5_13_reset;
logic [31:0] top_5_13_out;
logic top_5_13_done;
logic [31:0] left_5_13_in;
logic left_5_13_write_en;
logic left_5_13_clk;
logic left_5_13_reset;
logic [31:0] left_5_13_out;
logic left_5_13_done;
logic [31:0] pe_5_14_top;
logic [31:0] pe_5_14_left;
logic pe_5_14_mul_ready;
logic [31:0] pe_5_14_out;
logic pe_5_14_go;
logic pe_5_14_clk;
logic pe_5_14_reset;
logic pe_5_14_done;
logic [31:0] top_5_14_in;
logic top_5_14_write_en;
logic top_5_14_clk;
logic top_5_14_reset;
logic [31:0] top_5_14_out;
logic top_5_14_done;
logic [31:0] left_5_14_in;
logic left_5_14_write_en;
logic left_5_14_clk;
logic left_5_14_reset;
logic [31:0] left_5_14_out;
logic left_5_14_done;
logic [31:0] pe_5_15_top;
logic [31:0] pe_5_15_left;
logic pe_5_15_mul_ready;
logic [31:0] pe_5_15_out;
logic pe_5_15_go;
logic pe_5_15_clk;
logic pe_5_15_reset;
logic pe_5_15_done;
logic [31:0] top_5_15_in;
logic top_5_15_write_en;
logic top_5_15_clk;
logic top_5_15_reset;
logic [31:0] top_5_15_out;
logic top_5_15_done;
logic [31:0] left_5_15_in;
logic left_5_15_write_en;
logic left_5_15_clk;
logic left_5_15_reset;
logic [31:0] left_5_15_out;
logic left_5_15_done;
logic [31:0] pe_6_0_top;
logic [31:0] pe_6_0_left;
logic pe_6_0_mul_ready;
logic [31:0] pe_6_0_out;
logic pe_6_0_go;
logic pe_6_0_clk;
logic pe_6_0_reset;
logic pe_6_0_done;
logic [31:0] top_6_0_in;
logic top_6_0_write_en;
logic top_6_0_clk;
logic top_6_0_reset;
logic [31:0] top_6_0_out;
logic top_6_0_done;
logic [31:0] left_6_0_in;
logic left_6_0_write_en;
logic left_6_0_clk;
logic left_6_0_reset;
logic [31:0] left_6_0_out;
logic left_6_0_done;
logic [31:0] pe_6_1_top;
logic [31:0] pe_6_1_left;
logic pe_6_1_mul_ready;
logic [31:0] pe_6_1_out;
logic pe_6_1_go;
logic pe_6_1_clk;
logic pe_6_1_reset;
logic pe_6_1_done;
logic [31:0] top_6_1_in;
logic top_6_1_write_en;
logic top_6_1_clk;
logic top_6_1_reset;
logic [31:0] top_6_1_out;
logic top_6_1_done;
logic [31:0] left_6_1_in;
logic left_6_1_write_en;
logic left_6_1_clk;
logic left_6_1_reset;
logic [31:0] left_6_1_out;
logic left_6_1_done;
logic [31:0] pe_6_2_top;
logic [31:0] pe_6_2_left;
logic pe_6_2_mul_ready;
logic [31:0] pe_6_2_out;
logic pe_6_2_go;
logic pe_6_2_clk;
logic pe_6_2_reset;
logic pe_6_2_done;
logic [31:0] top_6_2_in;
logic top_6_2_write_en;
logic top_6_2_clk;
logic top_6_2_reset;
logic [31:0] top_6_2_out;
logic top_6_2_done;
logic [31:0] left_6_2_in;
logic left_6_2_write_en;
logic left_6_2_clk;
logic left_6_2_reset;
logic [31:0] left_6_2_out;
logic left_6_2_done;
logic [31:0] pe_6_3_top;
logic [31:0] pe_6_3_left;
logic pe_6_3_mul_ready;
logic [31:0] pe_6_3_out;
logic pe_6_3_go;
logic pe_6_3_clk;
logic pe_6_3_reset;
logic pe_6_3_done;
logic [31:0] top_6_3_in;
logic top_6_3_write_en;
logic top_6_3_clk;
logic top_6_3_reset;
logic [31:0] top_6_3_out;
logic top_6_3_done;
logic [31:0] left_6_3_in;
logic left_6_3_write_en;
logic left_6_3_clk;
logic left_6_3_reset;
logic [31:0] left_6_3_out;
logic left_6_3_done;
logic [31:0] pe_6_4_top;
logic [31:0] pe_6_4_left;
logic pe_6_4_mul_ready;
logic [31:0] pe_6_4_out;
logic pe_6_4_go;
logic pe_6_4_clk;
logic pe_6_4_reset;
logic pe_6_4_done;
logic [31:0] top_6_4_in;
logic top_6_4_write_en;
logic top_6_4_clk;
logic top_6_4_reset;
logic [31:0] top_6_4_out;
logic top_6_4_done;
logic [31:0] left_6_4_in;
logic left_6_4_write_en;
logic left_6_4_clk;
logic left_6_4_reset;
logic [31:0] left_6_4_out;
logic left_6_4_done;
logic [31:0] pe_6_5_top;
logic [31:0] pe_6_5_left;
logic pe_6_5_mul_ready;
logic [31:0] pe_6_5_out;
logic pe_6_5_go;
logic pe_6_5_clk;
logic pe_6_5_reset;
logic pe_6_5_done;
logic [31:0] top_6_5_in;
logic top_6_5_write_en;
logic top_6_5_clk;
logic top_6_5_reset;
logic [31:0] top_6_5_out;
logic top_6_5_done;
logic [31:0] left_6_5_in;
logic left_6_5_write_en;
logic left_6_5_clk;
logic left_6_5_reset;
logic [31:0] left_6_5_out;
logic left_6_5_done;
logic [31:0] pe_6_6_top;
logic [31:0] pe_6_6_left;
logic pe_6_6_mul_ready;
logic [31:0] pe_6_6_out;
logic pe_6_6_go;
logic pe_6_6_clk;
logic pe_6_6_reset;
logic pe_6_6_done;
logic [31:0] top_6_6_in;
logic top_6_6_write_en;
logic top_6_6_clk;
logic top_6_6_reset;
logic [31:0] top_6_6_out;
logic top_6_6_done;
logic [31:0] left_6_6_in;
logic left_6_6_write_en;
logic left_6_6_clk;
logic left_6_6_reset;
logic [31:0] left_6_6_out;
logic left_6_6_done;
logic [31:0] pe_6_7_top;
logic [31:0] pe_6_7_left;
logic pe_6_7_mul_ready;
logic [31:0] pe_6_7_out;
logic pe_6_7_go;
logic pe_6_7_clk;
logic pe_6_7_reset;
logic pe_6_7_done;
logic [31:0] top_6_7_in;
logic top_6_7_write_en;
logic top_6_7_clk;
logic top_6_7_reset;
logic [31:0] top_6_7_out;
logic top_6_7_done;
logic [31:0] left_6_7_in;
logic left_6_7_write_en;
logic left_6_7_clk;
logic left_6_7_reset;
logic [31:0] left_6_7_out;
logic left_6_7_done;
logic [31:0] pe_6_8_top;
logic [31:0] pe_6_8_left;
logic pe_6_8_mul_ready;
logic [31:0] pe_6_8_out;
logic pe_6_8_go;
logic pe_6_8_clk;
logic pe_6_8_reset;
logic pe_6_8_done;
logic [31:0] top_6_8_in;
logic top_6_8_write_en;
logic top_6_8_clk;
logic top_6_8_reset;
logic [31:0] top_6_8_out;
logic top_6_8_done;
logic [31:0] left_6_8_in;
logic left_6_8_write_en;
logic left_6_8_clk;
logic left_6_8_reset;
logic [31:0] left_6_8_out;
logic left_6_8_done;
logic [31:0] pe_6_9_top;
logic [31:0] pe_6_9_left;
logic pe_6_9_mul_ready;
logic [31:0] pe_6_9_out;
logic pe_6_9_go;
logic pe_6_9_clk;
logic pe_6_9_reset;
logic pe_6_9_done;
logic [31:0] top_6_9_in;
logic top_6_9_write_en;
logic top_6_9_clk;
logic top_6_9_reset;
logic [31:0] top_6_9_out;
logic top_6_9_done;
logic [31:0] left_6_9_in;
logic left_6_9_write_en;
logic left_6_9_clk;
logic left_6_9_reset;
logic [31:0] left_6_9_out;
logic left_6_9_done;
logic [31:0] pe_6_10_top;
logic [31:0] pe_6_10_left;
logic pe_6_10_mul_ready;
logic [31:0] pe_6_10_out;
logic pe_6_10_go;
logic pe_6_10_clk;
logic pe_6_10_reset;
logic pe_6_10_done;
logic [31:0] top_6_10_in;
logic top_6_10_write_en;
logic top_6_10_clk;
logic top_6_10_reset;
logic [31:0] top_6_10_out;
logic top_6_10_done;
logic [31:0] left_6_10_in;
logic left_6_10_write_en;
logic left_6_10_clk;
logic left_6_10_reset;
logic [31:0] left_6_10_out;
logic left_6_10_done;
logic [31:0] pe_6_11_top;
logic [31:0] pe_6_11_left;
logic pe_6_11_mul_ready;
logic [31:0] pe_6_11_out;
logic pe_6_11_go;
logic pe_6_11_clk;
logic pe_6_11_reset;
logic pe_6_11_done;
logic [31:0] top_6_11_in;
logic top_6_11_write_en;
logic top_6_11_clk;
logic top_6_11_reset;
logic [31:0] top_6_11_out;
logic top_6_11_done;
logic [31:0] left_6_11_in;
logic left_6_11_write_en;
logic left_6_11_clk;
logic left_6_11_reset;
logic [31:0] left_6_11_out;
logic left_6_11_done;
logic [31:0] pe_6_12_top;
logic [31:0] pe_6_12_left;
logic pe_6_12_mul_ready;
logic [31:0] pe_6_12_out;
logic pe_6_12_go;
logic pe_6_12_clk;
logic pe_6_12_reset;
logic pe_6_12_done;
logic [31:0] top_6_12_in;
logic top_6_12_write_en;
logic top_6_12_clk;
logic top_6_12_reset;
logic [31:0] top_6_12_out;
logic top_6_12_done;
logic [31:0] left_6_12_in;
logic left_6_12_write_en;
logic left_6_12_clk;
logic left_6_12_reset;
logic [31:0] left_6_12_out;
logic left_6_12_done;
logic [31:0] pe_6_13_top;
logic [31:0] pe_6_13_left;
logic pe_6_13_mul_ready;
logic [31:0] pe_6_13_out;
logic pe_6_13_go;
logic pe_6_13_clk;
logic pe_6_13_reset;
logic pe_6_13_done;
logic [31:0] top_6_13_in;
logic top_6_13_write_en;
logic top_6_13_clk;
logic top_6_13_reset;
logic [31:0] top_6_13_out;
logic top_6_13_done;
logic [31:0] left_6_13_in;
logic left_6_13_write_en;
logic left_6_13_clk;
logic left_6_13_reset;
logic [31:0] left_6_13_out;
logic left_6_13_done;
logic [31:0] pe_6_14_top;
logic [31:0] pe_6_14_left;
logic pe_6_14_mul_ready;
logic [31:0] pe_6_14_out;
logic pe_6_14_go;
logic pe_6_14_clk;
logic pe_6_14_reset;
logic pe_6_14_done;
logic [31:0] top_6_14_in;
logic top_6_14_write_en;
logic top_6_14_clk;
logic top_6_14_reset;
logic [31:0] top_6_14_out;
logic top_6_14_done;
logic [31:0] left_6_14_in;
logic left_6_14_write_en;
logic left_6_14_clk;
logic left_6_14_reset;
logic [31:0] left_6_14_out;
logic left_6_14_done;
logic [31:0] pe_6_15_top;
logic [31:0] pe_6_15_left;
logic pe_6_15_mul_ready;
logic [31:0] pe_6_15_out;
logic pe_6_15_go;
logic pe_6_15_clk;
logic pe_6_15_reset;
logic pe_6_15_done;
logic [31:0] top_6_15_in;
logic top_6_15_write_en;
logic top_6_15_clk;
logic top_6_15_reset;
logic [31:0] top_6_15_out;
logic top_6_15_done;
logic [31:0] left_6_15_in;
logic left_6_15_write_en;
logic left_6_15_clk;
logic left_6_15_reset;
logic [31:0] left_6_15_out;
logic left_6_15_done;
logic [31:0] pe_7_0_top;
logic [31:0] pe_7_0_left;
logic pe_7_0_mul_ready;
logic [31:0] pe_7_0_out;
logic pe_7_0_go;
logic pe_7_0_clk;
logic pe_7_0_reset;
logic pe_7_0_done;
logic [31:0] top_7_0_in;
logic top_7_0_write_en;
logic top_7_0_clk;
logic top_7_0_reset;
logic [31:0] top_7_0_out;
logic top_7_0_done;
logic [31:0] left_7_0_in;
logic left_7_0_write_en;
logic left_7_0_clk;
logic left_7_0_reset;
logic [31:0] left_7_0_out;
logic left_7_0_done;
logic [31:0] pe_7_1_top;
logic [31:0] pe_7_1_left;
logic pe_7_1_mul_ready;
logic [31:0] pe_7_1_out;
logic pe_7_1_go;
logic pe_7_1_clk;
logic pe_7_1_reset;
logic pe_7_1_done;
logic [31:0] top_7_1_in;
logic top_7_1_write_en;
logic top_7_1_clk;
logic top_7_1_reset;
logic [31:0] top_7_1_out;
logic top_7_1_done;
logic [31:0] left_7_1_in;
logic left_7_1_write_en;
logic left_7_1_clk;
logic left_7_1_reset;
logic [31:0] left_7_1_out;
logic left_7_1_done;
logic [31:0] pe_7_2_top;
logic [31:0] pe_7_2_left;
logic pe_7_2_mul_ready;
logic [31:0] pe_7_2_out;
logic pe_7_2_go;
logic pe_7_2_clk;
logic pe_7_2_reset;
logic pe_7_2_done;
logic [31:0] top_7_2_in;
logic top_7_2_write_en;
logic top_7_2_clk;
logic top_7_2_reset;
logic [31:0] top_7_2_out;
logic top_7_2_done;
logic [31:0] left_7_2_in;
logic left_7_2_write_en;
logic left_7_2_clk;
logic left_7_2_reset;
logic [31:0] left_7_2_out;
logic left_7_2_done;
logic [31:0] pe_7_3_top;
logic [31:0] pe_7_3_left;
logic pe_7_3_mul_ready;
logic [31:0] pe_7_3_out;
logic pe_7_3_go;
logic pe_7_3_clk;
logic pe_7_3_reset;
logic pe_7_3_done;
logic [31:0] top_7_3_in;
logic top_7_3_write_en;
logic top_7_3_clk;
logic top_7_3_reset;
logic [31:0] top_7_3_out;
logic top_7_3_done;
logic [31:0] left_7_3_in;
logic left_7_3_write_en;
logic left_7_3_clk;
logic left_7_3_reset;
logic [31:0] left_7_3_out;
logic left_7_3_done;
logic [31:0] pe_7_4_top;
logic [31:0] pe_7_4_left;
logic pe_7_4_mul_ready;
logic [31:0] pe_7_4_out;
logic pe_7_4_go;
logic pe_7_4_clk;
logic pe_7_4_reset;
logic pe_7_4_done;
logic [31:0] top_7_4_in;
logic top_7_4_write_en;
logic top_7_4_clk;
logic top_7_4_reset;
logic [31:0] top_7_4_out;
logic top_7_4_done;
logic [31:0] left_7_4_in;
logic left_7_4_write_en;
logic left_7_4_clk;
logic left_7_4_reset;
logic [31:0] left_7_4_out;
logic left_7_4_done;
logic [31:0] pe_7_5_top;
logic [31:0] pe_7_5_left;
logic pe_7_5_mul_ready;
logic [31:0] pe_7_5_out;
logic pe_7_5_go;
logic pe_7_5_clk;
logic pe_7_5_reset;
logic pe_7_5_done;
logic [31:0] top_7_5_in;
logic top_7_5_write_en;
logic top_7_5_clk;
logic top_7_5_reset;
logic [31:0] top_7_5_out;
logic top_7_5_done;
logic [31:0] left_7_5_in;
logic left_7_5_write_en;
logic left_7_5_clk;
logic left_7_5_reset;
logic [31:0] left_7_5_out;
logic left_7_5_done;
logic [31:0] pe_7_6_top;
logic [31:0] pe_7_6_left;
logic pe_7_6_mul_ready;
logic [31:0] pe_7_6_out;
logic pe_7_6_go;
logic pe_7_6_clk;
logic pe_7_6_reset;
logic pe_7_6_done;
logic [31:0] top_7_6_in;
logic top_7_6_write_en;
logic top_7_6_clk;
logic top_7_6_reset;
logic [31:0] top_7_6_out;
logic top_7_6_done;
logic [31:0] left_7_6_in;
logic left_7_6_write_en;
logic left_7_6_clk;
logic left_7_6_reset;
logic [31:0] left_7_6_out;
logic left_7_6_done;
logic [31:0] pe_7_7_top;
logic [31:0] pe_7_7_left;
logic pe_7_7_mul_ready;
logic [31:0] pe_7_7_out;
logic pe_7_7_go;
logic pe_7_7_clk;
logic pe_7_7_reset;
logic pe_7_7_done;
logic [31:0] top_7_7_in;
logic top_7_7_write_en;
logic top_7_7_clk;
logic top_7_7_reset;
logic [31:0] top_7_7_out;
logic top_7_7_done;
logic [31:0] left_7_7_in;
logic left_7_7_write_en;
logic left_7_7_clk;
logic left_7_7_reset;
logic [31:0] left_7_7_out;
logic left_7_7_done;
logic [31:0] pe_7_8_top;
logic [31:0] pe_7_8_left;
logic pe_7_8_mul_ready;
logic [31:0] pe_7_8_out;
logic pe_7_8_go;
logic pe_7_8_clk;
logic pe_7_8_reset;
logic pe_7_8_done;
logic [31:0] top_7_8_in;
logic top_7_8_write_en;
logic top_7_8_clk;
logic top_7_8_reset;
logic [31:0] top_7_8_out;
logic top_7_8_done;
logic [31:0] left_7_8_in;
logic left_7_8_write_en;
logic left_7_8_clk;
logic left_7_8_reset;
logic [31:0] left_7_8_out;
logic left_7_8_done;
logic [31:0] pe_7_9_top;
logic [31:0] pe_7_9_left;
logic pe_7_9_mul_ready;
logic [31:0] pe_7_9_out;
logic pe_7_9_go;
logic pe_7_9_clk;
logic pe_7_9_reset;
logic pe_7_9_done;
logic [31:0] top_7_9_in;
logic top_7_9_write_en;
logic top_7_9_clk;
logic top_7_9_reset;
logic [31:0] top_7_9_out;
logic top_7_9_done;
logic [31:0] left_7_9_in;
logic left_7_9_write_en;
logic left_7_9_clk;
logic left_7_9_reset;
logic [31:0] left_7_9_out;
logic left_7_9_done;
logic [31:0] pe_7_10_top;
logic [31:0] pe_7_10_left;
logic pe_7_10_mul_ready;
logic [31:0] pe_7_10_out;
logic pe_7_10_go;
logic pe_7_10_clk;
logic pe_7_10_reset;
logic pe_7_10_done;
logic [31:0] top_7_10_in;
logic top_7_10_write_en;
logic top_7_10_clk;
logic top_7_10_reset;
logic [31:0] top_7_10_out;
logic top_7_10_done;
logic [31:0] left_7_10_in;
logic left_7_10_write_en;
logic left_7_10_clk;
logic left_7_10_reset;
logic [31:0] left_7_10_out;
logic left_7_10_done;
logic [31:0] pe_7_11_top;
logic [31:0] pe_7_11_left;
logic pe_7_11_mul_ready;
logic [31:0] pe_7_11_out;
logic pe_7_11_go;
logic pe_7_11_clk;
logic pe_7_11_reset;
logic pe_7_11_done;
logic [31:0] top_7_11_in;
logic top_7_11_write_en;
logic top_7_11_clk;
logic top_7_11_reset;
logic [31:0] top_7_11_out;
logic top_7_11_done;
logic [31:0] left_7_11_in;
logic left_7_11_write_en;
logic left_7_11_clk;
logic left_7_11_reset;
logic [31:0] left_7_11_out;
logic left_7_11_done;
logic [31:0] pe_7_12_top;
logic [31:0] pe_7_12_left;
logic pe_7_12_mul_ready;
logic [31:0] pe_7_12_out;
logic pe_7_12_go;
logic pe_7_12_clk;
logic pe_7_12_reset;
logic pe_7_12_done;
logic [31:0] top_7_12_in;
logic top_7_12_write_en;
logic top_7_12_clk;
logic top_7_12_reset;
logic [31:0] top_7_12_out;
logic top_7_12_done;
logic [31:0] left_7_12_in;
logic left_7_12_write_en;
logic left_7_12_clk;
logic left_7_12_reset;
logic [31:0] left_7_12_out;
logic left_7_12_done;
logic [31:0] pe_7_13_top;
logic [31:0] pe_7_13_left;
logic pe_7_13_mul_ready;
logic [31:0] pe_7_13_out;
logic pe_7_13_go;
logic pe_7_13_clk;
logic pe_7_13_reset;
logic pe_7_13_done;
logic [31:0] top_7_13_in;
logic top_7_13_write_en;
logic top_7_13_clk;
logic top_7_13_reset;
logic [31:0] top_7_13_out;
logic top_7_13_done;
logic [31:0] left_7_13_in;
logic left_7_13_write_en;
logic left_7_13_clk;
logic left_7_13_reset;
logic [31:0] left_7_13_out;
logic left_7_13_done;
logic [31:0] pe_7_14_top;
logic [31:0] pe_7_14_left;
logic pe_7_14_mul_ready;
logic [31:0] pe_7_14_out;
logic pe_7_14_go;
logic pe_7_14_clk;
logic pe_7_14_reset;
logic pe_7_14_done;
logic [31:0] top_7_14_in;
logic top_7_14_write_en;
logic top_7_14_clk;
logic top_7_14_reset;
logic [31:0] top_7_14_out;
logic top_7_14_done;
logic [31:0] left_7_14_in;
logic left_7_14_write_en;
logic left_7_14_clk;
logic left_7_14_reset;
logic [31:0] left_7_14_out;
logic left_7_14_done;
logic [31:0] pe_7_15_top;
logic [31:0] pe_7_15_left;
logic pe_7_15_mul_ready;
logic [31:0] pe_7_15_out;
logic pe_7_15_go;
logic pe_7_15_clk;
logic pe_7_15_reset;
logic pe_7_15_done;
logic [31:0] top_7_15_in;
logic top_7_15_write_en;
logic top_7_15_clk;
logic top_7_15_reset;
logic [31:0] top_7_15_out;
logic top_7_15_done;
logic [31:0] left_7_15_in;
logic left_7_15_write_en;
logic left_7_15_clk;
logic left_7_15_reset;
logic [31:0] left_7_15_out;
logic left_7_15_done;
logic [31:0] pe_8_0_top;
logic [31:0] pe_8_0_left;
logic pe_8_0_mul_ready;
logic [31:0] pe_8_0_out;
logic pe_8_0_go;
logic pe_8_0_clk;
logic pe_8_0_reset;
logic pe_8_0_done;
logic [31:0] top_8_0_in;
logic top_8_0_write_en;
logic top_8_0_clk;
logic top_8_0_reset;
logic [31:0] top_8_0_out;
logic top_8_0_done;
logic [31:0] left_8_0_in;
logic left_8_0_write_en;
logic left_8_0_clk;
logic left_8_0_reset;
logic [31:0] left_8_0_out;
logic left_8_0_done;
logic [31:0] pe_8_1_top;
logic [31:0] pe_8_1_left;
logic pe_8_1_mul_ready;
logic [31:0] pe_8_1_out;
logic pe_8_1_go;
logic pe_8_1_clk;
logic pe_8_1_reset;
logic pe_8_1_done;
logic [31:0] top_8_1_in;
logic top_8_1_write_en;
logic top_8_1_clk;
logic top_8_1_reset;
logic [31:0] top_8_1_out;
logic top_8_1_done;
logic [31:0] left_8_1_in;
logic left_8_1_write_en;
logic left_8_1_clk;
logic left_8_1_reset;
logic [31:0] left_8_1_out;
logic left_8_1_done;
logic [31:0] pe_8_2_top;
logic [31:0] pe_8_2_left;
logic pe_8_2_mul_ready;
logic [31:0] pe_8_2_out;
logic pe_8_2_go;
logic pe_8_2_clk;
logic pe_8_2_reset;
logic pe_8_2_done;
logic [31:0] top_8_2_in;
logic top_8_2_write_en;
logic top_8_2_clk;
logic top_8_2_reset;
logic [31:0] top_8_2_out;
logic top_8_2_done;
logic [31:0] left_8_2_in;
logic left_8_2_write_en;
logic left_8_2_clk;
logic left_8_2_reset;
logic [31:0] left_8_2_out;
logic left_8_2_done;
logic [31:0] pe_8_3_top;
logic [31:0] pe_8_3_left;
logic pe_8_3_mul_ready;
logic [31:0] pe_8_3_out;
logic pe_8_3_go;
logic pe_8_3_clk;
logic pe_8_3_reset;
logic pe_8_3_done;
logic [31:0] top_8_3_in;
logic top_8_3_write_en;
logic top_8_3_clk;
logic top_8_3_reset;
logic [31:0] top_8_3_out;
logic top_8_3_done;
logic [31:0] left_8_3_in;
logic left_8_3_write_en;
logic left_8_3_clk;
logic left_8_3_reset;
logic [31:0] left_8_3_out;
logic left_8_3_done;
logic [31:0] pe_8_4_top;
logic [31:0] pe_8_4_left;
logic pe_8_4_mul_ready;
logic [31:0] pe_8_4_out;
logic pe_8_4_go;
logic pe_8_4_clk;
logic pe_8_4_reset;
logic pe_8_4_done;
logic [31:0] top_8_4_in;
logic top_8_4_write_en;
logic top_8_4_clk;
logic top_8_4_reset;
logic [31:0] top_8_4_out;
logic top_8_4_done;
logic [31:0] left_8_4_in;
logic left_8_4_write_en;
logic left_8_4_clk;
logic left_8_4_reset;
logic [31:0] left_8_4_out;
logic left_8_4_done;
logic [31:0] pe_8_5_top;
logic [31:0] pe_8_5_left;
logic pe_8_5_mul_ready;
logic [31:0] pe_8_5_out;
logic pe_8_5_go;
logic pe_8_5_clk;
logic pe_8_5_reset;
logic pe_8_5_done;
logic [31:0] top_8_5_in;
logic top_8_5_write_en;
logic top_8_5_clk;
logic top_8_5_reset;
logic [31:0] top_8_5_out;
logic top_8_5_done;
logic [31:0] left_8_5_in;
logic left_8_5_write_en;
logic left_8_5_clk;
logic left_8_5_reset;
logic [31:0] left_8_5_out;
logic left_8_5_done;
logic [31:0] pe_8_6_top;
logic [31:0] pe_8_6_left;
logic pe_8_6_mul_ready;
logic [31:0] pe_8_6_out;
logic pe_8_6_go;
logic pe_8_6_clk;
logic pe_8_6_reset;
logic pe_8_6_done;
logic [31:0] top_8_6_in;
logic top_8_6_write_en;
logic top_8_6_clk;
logic top_8_6_reset;
logic [31:0] top_8_6_out;
logic top_8_6_done;
logic [31:0] left_8_6_in;
logic left_8_6_write_en;
logic left_8_6_clk;
logic left_8_6_reset;
logic [31:0] left_8_6_out;
logic left_8_6_done;
logic [31:0] pe_8_7_top;
logic [31:0] pe_8_7_left;
logic pe_8_7_mul_ready;
logic [31:0] pe_8_7_out;
logic pe_8_7_go;
logic pe_8_7_clk;
logic pe_8_7_reset;
logic pe_8_7_done;
logic [31:0] top_8_7_in;
logic top_8_7_write_en;
logic top_8_7_clk;
logic top_8_7_reset;
logic [31:0] top_8_7_out;
logic top_8_7_done;
logic [31:0] left_8_7_in;
logic left_8_7_write_en;
logic left_8_7_clk;
logic left_8_7_reset;
logic [31:0] left_8_7_out;
logic left_8_7_done;
logic [31:0] pe_8_8_top;
logic [31:0] pe_8_8_left;
logic pe_8_8_mul_ready;
logic [31:0] pe_8_8_out;
logic pe_8_8_go;
logic pe_8_8_clk;
logic pe_8_8_reset;
logic pe_8_8_done;
logic [31:0] top_8_8_in;
logic top_8_8_write_en;
logic top_8_8_clk;
logic top_8_8_reset;
logic [31:0] top_8_8_out;
logic top_8_8_done;
logic [31:0] left_8_8_in;
logic left_8_8_write_en;
logic left_8_8_clk;
logic left_8_8_reset;
logic [31:0] left_8_8_out;
logic left_8_8_done;
logic [31:0] pe_8_9_top;
logic [31:0] pe_8_9_left;
logic pe_8_9_mul_ready;
logic [31:0] pe_8_9_out;
logic pe_8_9_go;
logic pe_8_9_clk;
logic pe_8_9_reset;
logic pe_8_9_done;
logic [31:0] top_8_9_in;
logic top_8_9_write_en;
logic top_8_9_clk;
logic top_8_9_reset;
logic [31:0] top_8_9_out;
logic top_8_9_done;
logic [31:0] left_8_9_in;
logic left_8_9_write_en;
logic left_8_9_clk;
logic left_8_9_reset;
logic [31:0] left_8_9_out;
logic left_8_9_done;
logic [31:0] pe_8_10_top;
logic [31:0] pe_8_10_left;
logic pe_8_10_mul_ready;
logic [31:0] pe_8_10_out;
logic pe_8_10_go;
logic pe_8_10_clk;
logic pe_8_10_reset;
logic pe_8_10_done;
logic [31:0] top_8_10_in;
logic top_8_10_write_en;
logic top_8_10_clk;
logic top_8_10_reset;
logic [31:0] top_8_10_out;
logic top_8_10_done;
logic [31:0] left_8_10_in;
logic left_8_10_write_en;
logic left_8_10_clk;
logic left_8_10_reset;
logic [31:0] left_8_10_out;
logic left_8_10_done;
logic [31:0] pe_8_11_top;
logic [31:0] pe_8_11_left;
logic pe_8_11_mul_ready;
logic [31:0] pe_8_11_out;
logic pe_8_11_go;
logic pe_8_11_clk;
logic pe_8_11_reset;
logic pe_8_11_done;
logic [31:0] top_8_11_in;
logic top_8_11_write_en;
logic top_8_11_clk;
logic top_8_11_reset;
logic [31:0] top_8_11_out;
logic top_8_11_done;
logic [31:0] left_8_11_in;
logic left_8_11_write_en;
logic left_8_11_clk;
logic left_8_11_reset;
logic [31:0] left_8_11_out;
logic left_8_11_done;
logic [31:0] pe_8_12_top;
logic [31:0] pe_8_12_left;
logic pe_8_12_mul_ready;
logic [31:0] pe_8_12_out;
logic pe_8_12_go;
logic pe_8_12_clk;
logic pe_8_12_reset;
logic pe_8_12_done;
logic [31:0] top_8_12_in;
logic top_8_12_write_en;
logic top_8_12_clk;
logic top_8_12_reset;
logic [31:0] top_8_12_out;
logic top_8_12_done;
logic [31:0] left_8_12_in;
logic left_8_12_write_en;
logic left_8_12_clk;
logic left_8_12_reset;
logic [31:0] left_8_12_out;
logic left_8_12_done;
logic [31:0] pe_8_13_top;
logic [31:0] pe_8_13_left;
logic pe_8_13_mul_ready;
logic [31:0] pe_8_13_out;
logic pe_8_13_go;
logic pe_8_13_clk;
logic pe_8_13_reset;
logic pe_8_13_done;
logic [31:0] top_8_13_in;
logic top_8_13_write_en;
logic top_8_13_clk;
logic top_8_13_reset;
logic [31:0] top_8_13_out;
logic top_8_13_done;
logic [31:0] left_8_13_in;
logic left_8_13_write_en;
logic left_8_13_clk;
logic left_8_13_reset;
logic [31:0] left_8_13_out;
logic left_8_13_done;
logic [31:0] pe_8_14_top;
logic [31:0] pe_8_14_left;
logic pe_8_14_mul_ready;
logic [31:0] pe_8_14_out;
logic pe_8_14_go;
logic pe_8_14_clk;
logic pe_8_14_reset;
logic pe_8_14_done;
logic [31:0] top_8_14_in;
logic top_8_14_write_en;
logic top_8_14_clk;
logic top_8_14_reset;
logic [31:0] top_8_14_out;
logic top_8_14_done;
logic [31:0] left_8_14_in;
logic left_8_14_write_en;
logic left_8_14_clk;
logic left_8_14_reset;
logic [31:0] left_8_14_out;
logic left_8_14_done;
logic [31:0] pe_8_15_top;
logic [31:0] pe_8_15_left;
logic pe_8_15_mul_ready;
logic [31:0] pe_8_15_out;
logic pe_8_15_go;
logic pe_8_15_clk;
logic pe_8_15_reset;
logic pe_8_15_done;
logic [31:0] top_8_15_in;
logic top_8_15_write_en;
logic top_8_15_clk;
logic top_8_15_reset;
logic [31:0] top_8_15_out;
logic top_8_15_done;
logic [31:0] left_8_15_in;
logic left_8_15_write_en;
logic left_8_15_clk;
logic left_8_15_reset;
logic [31:0] left_8_15_out;
logic left_8_15_done;
logic [31:0] pe_9_0_top;
logic [31:0] pe_9_0_left;
logic pe_9_0_mul_ready;
logic [31:0] pe_9_0_out;
logic pe_9_0_go;
logic pe_9_0_clk;
logic pe_9_0_reset;
logic pe_9_0_done;
logic [31:0] top_9_0_in;
logic top_9_0_write_en;
logic top_9_0_clk;
logic top_9_0_reset;
logic [31:0] top_9_0_out;
logic top_9_0_done;
logic [31:0] left_9_0_in;
logic left_9_0_write_en;
logic left_9_0_clk;
logic left_9_0_reset;
logic [31:0] left_9_0_out;
logic left_9_0_done;
logic [31:0] pe_9_1_top;
logic [31:0] pe_9_1_left;
logic pe_9_1_mul_ready;
logic [31:0] pe_9_1_out;
logic pe_9_1_go;
logic pe_9_1_clk;
logic pe_9_1_reset;
logic pe_9_1_done;
logic [31:0] top_9_1_in;
logic top_9_1_write_en;
logic top_9_1_clk;
logic top_9_1_reset;
logic [31:0] top_9_1_out;
logic top_9_1_done;
logic [31:0] left_9_1_in;
logic left_9_1_write_en;
logic left_9_1_clk;
logic left_9_1_reset;
logic [31:0] left_9_1_out;
logic left_9_1_done;
logic [31:0] pe_9_2_top;
logic [31:0] pe_9_2_left;
logic pe_9_2_mul_ready;
logic [31:0] pe_9_2_out;
logic pe_9_2_go;
logic pe_9_2_clk;
logic pe_9_2_reset;
logic pe_9_2_done;
logic [31:0] top_9_2_in;
logic top_9_2_write_en;
logic top_9_2_clk;
logic top_9_2_reset;
logic [31:0] top_9_2_out;
logic top_9_2_done;
logic [31:0] left_9_2_in;
logic left_9_2_write_en;
logic left_9_2_clk;
logic left_9_2_reset;
logic [31:0] left_9_2_out;
logic left_9_2_done;
logic [31:0] pe_9_3_top;
logic [31:0] pe_9_3_left;
logic pe_9_3_mul_ready;
logic [31:0] pe_9_3_out;
logic pe_9_3_go;
logic pe_9_3_clk;
logic pe_9_3_reset;
logic pe_9_3_done;
logic [31:0] top_9_3_in;
logic top_9_3_write_en;
logic top_9_3_clk;
logic top_9_3_reset;
logic [31:0] top_9_3_out;
logic top_9_3_done;
logic [31:0] left_9_3_in;
logic left_9_3_write_en;
logic left_9_3_clk;
logic left_9_3_reset;
logic [31:0] left_9_3_out;
logic left_9_3_done;
logic [31:0] pe_9_4_top;
logic [31:0] pe_9_4_left;
logic pe_9_4_mul_ready;
logic [31:0] pe_9_4_out;
logic pe_9_4_go;
logic pe_9_4_clk;
logic pe_9_4_reset;
logic pe_9_4_done;
logic [31:0] top_9_4_in;
logic top_9_4_write_en;
logic top_9_4_clk;
logic top_9_4_reset;
logic [31:0] top_9_4_out;
logic top_9_4_done;
logic [31:0] left_9_4_in;
logic left_9_4_write_en;
logic left_9_4_clk;
logic left_9_4_reset;
logic [31:0] left_9_4_out;
logic left_9_4_done;
logic [31:0] pe_9_5_top;
logic [31:0] pe_9_5_left;
logic pe_9_5_mul_ready;
logic [31:0] pe_9_5_out;
logic pe_9_5_go;
logic pe_9_5_clk;
logic pe_9_5_reset;
logic pe_9_5_done;
logic [31:0] top_9_5_in;
logic top_9_5_write_en;
logic top_9_5_clk;
logic top_9_5_reset;
logic [31:0] top_9_5_out;
logic top_9_5_done;
logic [31:0] left_9_5_in;
logic left_9_5_write_en;
logic left_9_5_clk;
logic left_9_5_reset;
logic [31:0] left_9_5_out;
logic left_9_5_done;
logic [31:0] pe_9_6_top;
logic [31:0] pe_9_6_left;
logic pe_9_6_mul_ready;
logic [31:0] pe_9_6_out;
logic pe_9_6_go;
logic pe_9_6_clk;
logic pe_9_6_reset;
logic pe_9_6_done;
logic [31:0] top_9_6_in;
logic top_9_6_write_en;
logic top_9_6_clk;
logic top_9_6_reset;
logic [31:0] top_9_6_out;
logic top_9_6_done;
logic [31:0] left_9_6_in;
logic left_9_6_write_en;
logic left_9_6_clk;
logic left_9_6_reset;
logic [31:0] left_9_6_out;
logic left_9_6_done;
logic [31:0] pe_9_7_top;
logic [31:0] pe_9_7_left;
logic pe_9_7_mul_ready;
logic [31:0] pe_9_7_out;
logic pe_9_7_go;
logic pe_9_7_clk;
logic pe_9_7_reset;
logic pe_9_7_done;
logic [31:0] top_9_7_in;
logic top_9_7_write_en;
logic top_9_7_clk;
logic top_9_7_reset;
logic [31:0] top_9_7_out;
logic top_9_7_done;
logic [31:0] left_9_7_in;
logic left_9_7_write_en;
logic left_9_7_clk;
logic left_9_7_reset;
logic [31:0] left_9_7_out;
logic left_9_7_done;
logic [31:0] pe_9_8_top;
logic [31:0] pe_9_8_left;
logic pe_9_8_mul_ready;
logic [31:0] pe_9_8_out;
logic pe_9_8_go;
logic pe_9_8_clk;
logic pe_9_8_reset;
logic pe_9_8_done;
logic [31:0] top_9_8_in;
logic top_9_8_write_en;
logic top_9_8_clk;
logic top_9_8_reset;
logic [31:0] top_9_8_out;
logic top_9_8_done;
logic [31:0] left_9_8_in;
logic left_9_8_write_en;
logic left_9_8_clk;
logic left_9_8_reset;
logic [31:0] left_9_8_out;
logic left_9_8_done;
logic [31:0] pe_9_9_top;
logic [31:0] pe_9_9_left;
logic pe_9_9_mul_ready;
logic [31:0] pe_9_9_out;
logic pe_9_9_go;
logic pe_9_9_clk;
logic pe_9_9_reset;
logic pe_9_9_done;
logic [31:0] top_9_9_in;
logic top_9_9_write_en;
logic top_9_9_clk;
logic top_9_9_reset;
logic [31:0] top_9_9_out;
logic top_9_9_done;
logic [31:0] left_9_9_in;
logic left_9_9_write_en;
logic left_9_9_clk;
logic left_9_9_reset;
logic [31:0] left_9_9_out;
logic left_9_9_done;
logic [31:0] pe_9_10_top;
logic [31:0] pe_9_10_left;
logic pe_9_10_mul_ready;
logic [31:0] pe_9_10_out;
logic pe_9_10_go;
logic pe_9_10_clk;
logic pe_9_10_reset;
logic pe_9_10_done;
logic [31:0] top_9_10_in;
logic top_9_10_write_en;
logic top_9_10_clk;
logic top_9_10_reset;
logic [31:0] top_9_10_out;
logic top_9_10_done;
logic [31:0] left_9_10_in;
logic left_9_10_write_en;
logic left_9_10_clk;
logic left_9_10_reset;
logic [31:0] left_9_10_out;
logic left_9_10_done;
logic [31:0] pe_9_11_top;
logic [31:0] pe_9_11_left;
logic pe_9_11_mul_ready;
logic [31:0] pe_9_11_out;
logic pe_9_11_go;
logic pe_9_11_clk;
logic pe_9_11_reset;
logic pe_9_11_done;
logic [31:0] top_9_11_in;
logic top_9_11_write_en;
logic top_9_11_clk;
logic top_9_11_reset;
logic [31:0] top_9_11_out;
logic top_9_11_done;
logic [31:0] left_9_11_in;
logic left_9_11_write_en;
logic left_9_11_clk;
logic left_9_11_reset;
logic [31:0] left_9_11_out;
logic left_9_11_done;
logic [31:0] pe_9_12_top;
logic [31:0] pe_9_12_left;
logic pe_9_12_mul_ready;
logic [31:0] pe_9_12_out;
logic pe_9_12_go;
logic pe_9_12_clk;
logic pe_9_12_reset;
logic pe_9_12_done;
logic [31:0] top_9_12_in;
logic top_9_12_write_en;
logic top_9_12_clk;
logic top_9_12_reset;
logic [31:0] top_9_12_out;
logic top_9_12_done;
logic [31:0] left_9_12_in;
logic left_9_12_write_en;
logic left_9_12_clk;
logic left_9_12_reset;
logic [31:0] left_9_12_out;
logic left_9_12_done;
logic [31:0] pe_9_13_top;
logic [31:0] pe_9_13_left;
logic pe_9_13_mul_ready;
logic [31:0] pe_9_13_out;
logic pe_9_13_go;
logic pe_9_13_clk;
logic pe_9_13_reset;
logic pe_9_13_done;
logic [31:0] top_9_13_in;
logic top_9_13_write_en;
logic top_9_13_clk;
logic top_9_13_reset;
logic [31:0] top_9_13_out;
logic top_9_13_done;
logic [31:0] left_9_13_in;
logic left_9_13_write_en;
logic left_9_13_clk;
logic left_9_13_reset;
logic [31:0] left_9_13_out;
logic left_9_13_done;
logic [31:0] pe_9_14_top;
logic [31:0] pe_9_14_left;
logic pe_9_14_mul_ready;
logic [31:0] pe_9_14_out;
logic pe_9_14_go;
logic pe_9_14_clk;
logic pe_9_14_reset;
logic pe_9_14_done;
logic [31:0] top_9_14_in;
logic top_9_14_write_en;
logic top_9_14_clk;
logic top_9_14_reset;
logic [31:0] top_9_14_out;
logic top_9_14_done;
logic [31:0] left_9_14_in;
logic left_9_14_write_en;
logic left_9_14_clk;
logic left_9_14_reset;
logic [31:0] left_9_14_out;
logic left_9_14_done;
logic [31:0] pe_9_15_top;
logic [31:0] pe_9_15_left;
logic pe_9_15_mul_ready;
logic [31:0] pe_9_15_out;
logic pe_9_15_go;
logic pe_9_15_clk;
logic pe_9_15_reset;
logic pe_9_15_done;
logic [31:0] top_9_15_in;
logic top_9_15_write_en;
logic top_9_15_clk;
logic top_9_15_reset;
logic [31:0] top_9_15_out;
logic top_9_15_done;
logic [31:0] left_9_15_in;
logic left_9_15_write_en;
logic left_9_15_clk;
logic left_9_15_reset;
logic [31:0] left_9_15_out;
logic left_9_15_done;
logic [31:0] pe_10_0_top;
logic [31:0] pe_10_0_left;
logic pe_10_0_mul_ready;
logic [31:0] pe_10_0_out;
logic pe_10_0_go;
logic pe_10_0_clk;
logic pe_10_0_reset;
logic pe_10_0_done;
logic [31:0] top_10_0_in;
logic top_10_0_write_en;
logic top_10_0_clk;
logic top_10_0_reset;
logic [31:0] top_10_0_out;
logic top_10_0_done;
logic [31:0] left_10_0_in;
logic left_10_0_write_en;
logic left_10_0_clk;
logic left_10_0_reset;
logic [31:0] left_10_0_out;
logic left_10_0_done;
logic [31:0] pe_10_1_top;
logic [31:0] pe_10_1_left;
logic pe_10_1_mul_ready;
logic [31:0] pe_10_1_out;
logic pe_10_1_go;
logic pe_10_1_clk;
logic pe_10_1_reset;
logic pe_10_1_done;
logic [31:0] top_10_1_in;
logic top_10_1_write_en;
logic top_10_1_clk;
logic top_10_1_reset;
logic [31:0] top_10_1_out;
logic top_10_1_done;
logic [31:0] left_10_1_in;
logic left_10_1_write_en;
logic left_10_1_clk;
logic left_10_1_reset;
logic [31:0] left_10_1_out;
logic left_10_1_done;
logic [31:0] pe_10_2_top;
logic [31:0] pe_10_2_left;
logic pe_10_2_mul_ready;
logic [31:0] pe_10_2_out;
logic pe_10_2_go;
logic pe_10_2_clk;
logic pe_10_2_reset;
logic pe_10_2_done;
logic [31:0] top_10_2_in;
logic top_10_2_write_en;
logic top_10_2_clk;
logic top_10_2_reset;
logic [31:0] top_10_2_out;
logic top_10_2_done;
logic [31:0] left_10_2_in;
logic left_10_2_write_en;
logic left_10_2_clk;
logic left_10_2_reset;
logic [31:0] left_10_2_out;
logic left_10_2_done;
logic [31:0] pe_10_3_top;
logic [31:0] pe_10_3_left;
logic pe_10_3_mul_ready;
logic [31:0] pe_10_3_out;
logic pe_10_3_go;
logic pe_10_3_clk;
logic pe_10_3_reset;
logic pe_10_3_done;
logic [31:0] top_10_3_in;
logic top_10_3_write_en;
logic top_10_3_clk;
logic top_10_3_reset;
logic [31:0] top_10_3_out;
logic top_10_3_done;
logic [31:0] left_10_3_in;
logic left_10_3_write_en;
logic left_10_3_clk;
logic left_10_3_reset;
logic [31:0] left_10_3_out;
logic left_10_3_done;
logic [31:0] pe_10_4_top;
logic [31:0] pe_10_4_left;
logic pe_10_4_mul_ready;
logic [31:0] pe_10_4_out;
logic pe_10_4_go;
logic pe_10_4_clk;
logic pe_10_4_reset;
logic pe_10_4_done;
logic [31:0] top_10_4_in;
logic top_10_4_write_en;
logic top_10_4_clk;
logic top_10_4_reset;
logic [31:0] top_10_4_out;
logic top_10_4_done;
logic [31:0] left_10_4_in;
logic left_10_4_write_en;
logic left_10_4_clk;
logic left_10_4_reset;
logic [31:0] left_10_4_out;
logic left_10_4_done;
logic [31:0] pe_10_5_top;
logic [31:0] pe_10_5_left;
logic pe_10_5_mul_ready;
logic [31:0] pe_10_5_out;
logic pe_10_5_go;
logic pe_10_5_clk;
logic pe_10_5_reset;
logic pe_10_5_done;
logic [31:0] top_10_5_in;
logic top_10_5_write_en;
logic top_10_5_clk;
logic top_10_5_reset;
logic [31:0] top_10_5_out;
logic top_10_5_done;
logic [31:0] left_10_5_in;
logic left_10_5_write_en;
logic left_10_5_clk;
logic left_10_5_reset;
logic [31:0] left_10_5_out;
logic left_10_5_done;
logic [31:0] pe_10_6_top;
logic [31:0] pe_10_6_left;
logic pe_10_6_mul_ready;
logic [31:0] pe_10_6_out;
logic pe_10_6_go;
logic pe_10_6_clk;
logic pe_10_6_reset;
logic pe_10_6_done;
logic [31:0] top_10_6_in;
logic top_10_6_write_en;
logic top_10_6_clk;
logic top_10_6_reset;
logic [31:0] top_10_6_out;
logic top_10_6_done;
logic [31:0] left_10_6_in;
logic left_10_6_write_en;
logic left_10_6_clk;
logic left_10_6_reset;
logic [31:0] left_10_6_out;
logic left_10_6_done;
logic [31:0] pe_10_7_top;
logic [31:0] pe_10_7_left;
logic pe_10_7_mul_ready;
logic [31:0] pe_10_7_out;
logic pe_10_7_go;
logic pe_10_7_clk;
logic pe_10_7_reset;
logic pe_10_7_done;
logic [31:0] top_10_7_in;
logic top_10_7_write_en;
logic top_10_7_clk;
logic top_10_7_reset;
logic [31:0] top_10_7_out;
logic top_10_7_done;
logic [31:0] left_10_7_in;
logic left_10_7_write_en;
logic left_10_7_clk;
logic left_10_7_reset;
logic [31:0] left_10_7_out;
logic left_10_7_done;
logic [31:0] pe_10_8_top;
logic [31:0] pe_10_8_left;
logic pe_10_8_mul_ready;
logic [31:0] pe_10_8_out;
logic pe_10_8_go;
logic pe_10_8_clk;
logic pe_10_8_reset;
logic pe_10_8_done;
logic [31:0] top_10_8_in;
logic top_10_8_write_en;
logic top_10_8_clk;
logic top_10_8_reset;
logic [31:0] top_10_8_out;
logic top_10_8_done;
logic [31:0] left_10_8_in;
logic left_10_8_write_en;
logic left_10_8_clk;
logic left_10_8_reset;
logic [31:0] left_10_8_out;
logic left_10_8_done;
logic [31:0] pe_10_9_top;
logic [31:0] pe_10_9_left;
logic pe_10_9_mul_ready;
logic [31:0] pe_10_9_out;
logic pe_10_9_go;
logic pe_10_9_clk;
logic pe_10_9_reset;
logic pe_10_9_done;
logic [31:0] top_10_9_in;
logic top_10_9_write_en;
logic top_10_9_clk;
logic top_10_9_reset;
logic [31:0] top_10_9_out;
logic top_10_9_done;
logic [31:0] left_10_9_in;
logic left_10_9_write_en;
logic left_10_9_clk;
logic left_10_9_reset;
logic [31:0] left_10_9_out;
logic left_10_9_done;
logic [31:0] pe_10_10_top;
logic [31:0] pe_10_10_left;
logic pe_10_10_mul_ready;
logic [31:0] pe_10_10_out;
logic pe_10_10_go;
logic pe_10_10_clk;
logic pe_10_10_reset;
logic pe_10_10_done;
logic [31:0] top_10_10_in;
logic top_10_10_write_en;
logic top_10_10_clk;
logic top_10_10_reset;
logic [31:0] top_10_10_out;
logic top_10_10_done;
logic [31:0] left_10_10_in;
logic left_10_10_write_en;
logic left_10_10_clk;
logic left_10_10_reset;
logic [31:0] left_10_10_out;
logic left_10_10_done;
logic [31:0] pe_10_11_top;
logic [31:0] pe_10_11_left;
logic pe_10_11_mul_ready;
logic [31:0] pe_10_11_out;
logic pe_10_11_go;
logic pe_10_11_clk;
logic pe_10_11_reset;
logic pe_10_11_done;
logic [31:0] top_10_11_in;
logic top_10_11_write_en;
logic top_10_11_clk;
logic top_10_11_reset;
logic [31:0] top_10_11_out;
logic top_10_11_done;
logic [31:0] left_10_11_in;
logic left_10_11_write_en;
logic left_10_11_clk;
logic left_10_11_reset;
logic [31:0] left_10_11_out;
logic left_10_11_done;
logic [31:0] pe_10_12_top;
logic [31:0] pe_10_12_left;
logic pe_10_12_mul_ready;
logic [31:0] pe_10_12_out;
logic pe_10_12_go;
logic pe_10_12_clk;
logic pe_10_12_reset;
logic pe_10_12_done;
logic [31:0] top_10_12_in;
logic top_10_12_write_en;
logic top_10_12_clk;
logic top_10_12_reset;
logic [31:0] top_10_12_out;
logic top_10_12_done;
logic [31:0] left_10_12_in;
logic left_10_12_write_en;
logic left_10_12_clk;
logic left_10_12_reset;
logic [31:0] left_10_12_out;
logic left_10_12_done;
logic [31:0] pe_10_13_top;
logic [31:0] pe_10_13_left;
logic pe_10_13_mul_ready;
logic [31:0] pe_10_13_out;
logic pe_10_13_go;
logic pe_10_13_clk;
logic pe_10_13_reset;
logic pe_10_13_done;
logic [31:0] top_10_13_in;
logic top_10_13_write_en;
logic top_10_13_clk;
logic top_10_13_reset;
logic [31:0] top_10_13_out;
logic top_10_13_done;
logic [31:0] left_10_13_in;
logic left_10_13_write_en;
logic left_10_13_clk;
logic left_10_13_reset;
logic [31:0] left_10_13_out;
logic left_10_13_done;
logic [31:0] pe_10_14_top;
logic [31:0] pe_10_14_left;
logic pe_10_14_mul_ready;
logic [31:0] pe_10_14_out;
logic pe_10_14_go;
logic pe_10_14_clk;
logic pe_10_14_reset;
logic pe_10_14_done;
logic [31:0] top_10_14_in;
logic top_10_14_write_en;
logic top_10_14_clk;
logic top_10_14_reset;
logic [31:0] top_10_14_out;
logic top_10_14_done;
logic [31:0] left_10_14_in;
logic left_10_14_write_en;
logic left_10_14_clk;
logic left_10_14_reset;
logic [31:0] left_10_14_out;
logic left_10_14_done;
logic [31:0] pe_10_15_top;
logic [31:0] pe_10_15_left;
logic pe_10_15_mul_ready;
logic [31:0] pe_10_15_out;
logic pe_10_15_go;
logic pe_10_15_clk;
logic pe_10_15_reset;
logic pe_10_15_done;
logic [31:0] top_10_15_in;
logic top_10_15_write_en;
logic top_10_15_clk;
logic top_10_15_reset;
logic [31:0] top_10_15_out;
logic top_10_15_done;
logic [31:0] left_10_15_in;
logic left_10_15_write_en;
logic left_10_15_clk;
logic left_10_15_reset;
logic [31:0] left_10_15_out;
logic left_10_15_done;
logic [31:0] pe_11_0_top;
logic [31:0] pe_11_0_left;
logic pe_11_0_mul_ready;
logic [31:0] pe_11_0_out;
logic pe_11_0_go;
logic pe_11_0_clk;
logic pe_11_0_reset;
logic pe_11_0_done;
logic [31:0] top_11_0_in;
logic top_11_0_write_en;
logic top_11_0_clk;
logic top_11_0_reset;
logic [31:0] top_11_0_out;
logic top_11_0_done;
logic [31:0] left_11_0_in;
logic left_11_0_write_en;
logic left_11_0_clk;
logic left_11_0_reset;
logic [31:0] left_11_0_out;
logic left_11_0_done;
logic [31:0] pe_11_1_top;
logic [31:0] pe_11_1_left;
logic pe_11_1_mul_ready;
logic [31:0] pe_11_1_out;
logic pe_11_1_go;
logic pe_11_1_clk;
logic pe_11_1_reset;
logic pe_11_1_done;
logic [31:0] top_11_1_in;
logic top_11_1_write_en;
logic top_11_1_clk;
logic top_11_1_reset;
logic [31:0] top_11_1_out;
logic top_11_1_done;
logic [31:0] left_11_1_in;
logic left_11_1_write_en;
logic left_11_1_clk;
logic left_11_1_reset;
logic [31:0] left_11_1_out;
logic left_11_1_done;
logic [31:0] pe_11_2_top;
logic [31:0] pe_11_2_left;
logic pe_11_2_mul_ready;
logic [31:0] pe_11_2_out;
logic pe_11_2_go;
logic pe_11_2_clk;
logic pe_11_2_reset;
logic pe_11_2_done;
logic [31:0] top_11_2_in;
logic top_11_2_write_en;
logic top_11_2_clk;
logic top_11_2_reset;
logic [31:0] top_11_2_out;
logic top_11_2_done;
logic [31:0] left_11_2_in;
logic left_11_2_write_en;
logic left_11_2_clk;
logic left_11_2_reset;
logic [31:0] left_11_2_out;
logic left_11_2_done;
logic [31:0] pe_11_3_top;
logic [31:0] pe_11_3_left;
logic pe_11_3_mul_ready;
logic [31:0] pe_11_3_out;
logic pe_11_3_go;
logic pe_11_3_clk;
logic pe_11_3_reset;
logic pe_11_3_done;
logic [31:0] top_11_3_in;
logic top_11_3_write_en;
logic top_11_3_clk;
logic top_11_3_reset;
logic [31:0] top_11_3_out;
logic top_11_3_done;
logic [31:0] left_11_3_in;
logic left_11_3_write_en;
logic left_11_3_clk;
logic left_11_3_reset;
logic [31:0] left_11_3_out;
logic left_11_3_done;
logic [31:0] pe_11_4_top;
logic [31:0] pe_11_4_left;
logic pe_11_4_mul_ready;
logic [31:0] pe_11_4_out;
logic pe_11_4_go;
logic pe_11_4_clk;
logic pe_11_4_reset;
logic pe_11_4_done;
logic [31:0] top_11_4_in;
logic top_11_4_write_en;
logic top_11_4_clk;
logic top_11_4_reset;
logic [31:0] top_11_4_out;
logic top_11_4_done;
logic [31:0] left_11_4_in;
logic left_11_4_write_en;
logic left_11_4_clk;
logic left_11_4_reset;
logic [31:0] left_11_4_out;
logic left_11_4_done;
logic [31:0] pe_11_5_top;
logic [31:0] pe_11_5_left;
logic pe_11_5_mul_ready;
logic [31:0] pe_11_5_out;
logic pe_11_5_go;
logic pe_11_5_clk;
logic pe_11_5_reset;
logic pe_11_5_done;
logic [31:0] top_11_5_in;
logic top_11_5_write_en;
logic top_11_5_clk;
logic top_11_5_reset;
logic [31:0] top_11_5_out;
logic top_11_5_done;
logic [31:0] left_11_5_in;
logic left_11_5_write_en;
logic left_11_5_clk;
logic left_11_5_reset;
logic [31:0] left_11_5_out;
logic left_11_5_done;
logic [31:0] pe_11_6_top;
logic [31:0] pe_11_6_left;
logic pe_11_6_mul_ready;
logic [31:0] pe_11_6_out;
logic pe_11_6_go;
logic pe_11_6_clk;
logic pe_11_6_reset;
logic pe_11_6_done;
logic [31:0] top_11_6_in;
logic top_11_6_write_en;
logic top_11_6_clk;
logic top_11_6_reset;
logic [31:0] top_11_6_out;
logic top_11_6_done;
logic [31:0] left_11_6_in;
logic left_11_6_write_en;
logic left_11_6_clk;
logic left_11_6_reset;
logic [31:0] left_11_6_out;
logic left_11_6_done;
logic [31:0] pe_11_7_top;
logic [31:0] pe_11_7_left;
logic pe_11_7_mul_ready;
logic [31:0] pe_11_7_out;
logic pe_11_7_go;
logic pe_11_7_clk;
logic pe_11_7_reset;
logic pe_11_7_done;
logic [31:0] top_11_7_in;
logic top_11_7_write_en;
logic top_11_7_clk;
logic top_11_7_reset;
logic [31:0] top_11_7_out;
logic top_11_7_done;
logic [31:0] left_11_7_in;
logic left_11_7_write_en;
logic left_11_7_clk;
logic left_11_7_reset;
logic [31:0] left_11_7_out;
logic left_11_7_done;
logic [31:0] pe_11_8_top;
logic [31:0] pe_11_8_left;
logic pe_11_8_mul_ready;
logic [31:0] pe_11_8_out;
logic pe_11_8_go;
logic pe_11_8_clk;
logic pe_11_8_reset;
logic pe_11_8_done;
logic [31:0] top_11_8_in;
logic top_11_8_write_en;
logic top_11_8_clk;
logic top_11_8_reset;
logic [31:0] top_11_8_out;
logic top_11_8_done;
logic [31:0] left_11_8_in;
logic left_11_8_write_en;
logic left_11_8_clk;
logic left_11_8_reset;
logic [31:0] left_11_8_out;
logic left_11_8_done;
logic [31:0] pe_11_9_top;
logic [31:0] pe_11_9_left;
logic pe_11_9_mul_ready;
logic [31:0] pe_11_9_out;
logic pe_11_9_go;
logic pe_11_9_clk;
logic pe_11_9_reset;
logic pe_11_9_done;
logic [31:0] top_11_9_in;
logic top_11_9_write_en;
logic top_11_9_clk;
logic top_11_9_reset;
logic [31:0] top_11_9_out;
logic top_11_9_done;
logic [31:0] left_11_9_in;
logic left_11_9_write_en;
logic left_11_9_clk;
logic left_11_9_reset;
logic [31:0] left_11_9_out;
logic left_11_9_done;
logic [31:0] pe_11_10_top;
logic [31:0] pe_11_10_left;
logic pe_11_10_mul_ready;
logic [31:0] pe_11_10_out;
logic pe_11_10_go;
logic pe_11_10_clk;
logic pe_11_10_reset;
logic pe_11_10_done;
logic [31:0] top_11_10_in;
logic top_11_10_write_en;
logic top_11_10_clk;
logic top_11_10_reset;
logic [31:0] top_11_10_out;
logic top_11_10_done;
logic [31:0] left_11_10_in;
logic left_11_10_write_en;
logic left_11_10_clk;
logic left_11_10_reset;
logic [31:0] left_11_10_out;
logic left_11_10_done;
logic [31:0] pe_11_11_top;
logic [31:0] pe_11_11_left;
logic pe_11_11_mul_ready;
logic [31:0] pe_11_11_out;
logic pe_11_11_go;
logic pe_11_11_clk;
logic pe_11_11_reset;
logic pe_11_11_done;
logic [31:0] top_11_11_in;
logic top_11_11_write_en;
logic top_11_11_clk;
logic top_11_11_reset;
logic [31:0] top_11_11_out;
logic top_11_11_done;
logic [31:0] left_11_11_in;
logic left_11_11_write_en;
logic left_11_11_clk;
logic left_11_11_reset;
logic [31:0] left_11_11_out;
logic left_11_11_done;
logic [31:0] pe_11_12_top;
logic [31:0] pe_11_12_left;
logic pe_11_12_mul_ready;
logic [31:0] pe_11_12_out;
logic pe_11_12_go;
logic pe_11_12_clk;
logic pe_11_12_reset;
logic pe_11_12_done;
logic [31:0] top_11_12_in;
logic top_11_12_write_en;
logic top_11_12_clk;
logic top_11_12_reset;
logic [31:0] top_11_12_out;
logic top_11_12_done;
logic [31:0] left_11_12_in;
logic left_11_12_write_en;
logic left_11_12_clk;
logic left_11_12_reset;
logic [31:0] left_11_12_out;
logic left_11_12_done;
logic [31:0] pe_11_13_top;
logic [31:0] pe_11_13_left;
logic pe_11_13_mul_ready;
logic [31:0] pe_11_13_out;
logic pe_11_13_go;
logic pe_11_13_clk;
logic pe_11_13_reset;
logic pe_11_13_done;
logic [31:0] top_11_13_in;
logic top_11_13_write_en;
logic top_11_13_clk;
logic top_11_13_reset;
logic [31:0] top_11_13_out;
logic top_11_13_done;
logic [31:0] left_11_13_in;
logic left_11_13_write_en;
logic left_11_13_clk;
logic left_11_13_reset;
logic [31:0] left_11_13_out;
logic left_11_13_done;
logic [31:0] pe_11_14_top;
logic [31:0] pe_11_14_left;
logic pe_11_14_mul_ready;
logic [31:0] pe_11_14_out;
logic pe_11_14_go;
logic pe_11_14_clk;
logic pe_11_14_reset;
logic pe_11_14_done;
logic [31:0] top_11_14_in;
logic top_11_14_write_en;
logic top_11_14_clk;
logic top_11_14_reset;
logic [31:0] top_11_14_out;
logic top_11_14_done;
logic [31:0] left_11_14_in;
logic left_11_14_write_en;
logic left_11_14_clk;
logic left_11_14_reset;
logic [31:0] left_11_14_out;
logic left_11_14_done;
logic [31:0] pe_11_15_top;
logic [31:0] pe_11_15_left;
logic pe_11_15_mul_ready;
logic [31:0] pe_11_15_out;
logic pe_11_15_go;
logic pe_11_15_clk;
logic pe_11_15_reset;
logic pe_11_15_done;
logic [31:0] top_11_15_in;
logic top_11_15_write_en;
logic top_11_15_clk;
logic top_11_15_reset;
logic [31:0] top_11_15_out;
logic top_11_15_done;
logic [31:0] left_11_15_in;
logic left_11_15_write_en;
logic left_11_15_clk;
logic left_11_15_reset;
logic [31:0] left_11_15_out;
logic left_11_15_done;
logic [31:0] pe_12_0_top;
logic [31:0] pe_12_0_left;
logic pe_12_0_mul_ready;
logic [31:0] pe_12_0_out;
logic pe_12_0_go;
logic pe_12_0_clk;
logic pe_12_0_reset;
logic pe_12_0_done;
logic [31:0] top_12_0_in;
logic top_12_0_write_en;
logic top_12_0_clk;
logic top_12_0_reset;
logic [31:0] top_12_0_out;
logic top_12_0_done;
logic [31:0] left_12_0_in;
logic left_12_0_write_en;
logic left_12_0_clk;
logic left_12_0_reset;
logic [31:0] left_12_0_out;
logic left_12_0_done;
logic [31:0] pe_12_1_top;
logic [31:0] pe_12_1_left;
logic pe_12_1_mul_ready;
logic [31:0] pe_12_1_out;
logic pe_12_1_go;
logic pe_12_1_clk;
logic pe_12_1_reset;
logic pe_12_1_done;
logic [31:0] top_12_1_in;
logic top_12_1_write_en;
logic top_12_1_clk;
logic top_12_1_reset;
logic [31:0] top_12_1_out;
logic top_12_1_done;
logic [31:0] left_12_1_in;
logic left_12_1_write_en;
logic left_12_1_clk;
logic left_12_1_reset;
logic [31:0] left_12_1_out;
logic left_12_1_done;
logic [31:0] pe_12_2_top;
logic [31:0] pe_12_2_left;
logic pe_12_2_mul_ready;
logic [31:0] pe_12_2_out;
logic pe_12_2_go;
logic pe_12_2_clk;
logic pe_12_2_reset;
logic pe_12_2_done;
logic [31:0] top_12_2_in;
logic top_12_2_write_en;
logic top_12_2_clk;
logic top_12_2_reset;
logic [31:0] top_12_2_out;
logic top_12_2_done;
logic [31:0] left_12_2_in;
logic left_12_2_write_en;
logic left_12_2_clk;
logic left_12_2_reset;
logic [31:0] left_12_2_out;
logic left_12_2_done;
logic [31:0] pe_12_3_top;
logic [31:0] pe_12_3_left;
logic pe_12_3_mul_ready;
logic [31:0] pe_12_3_out;
logic pe_12_3_go;
logic pe_12_3_clk;
logic pe_12_3_reset;
logic pe_12_3_done;
logic [31:0] top_12_3_in;
logic top_12_3_write_en;
logic top_12_3_clk;
logic top_12_3_reset;
logic [31:0] top_12_3_out;
logic top_12_3_done;
logic [31:0] left_12_3_in;
logic left_12_3_write_en;
logic left_12_3_clk;
logic left_12_3_reset;
logic [31:0] left_12_3_out;
logic left_12_3_done;
logic [31:0] pe_12_4_top;
logic [31:0] pe_12_4_left;
logic pe_12_4_mul_ready;
logic [31:0] pe_12_4_out;
logic pe_12_4_go;
logic pe_12_4_clk;
logic pe_12_4_reset;
logic pe_12_4_done;
logic [31:0] top_12_4_in;
logic top_12_4_write_en;
logic top_12_4_clk;
logic top_12_4_reset;
logic [31:0] top_12_4_out;
logic top_12_4_done;
logic [31:0] left_12_4_in;
logic left_12_4_write_en;
logic left_12_4_clk;
logic left_12_4_reset;
logic [31:0] left_12_4_out;
logic left_12_4_done;
logic [31:0] pe_12_5_top;
logic [31:0] pe_12_5_left;
logic pe_12_5_mul_ready;
logic [31:0] pe_12_5_out;
logic pe_12_5_go;
logic pe_12_5_clk;
logic pe_12_5_reset;
logic pe_12_5_done;
logic [31:0] top_12_5_in;
logic top_12_5_write_en;
logic top_12_5_clk;
logic top_12_5_reset;
logic [31:0] top_12_5_out;
logic top_12_5_done;
logic [31:0] left_12_5_in;
logic left_12_5_write_en;
logic left_12_5_clk;
logic left_12_5_reset;
logic [31:0] left_12_5_out;
logic left_12_5_done;
logic [31:0] pe_12_6_top;
logic [31:0] pe_12_6_left;
logic pe_12_6_mul_ready;
logic [31:0] pe_12_6_out;
logic pe_12_6_go;
logic pe_12_6_clk;
logic pe_12_6_reset;
logic pe_12_6_done;
logic [31:0] top_12_6_in;
logic top_12_6_write_en;
logic top_12_6_clk;
logic top_12_6_reset;
logic [31:0] top_12_6_out;
logic top_12_6_done;
logic [31:0] left_12_6_in;
logic left_12_6_write_en;
logic left_12_6_clk;
logic left_12_6_reset;
logic [31:0] left_12_6_out;
logic left_12_6_done;
logic [31:0] pe_12_7_top;
logic [31:0] pe_12_7_left;
logic pe_12_7_mul_ready;
logic [31:0] pe_12_7_out;
logic pe_12_7_go;
logic pe_12_7_clk;
logic pe_12_7_reset;
logic pe_12_7_done;
logic [31:0] top_12_7_in;
logic top_12_7_write_en;
logic top_12_7_clk;
logic top_12_7_reset;
logic [31:0] top_12_7_out;
logic top_12_7_done;
logic [31:0] left_12_7_in;
logic left_12_7_write_en;
logic left_12_7_clk;
logic left_12_7_reset;
logic [31:0] left_12_7_out;
logic left_12_7_done;
logic [31:0] pe_12_8_top;
logic [31:0] pe_12_8_left;
logic pe_12_8_mul_ready;
logic [31:0] pe_12_8_out;
logic pe_12_8_go;
logic pe_12_8_clk;
logic pe_12_8_reset;
logic pe_12_8_done;
logic [31:0] top_12_8_in;
logic top_12_8_write_en;
logic top_12_8_clk;
logic top_12_8_reset;
logic [31:0] top_12_8_out;
logic top_12_8_done;
logic [31:0] left_12_8_in;
logic left_12_8_write_en;
logic left_12_8_clk;
logic left_12_8_reset;
logic [31:0] left_12_8_out;
logic left_12_8_done;
logic [31:0] pe_12_9_top;
logic [31:0] pe_12_9_left;
logic pe_12_9_mul_ready;
logic [31:0] pe_12_9_out;
logic pe_12_9_go;
logic pe_12_9_clk;
logic pe_12_9_reset;
logic pe_12_9_done;
logic [31:0] top_12_9_in;
logic top_12_9_write_en;
logic top_12_9_clk;
logic top_12_9_reset;
logic [31:0] top_12_9_out;
logic top_12_9_done;
logic [31:0] left_12_9_in;
logic left_12_9_write_en;
logic left_12_9_clk;
logic left_12_9_reset;
logic [31:0] left_12_9_out;
logic left_12_9_done;
logic [31:0] pe_12_10_top;
logic [31:0] pe_12_10_left;
logic pe_12_10_mul_ready;
logic [31:0] pe_12_10_out;
logic pe_12_10_go;
logic pe_12_10_clk;
logic pe_12_10_reset;
logic pe_12_10_done;
logic [31:0] top_12_10_in;
logic top_12_10_write_en;
logic top_12_10_clk;
logic top_12_10_reset;
logic [31:0] top_12_10_out;
logic top_12_10_done;
logic [31:0] left_12_10_in;
logic left_12_10_write_en;
logic left_12_10_clk;
logic left_12_10_reset;
logic [31:0] left_12_10_out;
logic left_12_10_done;
logic [31:0] pe_12_11_top;
logic [31:0] pe_12_11_left;
logic pe_12_11_mul_ready;
logic [31:0] pe_12_11_out;
logic pe_12_11_go;
logic pe_12_11_clk;
logic pe_12_11_reset;
logic pe_12_11_done;
logic [31:0] top_12_11_in;
logic top_12_11_write_en;
logic top_12_11_clk;
logic top_12_11_reset;
logic [31:0] top_12_11_out;
logic top_12_11_done;
logic [31:0] left_12_11_in;
logic left_12_11_write_en;
logic left_12_11_clk;
logic left_12_11_reset;
logic [31:0] left_12_11_out;
logic left_12_11_done;
logic [31:0] pe_12_12_top;
logic [31:0] pe_12_12_left;
logic pe_12_12_mul_ready;
logic [31:0] pe_12_12_out;
logic pe_12_12_go;
logic pe_12_12_clk;
logic pe_12_12_reset;
logic pe_12_12_done;
logic [31:0] top_12_12_in;
logic top_12_12_write_en;
logic top_12_12_clk;
logic top_12_12_reset;
logic [31:0] top_12_12_out;
logic top_12_12_done;
logic [31:0] left_12_12_in;
logic left_12_12_write_en;
logic left_12_12_clk;
logic left_12_12_reset;
logic [31:0] left_12_12_out;
logic left_12_12_done;
logic [31:0] pe_12_13_top;
logic [31:0] pe_12_13_left;
logic pe_12_13_mul_ready;
logic [31:0] pe_12_13_out;
logic pe_12_13_go;
logic pe_12_13_clk;
logic pe_12_13_reset;
logic pe_12_13_done;
logic [31:0] top_12_13_in;
logic top_12_13_write_en;
logic top_12_13_clk;
logic top_12_13_reset;
logic [31:0] top_12_13_out;
logic top_12_13_done;
logic [31:0] left_12_13_in;
logic left_12_13_write_en;
logic left_12_13_clk;
logic left_12_13_reset;
logic [31:0] left_12_13_out;
logic left_12_13_done;
logic [31:0] pe_12_14_top;
logic [31:0] pe_12_14_left;
logic pe_12_14_mul_ready;
logic [31:0] pe_12_14_out;
logic pe_12_14_go;
logic pe_12_14_clk;
logic pe_12_14_reset;
logic pe_12_14_done;
logic [31:0] top_12_14_in;
logic top_12_14_write_en;
logic top_12_14_clk;
logic top_12_14_reset;
logic [31:0] top_12_14_out;
logic top_12_14_done;
logic [31:0] left_12_14_in;
logic left_12_14_write_en;
logic left_12_14_clk;
logic left_12_14_reset;
logic [31:0] left_12_14_out;
logic left_12_14_done;
logic [31:0] pe_12_15_top;
logic [31:0] pe_12_15_left;
logic pe_12_15_mul_ready;
logic [31:0] pe_12_15_out;
logic pe_12_15_go;
logic pe_12_15_clk;
logic pe_12_15_reset;
logic pe_12_15_done;
logic [31:0] top_12_15_in;
logic top_12_15_write_en;
logic top_12_15_clk;
logic top_12_15_reset;
logic [31:0] top_12_15_out;
logic top_12_15_done;
logic [31:0] left_12_15_in;
logic left_12_15_write_en;
logic left_12_15_clk;
logic left_12_15_reset;
logic [31:0] left_12_15_out;
logic left_12_15_done;
logic [31:0] pe_13_0_top;
logic [31:0] pe_13_0_left;
logic pe_13_0_mul_ready;
logic [31:0] pe_13_0_out;
logic pe_13_0_go;
logic pe_13_0_clk;
logic pe_13_0_reset;
logic pe_13_0_done;
logic [31:0] top_13_0_in;
logic top_13_0_write_en;
logic top_13_0_clk;
logic top_13_0_reset;
logic [31:0] top_13_0_out;
logic top_13_0_done;
logic [31:0] left_13_0_in;
logic left_13_0_write_en;
logic left_13_0_clk;
logic left_13_0_reset;
logic [31:0] left_13_0_out;
logic left_13_0_done;
logic [31:0] pe_13_1_top;
logic [31:0] pe_13_1_left;
logic pe_13_1_mul_ready;
logic [31:0] pe_13_1_out;
logic pe_13_1_go;
logic pe_13_1_clk;
logic pe_13_1_reset;
logic pe_13_1_done;
logic [31:0] top_13_1_in;
logic top_13_1_write_en;
logic top_13_1_clk;
logic top_13_1_reset;
logic [31:0] top_13_1_out;
logic top_13_1_done;
logic [31:0] left_13_1_in;
logic left_13_1_write_en;
logic left_13_1_clk;
logic left_13_1_reset;
logic [31:0] left_13_1_out;
logic left_13_1_done;
logic [31:0] pe_13_2_top;
logic [31:0] pe_13_2_left;
logic pe_13_2_mul_ready;
logic [31:0] pe_13_2_out;
logic pe_13_2_go;
logic pe_13_2_clk;
logic pe_13_2_reset;
logic pe_13_2_done;
logic [31:0] top_13_2_in;
logic top_13_2_write_en;
logic top_13_2_clk;
logic top_13_2_reset;
logic [31:0] top_13_2_out;
logic top_13_2_done;
logic [31:0] left_13_2_in;
logic left_13_2_write_en;
logic left_13_2_clk;
logic left_13_2_reset;
logic [31:0] left_13_2_out;
logic left_13_2_done;
logic [31:0] pe_13_3_top;
logic [31:0] pe_13_3_left;
logic pe_13_3_mul_ready;
logic [31:0] pe_13_3_out;
logic pe_13_3_go;
logic pe_13_3_clk;
logic pe_13_3_reset;
logic pe_13_3_done;
logic [31:0] top_13_3_in;
logic top_13_3_write_en;
logic top_13_3_clk;
logic top_13_3_reset;
logic [31:0] top_13_3_out;
logic top_13_3_done;
logic [31:0] left_13_3_in;
logic left_13_3_write_en;
logic left_13_3_clk;
logic left_13_3_reset;
logic [31:0] left_13_3_out;
logic left_13_3_done;
logic [31:0] pe_13_4_top;
logic [31:0] pe_13_4_left;
logic pe_13_4_mul_ready;
logic [31:0] pe_13_4_out;
logic pe_13_4_go;
logic pe_13_4_clk;
logic pe_13_4_reset;
logic pe_13_4_done;
logic [31:0] top_13_4_in;
logic top_13_4_write_en;
logic top_13_4_clk;
logic top_13_4_reset;
logic [31:0] top_13_4_out;
logic top_13_4_done;
logic [31:0] left_13_4_in;
logic left_13_4_write_en;
logic left_13_4_clk;
logic left_13_4_reset;
logic [31:0] left_13_4_out;
logic left_13_4_done;
logic [31:0] pe_13_5_top;
logic [31:0] pe_13_5_left;
logic pe_13_5_mul_ready;
logic [31:0] pe_13_5_out;
logic pe_13_5_go;
logic pe_13_5_clk;
logic pe_13_5_reset;
logic pe_13_5_done;
logic [31:0] top_13_5_in;
logic top_13_5_write_en;
logic top_13_5_clk;
logic top_13_5_reset;
logic [31:0] top_13_5_out;
logic top_13_5_done;
logic [31:0] left_13_5_in;
logic left_13_5_write_en;
logic left_13_5_clk;
logic left_13_5_reset;
logic [31:0] left_13_5_out;
logic left_13_5_done;
logic [31:0] pe_13_6_top;
logic [31:0] pe_13_6_left;
logic pe_13_6_mul_ready;
logic [31:0] pe_13_6_out;
logic pe_13_6_go;
logic pe_13_6_clk;
logic pe_13_6_reset;
logic pe_13_6_done;
logic [31:0] top_13_6_in;
logic top_13_6_write_en;
logic top_13_6_clk;
logic top_13_6_reset;
logic [31:0] top_13_6_out;
logic top_13_6_done;
logic [31:0] left_13_6_in;
logic left_13_6_write_en;
logic left_13_6_clk;
logic left_13_6_reset;
logic [31:0] left_13_6_out;
logic left_13_6_done;
logic [31:0] pe_13_7_top;
logic [31:0] pe_13_7_left;
logic pe_13_7_mul_ready;
logic [31:0] pe_13_7_out;
logic pe_13_7_go;
logic pe_13_7_clk;
logic pe_13_7_reset;
logic pe_13_7_done;
logic [31:0] top_13_7_in;
logic top_13_7_write_en;
logic top_13_7_clk;
logic top_13_7_reset;
logic [31:0] top_13_7_out;
logic top_13_7_done;
logic [31:0] left_13_7_in;
logic left_13_7_write_en;
logic left_13_7_clk;
logic left_13_7_reset;
logic [31:0] left_13_7_out;
logic left_13_7_done;
logic [31:0] pe_13_8_top;
logic [31:0] pe_13_8_left;
logic pe_13_8_mul_ready;
logic [31:0] pe_13_8_out;
logic pe_13_8_go;
logic pe_13_8_clk;
logic pe_13_8_reset;
logic pe_13_8_done;
logic [31:0] top_13_8_in;
logic top_13_8_write_en;
logic top_13_8_clk;
logic top_13_8_reset;
logic [31:0] top_13_8_out;
logic top_13_8_done;
logic [31:0] left_13_8_in;
logic left_13_8_write_en;
logic left_13_8_clk;
logic left_13_8_reset;
logic [31:0] left_13_8_out;
logic left_13_8_done;
logic [31:0] pe_13_9_top;
logic [31:0] pe_13_9_left;
logic pe_13_9_mul_ready;
logic [31:0] pe_13_9_out;
logic pe_13_9_go;
logic pe_13_9_clk;
logic pe_13_9_reset;
logic pe_13_9_done;
logic [31:0] top_13_9_in;
logic top_13_9_write_en;
logic top_13_9_clk;
logic top_13_9_reset;
logic [31:0] top_13_9_out;
logic top_13_9_done;
logic [31:0] left_13_9_in;
logic left_13_9_write_en;
logic left_13_9_clk;
logic left_13_9_reset;
logic [31:0] left_13_9_out;
logic left_13_9_done;
logic [31:0] pe_13_10_top;
logic [31:0] pe_13_10_left;
logic pe_13_10_mul_ready;
logic [31:0] pe_13_10_out;
logic pe_13_10_go;
logic pe_13_10_clk;
logic pe_13_10_reset;
logic pe_13_10_done;
logic [31:0] top_13_10_in;
logic top_13_10_write_en;
logic top_13_10_clk;
logic top_13_10_reset;
logic [31:0] top_13_10_out;
logic top_13_10_done;
logic [31:0] left_13_10_in;
logic left_13_10_write_en;
logic left_13_10_clk;
logic left_13_10_reset;
logic [31:0] left_13_10_out;
logic left_13_10_done;
logic [31:0] pe_13_11_top;
logic [31:0] pe_13_11_left;
logic pe_13_11_mul_ready;
logic [31:0] pe_13_11_out;
logic pe_13_11_go;
logic pe_13_11_clk;
logic pe_13_11_reset;
logic pe_13_11_done;
logic [31:0] top_13_11_in;
logic top_13_11_write_en;
logic top_13_11_clk;
logic top_13_11_reset;
logic [31:0] top_13_11_out;
logic top_13_11_done;
logic [31:0] left_13_11_in;
logic left_13_11_write_en;
logic left_13_11_clk;
logic left_13_11_reset;
logic [31:0] left_13_11_out;
logic left_13_11_done;
logic [31:0] pe_13_12_top;
logic [31:0] pe_13_12_left;
logic pe_13_12_mul_ready;
logic [31:0] pe_13_12_out;
logic pe_13_12_go;
logic pe_13_12_clk;
logic pe_13_12_reset;
logic pe_13_12_done;
logic [31:0] top_13_12_in;
logic top_13_12_write_en;
logic top_13_12_clk;
logic top_13_12_reset;
logic [31:0] top_13_12_out;
logic top_13_12_done;
logic [31:0] left_13_12_in;
logic left_13_12_write_en;
logic left_13_12_clk;
logic left_13_12_reset;
logic [31:0] left_13_12_out;
logic left_13_12_done;
logic [31:0] pe_13_13_top;
logic [31:0] pe_13_13_left;
logic pe_13_13_mul_ready;
logic [31:0] pe_13_13_out;
logic pe_13_13_go;
logic pe_13_13_clk;
logic pe_13_13_reset;
logic pe_13_13_done;
logic [31:0] top_13_13_in;
logic top_13_13_write_en;
logic top_13_13_clk;
logic top_13_13_reset;
logic [31:0] top_13_13_out;
logic top_13_13_done;
logic [31:0] left_13_13_in;
logic left_13_13_write_en;
logic left_13_13_clk;
logic left_13_13_reset;
logic [31:0] left_13_13_out;
logic left_13_13_done;
logic [31:0] pe_13_14_top;
logic [31:0] pe_13_14_left;
logic pe_13_14_mul_ready;
logic [31:0] pe_13_14_out;
logic pe_13_14_go;
logic pe_13_14_clk;
logic pe_13_14_reset;
logic pe_13_14_done;
logic [31:0] top_13_14_in;
logic top_13_14_write_en;
logic top_13_14_clk;
logic top_13_14_reset;
logic [31:0] top_13_14_out;
logic top_13_14_done;
logic [31:0] left_13_14_in;
logic left_13_14_write_en;
logic left_13_14_clk;
logic left_13_14_reset;
logic [31:0] left_13_14_out;
logic left_13_14_done;
logic [31:0] pe_13_15_top;
logic [31:0] pe_13_15_left;
logic pe_13_15_mul_ready;
logic [31:0] pe_13_15_out;
logic pe_13_15_go;
logic pe_13_15_clk;
logic pe_13_15_reset;
logic pe_13_15_done;
logic [31:0] top_13_15_in;
logic top_13_15_write_en;
logic top_13_15_clk;
logic top_13_15_reset;
logic [31:0] top_13_15_out;
logic top_13_15_done;
logic [31:0] left_13_15_in;
logic left_13_15_write_en;
logic left_13_15_clk;
logic left_13_15_reset;
logic [31:0] left_13_15_out;
logic left_13_15_done;
logic [31:0] pe_14_0_top;
logic [31:0] pe_14_0_left;
logic pe_14_0_mul_ready;
logic [31:0] pe_14_0_out;
logic pe_14_0_go;
logic pe_14_0_clk;
logic pe_14_0_reset;
logic pe_14_0_done;
logic [31:0] top_14_0_in;
logic top_14_0_write_en;
logic top_14_0_clk;
logic top_14_0_reset;
logic [31:0] top_14_0_out;
logic top_14_0_done;
logic [31:0] left_14_0_in;
logic left_14_0_write_en;
logic left_14_0_clk;
logic left_14_0_reset;
logic [31:0] left_14_0_out;
logic left_14_0_done;
logic [31:0] pe_14_1_top;
logic [31:0] pe_14_1_left;
logic pe_14_1_mul_ready;
logic [31:0] pe_14_1_out;
logic pe_14_1_go;
logic pe_14_1_clk;
logic pe_14_1_reset;
logic pe_14_1_done;
logic [31:0] top_14_1_in;
logic top_14_1_write_en;
logic top_14_1_clk;
logic top_14_1_reset;
logic [31:0] top_14_1_out;
logic top_14_1_done;
logic [31:0] left_14_1_in;
logic left_14_1_write_en;
logic left_14_1_clk;
logic left_14_1_reset;
logic [31:0] left_14_1_out;
logic left_14_1_done;
logic [31:0] pe_14_2_top;
logic [31:0] pe_14_2_left;
logic pe_14_2_mul_ready;
logic [31:0] pe_14_2_out;
logic pe_14_2_go;
logic pe_14_2_clk;
logic pe_14_2_reset;
logic pe_14_2_done;
logic [31:0] top_14_2_in;
logic top_14_2_write_en;
logic top_14_2_clk;
logic top_14_2_reset;
logic [31:0] top_14_2_out;
logic top_14_2_done;
logic [31:0] left_14_2_in;
logic left_14_2_write_en;
logic left_14_2_clk;
logic left_14_2_reset;
logic [31:0] left_14_2_out;
logic left_14_2_done;
logic [31:0] pe_14_3_top;
logic [31:0] pe_14_3_left;
logic pe_14_3_mul_ready;
logic [31:0] pe_14_3_out;
logic pe_14_3_go;
logic pe_14_3_clk;
logic pe_14_3_reset;
logic pe_14_3_done;
logic [31:0] top_14_3_in;
logic top_14_3_write_en;
logic top_14_3_clk;
logic top_14_3_reset;
logic [31:0] top_14_3_out;
logic top_14_3_done;
logic [31:0] left_14_3_in;
logic left_14_3_write_en;
logic left_14_3_clk;
logic left_14_3_reset;
logic [31:0] left_14_3_out;
logic left_14_3_done;
logic [31:0] pe_14_4_top;
logic [31:0] pe_14_4_left;
logic pe_14_4_mul_ready;
logic [31:0] pe_14_4_out;
logic pe_14_4_go;
logic pe_14_4_clk;
logic pe_14_4_reset;
logic pe_14_4_done;
logic [31:0] top_14_4_in;
logic top_14_4_write_en;
logic top_14_4_clk;
logic top_14_4_reset;
logic [31:0] top_14_4_out;
logic top_14_4_done;
logic [31:0] left_14_4_in;
logic left_14_4_write_en;
logic left_14_4_clk;
logic left_14_4_reset;
logic [31:0] left_14_4_out;
logic left_14_4_done;
logic [31:0] pe_14_5_top;
logic [31:0] pe_14_5_left;
logic pe_14_5_mul_ready;
logic [31:0] pe_14_5_out;
logic pe_14_5_go;
logic pe_14_5_clk;
logic pe_14_5_reset;
logic pe_14_5_done;
logic [31:0] top_14_5_in;
logic top_14_5_write_en;
logic top_14_5_clk;
logic top_14_5_reset;
logic [31:0] top_14_5_out;
logic top_14_5_done;
logic [31:0] left_14_5_in;
logic left_14_5_write_en;
logic left_14_5_clk;
logic left_14_5_reset;
logic [31:0] left_14_5_out;
logic left_14_5_done;
logic [31:0] pe_14_6_top;
logic [31:0] pe_14_6_left;
logic pe_14_6_mul_ready;
logic [31:0] pe_14_6_out;
logic pe_14_6_go;
logic pe_14_6_clk;
logic pe_14_6_reset;
logic pe_14_6_done;
logic [31:0] top_14_6_in;
logic top_14_6_write_en;
logic top_14_6_clk;
logic top_14_6_reset;
logic [31:0] top_14_6_out;
logic top_14_6_done;
logic [31:0] left_14_6_in;
logic left_14_6_write_en;
logic left_14_6_clk;
logic left_14_6_reset;
logic [31:0] left_14_6_out;
logic left_14_6_done;
logic [31:0] pe_14_7_top;
logic [31:0] pe_14_7_left;
logic pe_14_7_mul_ready;
logic [31:0] pe_14_7_out;
logic pe_14_7_go;
logic pe_14_7_clk;
logic pe_14_7_reset;
logic pe_14_7_done;
logic [31:0] top_14_7_in;
logic top_14_7_write_en;
logic top_14_7_clk;
logic top_14_7_reset;
logic [31:0] top_14_7_out;
logic top_14_7_done;
logic [31:0] left_14_7_in;
logic left_14_7_write_en;
logic left_14_7_clk;
logic left_14_7_reset;
logic [31:0] left_14_7_out;
logic left_14_7_done;
logic [31:0] pe_14_8_top;
logic [31:0] pe_14_8_left;
logic pe_14_8_mul_ready;
logic [31:0] pe_14_8_out;
logic pe_14_8_go;
logic pe_14_8_clk;
logic pe_14_8_reset;
logic pe_14_8_done;
logic [31:0] top_14_8_in;
logic top_14_8_write_en;
logic top_14_8_clk;
logic top_14_8_reset;
logic [31:0] top_14_8_out;
logic top_14_8_done;
logic [31:0] left_14_8_in;
logic left_14_8_write_en;
logic left_14_8_clk;
logic left_14_8_reset;
logic [31:0] left_14_8_out;
logic left_14_8_done;
logic [31:0] pe_14_9_top;
logic [31:0] pe_14_9_left;
logic pe_14_9_mul_ready;
logic [31:0] pe_14_9_out;
logic pe_14_9_go;
logic pe_14_9_clk;
logic pe_14_9_reset;
logic pe_14_9_done;
logic [31:0] top_14_9_in;
logic top_14_9_write_en;
logic top_14_9_clk;
logic top_14_9_reset;
logic [31:0] top_14_9_out;
logic top_14_9_done;
logic [31:0] left_14_9_in;
logic left_14_9_write_en;
logic left_14_9_clk;
logic left_14_9_reset;
logic [31:0] left_14_9_out;
logic left_14_9_done;
logic [31:0] pe_14_10_top;
logic [31:0] pe_14_10_left;
logic pe_14_10_mul_ready;
logic [31:0] pe_14_10_out;
logic pe_14_10_go;
logic pe_14_10_clk;
logic pe_14_10_reset;
logic pe_14_10_done;
logic [31:0] top_14_10_in;
logic top_14_10_write_en;
logic top_14_10_clk;
logic top_14_10_reset;
logic [31:0] top_14_10_out;
logic top_14_10_done;
logic [31:0] left_14_10_in;
logic left_14_10_write_en;
logic left_14_10_clk;
logic left_14_10_reset;
logic [31:0] left_14_10_out;
logic left_14_10_done;
logic [31:0] pe_14_11_top;
logic [31:0] pe_14_11_left;
logic pe_14_11_mul_ready;
logic [31:0] pe_14_11_out;
logic pe_14_11_go;
logic pe_14_11_clk;
logic pe_14_11_reset;
logic pe_14_11_done;
logic [31:0] top_14_11_in;
logic top_14_11_write_en;
logic top_14_11_clk;
logic top_14_11_reset;
logic [31:0] top_14_11_out;
logic top_14_11_done;
logic [31:0] left_14_11_in;
logic left_14_11_write_en;
logic left_14_11_clk;
logic left_14_11_reset;
logic [31:0] left_14_11_out;
logic left_14_11_done;
logic [31:0] pe_14_12_top;
logic [31:0] pe_14_12_left;
logic pe_14_12_mul_ready;
logic [31:0] pe_14_12_out;
logic pe_14_12_go;
logic pe_14_12_clk;
logic pe_14_12_reset;
logic pe_14_12_done;
logic [31:0] top_14_12_in;
logic top_14_12_write_en;
logic top_14_12_clk;
logic top_14_12_reset;
logic [31:0] top_14_12_out;
logic top_14_12_done;
logic [31:0] left_14_12_in;
logic left_14_12_write_en;
logic left_14_12_clk;
logic left_14_12_reset;
logic [31:0] left_14_12_out;
logic left_14_12_done;
logic [31:0] pe_14_13_top;
logic [31:0] pe_14_13_left;
logic pe_14_13_mul_ready;
logic [31:0] pe_14_13_out;
logic pe_14_13_go;
logic pe_14_13_clk;
logic pe_14_13_reset;
logic pe_14_13_done;
logic [31:0] top_14_13_in;
logic top_14_13_write_en;
logic top_14_13_clk;
logic top_14_13_reset;
logic [31:0] top_14_13_out;
logic top_14_13_done;
logic [31:0] left_14_13_in;
logic left_14_13_write_en;
logic left_14_13_clk;
logic left_14_13_reset;
logic [31:0] left_14_13_out;
logic left_14_13_done;
logic [31:0] pe_14_14_top;
logic [31:0] pe_14_14_left;
logic pe_14_14_mul_ready;
logic [31:0] pe_14_14_out;
logic pe_14_14_go;
logic pe_14_14_clk;
logic pe_14_14_reset;
logic pe_14_14_done;
logic [31:0] top_14_14_in;
logic top_14_14_write_en;
logic top_14_14_clk;
logic top_14_14_reset;
logic [31:0] top_14_14_out;
logic top_14_14_done;
logic [31:0] left_14_14_in;
logic left_14_14_write_en;
logic left_14_14_clk;
logic left_14_14_reset;
logic [31:0] left_14_14_out;
logic left_14_14_done;
logic [31:0] pe_14_15_top;
logic [31:0] pe_14_15_left;
logic pe_14_15_mul_ready;
logic [31:0] pe_14_15_out;
logic pe_14_15_go;
logic pe_14_15_clk;
logic pe_14_15_reset;
logic pe_14_15_done;
logic [31:0] top_14_15_in;
logic top_14_15_write_en;
logic top_14_15_clk;
logic top_14_15_reset;
logic [31:0] top_14_15_out;
logic top_14_15_done;
logic [31:0] left_14_15_in;
logic left_14_15_write_en;
logic left_14_15_clk;
logic left_14_15_reset;
logic [31:0] left_14_15_out;
logic left_14_15_done;
logic [31:0] pe_15_0_top;
logic [31:0] pe_15_0_left;
logic pe_15_0_mul_ready;
logic [31:0] pe_15_0_out;
logic pe_15_0_go;
logic pe_15_0_clk;
logic pe_15_0_reset;
logic pe_15_0_done;
logic [31:0] top_15_0_in;
logic top_15_0_write_en;
logic top_15_0_clk;
logic top_15_0_reset;
logic [31:0] top_15_0_out;
logic top_15_0_done;
logic [31:0] left_15_0_in;
logic left_15_0_write_en;
logic left_15_0_clk;
logic left_15_0_reset;
logic [31:0] left_15_0_out;
logic left_15_0_done;
logic [31:0] pe_15_1_top;
logic [31:0] pe_15_1_left;
logic pe_15_1_mul_ready;
logic [31:0] pe_15_1_out;
logic pe_15_1_go;
logic pe_15_1_clk;
logic pe_15_1_reset;
logic pe_15_1_done;
logic [31:0] top_15_1_in;
logic top_15_1_write_en;
logic top_15_1_clk;
logic top_15_1_reset;
logic [31:0] top_15_1_out;
logic top_15_1_done;
logic [31:0] left_15_1_in;
logic left_15_1_write_en;
logic left_15_1_clk;
logic left_15_1_reset;
logic [31:0] left_15_1_out;
logic left_15_1_done;
logic [31:0] pe_15_2_top;
logic [31:0] pe_15_2_left;
logic pe_15_2_mul_ready;
logic [31:0] pe_15_2_out;
logic pe_15_2_go;
logic pe_15_2_clk;
logic pe_15_2_reset;
logic pe_15_2_done;
logic [31:0] top_15_2_in;
logic top_15_2_write_en;
logic top_15_2_clk;
logic top_15_2_reset;
logic [31:0] top_15_2_out;
logic top_15_2_done;
logic [31:0] left_15_2_in;
logic left_15_2_write_en;
logic left_15_2_clk;
logic left_15_2_reset;
logic [31:0] left_15_2_out;
logic left_15_2_done;
logic [31:0] pe_15_3_top;
logic [31:0] pe_15_3_left;
logic pe_15_3_mul_ready;
logic [31:0] pe_15_3_out;
logic pe_15_3_go;
logic pe_15_3_clk;
logic pe_15_3_reset;
logic pe_15_3_done;
logic [31:0] top_15_3_in;
logic top_15_3_write_en;
logic top_15_3_clk;
logic top_15_3_reset;
logic [31:0] top_15_3_out;
logic top_15_3_done;
logic [31:0] left_15_3_in;
logic left_15_3_write_en;
logic left_15_3_clk;
logic left_15_3_reset;
logic [31:0] left_15_3_out;
logic left_15_3_done;
logic [31:0] pe_15_4_top;
logic [31:0] pe_15_4_left;
logic pe_15_4_mul_ready;
logic [31:0] pe_15_4_out;
logic pe_15_4_go;
logic pe_15_4_clk;
logic pe_15_4_reset;
logic pe_15_4_done;
logic [31:0] top_15_4_in;
logic top_15_4_write_en;
logic top_15_4_clk;
logic top_15_4_reset;
logic [31:0] top_15_4_out;
logic top_15_4_done;
logic [31:0] left_15_4_in;
logic left_15_4_write_en;
logic left_15_4_clk;
logic left_15_4_reset;
logic [31:0] left_15_4_out;
logic left_15_4_done;
logic [31:0] pe_15_5_top;
logic [31:0] pe_15_5_left;
logic pe_15_5_mul_ready;
logic [31:0] pe_15_5_out;
logic pe_15_5_go;
logic pe_15_5_clk;
logic pe_15_5_reset;
logic pe_15_5_done;
logic [31:0] top_15_5_in;
logic top_15_5_write_en;
logic top_15_5_clk;
logic top_15_5_reset;
logic [31:0] top_15_5_out;
logic top_15_5_done;
logic [31:0] left_15_5_in;
logic left_15_5_write_en;
logic left_15_5_clk;
logic left_15_5_reset;
logic [31:0] left_15_5_out;
logic left_15_5_done;
logic [31:0] pe_15_6_top;
logic [31:0] pe_15_6_left;
logic pe_15_6_mul_ready;
logic [31:0] pe_15_6_out;
logic pe_15_6_go;
logic pe_15_6_clk;
logic pe_15_6_reset;
logic pe_15_6_done;
logic [31:0] top_15_6_in;
logic top_15_6_write_en;
logic top_15_6_clk;
logic top_15_6_reset;
logic [31:0] top_15_6_out;
logic top_15_6_done;
logic [31:0] left_15_6_in;
logic left_15_6_write_en;
logic left_15_6_clk;
logic left_15_6_reset;
logic [31:0] left_15_6_out;
logic left_15_6_done;
logic [31:0] pe_15_7_top;
logic [31:0] pe_15_7_left;
logic pe_15_7_mul_ready;
logic [31:0] pe_15_7_out;
logic pe_15_7_go;
logic pe_15_7_clk;
logic pe_15_7_reset;
logic pe_15_7_done;
logic [31:0] top_15_7_in;
logic top_15_7_write_en;
logic top_15_7_clk;
logic top_15_7_reset;
logic [31:0] top_15_7_out;
logic top_15_7_done;
logic [31:0] left_15_7_in;
logic left_15_7_write_en;
logic left_15_7_clk;
logic left_15_7_reset;
logic [31:0] left_15_7_out;
logic left_15_7_done;
logic [31:0] pe_15_8_top;
logic [31:0] pe_15_8_left;
logic pe_15_8_mul_ready;
logic [31:0] pe_15_8_out;
logic pe_15_8_go;
logic pe_15_8_clk;
logic pe_15_8_reset;
logic pe_15_8_done;
logic [31:0] top_15_8_in;
logic top_15_8_write_en;
logic top_15_8_clk;
logic top_15_8_reset;
logic [31:0] top_15_8_out;
logic top_15_8_done;
logic [31:0] left_15_8_in;
logic left_15_8_write_en;
logic left_15_8_clk;
logic left_15_8_reset;
logic [31:0] left_15_8_out;
logic left_15_8_done;
logic [31:0] pe_15_9_top;
logic [31:0] pe_15_9_left;
logic pe_15_9_mul_ready;
logic [31:0] pe_15_9_out;
logic pe_15_9_go;
logic pe_15_9_clk;
logic pe_15_9_reset;
logic pe_15_9_done;
logic [31:0] top_15_9_in;
logic top_15_9_write_en;
logic top_15_9_clk;
logic top_15_9_reset;
logic [31:0] top_15_9_out;
logic top_15_9_done;
logic [31:0] left_15_9_in;
logic left_15_9_write_en;
logic left_15_9_clk;
logic left_15_9_reset;
logic [31:0] left_15_9_out;
logic left_15_9_done;
logic [31:0] pe_15_10_top;
logic [31:0] pe_15_10_left;
logic pe_15_10_mul_ready;
logic [31:0] pe_15_10_out;
logic pe_15_10_go;
logic pe_15_10_clk;
logic pe_15_10_reset;
logic pe_15_10_done;
logic [31:0] top_15_10_in;
logic top_15_10_write_en;
logic top_15_10_clk;
logic top_15_10_reset;
logic [31:0] top_15_10_out;
logic top_15_10_done;
logic [31:0] left_15_10_in;
logic left_15_10_write_en;
logic left_15_10_clk;
logic left_15_10_reset;
logic [31:0] left_15_10_out;
logic left_15_10_done;
logic [31:0] pe_15_11_top;
logic [31:0] pe_15_11_left;
logic pe_15_11_mul_ready;
logic [31:0] pe_15_11_out;
logic pe_15_11_go;
logic pe_15_11_clk;
logic pe_15_11_reset;
logic pe_15_11_done;
logic [31:0] top_15_11_in;
logic top_15_11_write_en;
logic top_15_11_clk;
logic top_15_11_reset;
logic [31:0] top_15_11_out;
logic top_15_11_done;
logic [31:0] left_15_11_in;
logic left_15_11_write_en;
logic left_15_11_clk;
logic left_15_11_reset;
logic [31:0] left_15_11_out;
logic left_15_11_done;
logic [31:0] pe_15_12_top;
logic [31:0] pe_15_12_left;
logic pe_15_12_mul_ready;
logic [31:0] pe_15_12_out;
logic pe_15_12_go;
logic pe_15_12_clk;
logic pe_15_12_reset;
logic pe_15_12_done;
logic [31:0] top_15_12_in;
logic top_15_12_write_en;
logic top_15_12_clk;
logic top_15_12_reset;
logic [31:0] top_15_12_out;
logic top_15_12_done;
logic [31:0] left_15_12_in;
logic left_15_12_write_en;
logic left_15_12_clk;
logic left_15_12_reset;
logic [31:0] left_15_12_out;
logic left_15_12_done;
logic [31:0] pe_15_13_top;
logic [31:0] pe_15_13_left;
logic pe_15_13_mul_ready;
logic [31:0] pe_15_13_out;
logic pe_15_13_go;
logic pe_15_13_clk;
logic pe_15_13_reset;
logic pe_15_13_done;
logic [31:0] top_15_13_in;
logic top_15_13_write_en;
logic top_15_13_clk;
logic top_15_13_reset;
logic [31:0] top_15_13_out;
logic top_15_13_done;
logic [31:0] left_15_13_in;
logic left_15_13_write_en;
logic left_15_13_clk;
logic left_15_13_reset;
logic [31:0] left_15_13_out;
logic left_15_13_done;
logic [31:0] pe_15_14_top;
logic [31:0] pe_15_14_left;
logic pe_15_14_mul_ready;
logic [31:0] pe_15_14_out;
logic pe_15_14_go;
logic pe_15_14_clk;
logic pe_15_14_reset;
logic pe_15_14_done;
logic [31:0] top_15_14_in;
logic top_15_14_write_en;
logic top_15_14_clk;
logic top_15_14_reset;
logic [31:0] top_15_14_out;
logic top_15_14_done;
logic [31:0] left_15_14_in;
logic left_15_14_write_en;
logic left_15_14_clk;
logic left_15_14_reset;
logic [31:0] left_15_14_out;
logic left_15_14_done;
logic [31:0] pe_15_15_top;
logic [31:0] pe_15_15_left;
logic pe_15_15_mul_ready;
logic [31:0] pe_15_15_out;
logic pe_15_15_go;
logic pe_15_15_clk;
logic pe_15_15_reset;
logic pe_15_15_done;
logic [31:0] top_15_15_in;
logic top_15_15_write_en;
logic top_15_15_clk;
logic top_15_15_reset;
logic [31:0] top_15_15_out;
logic top_15_15_done;
logic [31:0] left_15_15_in;
logic left_15_15_write_en;
logic left_15_15_clk;
logic left_15_15_reset;
logic [31:0] left_15_15_out;
logic left_15_15_done;
logic [4:0] t0_idx_in;
logic t0_idx_write_en;
logic t0_idx_clk;
logic t0_idx_reset;
logic [4:0] t0_idx_out;
logic t0_idx_done;
logic [4:0] t0_add_left;
logic [4:0] t0_add_right;
logic [4:0] t0_add_out;
logic [4:0] t1_idx_in;
logic t1_idx_write_en;
logic t1_idx_clk;
logic t1_idx_reset;
logic [4:0] t1_idx_out;
logic t1_idx_done;
logic [4:0] t1_add_left;
logic [4:0] t1_add_right;
logic [4:0] t1_add_out;
logic [4:0] t2_idx_in;
logic t2_idx_write_en;
logic t2_idx_clk;
logic t2_idx_reset;
logic [4:0] t2_idx_out;
logic t2_idx_done;
logic [4:0] t2_add_left;
logic [4:0] t2_add_right;
logic [4:0] t2_add_out;
logic [4:0] t3_idx_in;
logic t3_idx_write_en;
logic t3_idx_clk;
logic t3_idx_reset;
logic [4:0] t3_idx_out;
logic t3_idx_done;
logic [4:0] t3_add_left;
logic [4:0] t3_add_right;
logic [4:0] t3_add_out;
logic [4:0] t4_idx_in;
logic t4_idx_write_en;
logic t4_idx_clk;
logic t4_idx_reset;
logic [4:0] t4_idx_out;
logic t4_idx_done;
logic [4:0] t4_add_left;
logic [4:0] t4_add_right;
logic [4:0] t4_add_out;
logic [4:0] t5_idx_in;
logic t5_idx_write_en;
logic t5_idx_clk;
logic t5_idx_reset;
logic [4:0] t5_idx_out;
logic t5_idx_done;
logic [4:0] t5_add_left;
logic [4:0] t5_add_right;
logic [4:0] t5_add_out;
logic [4:0] t6_idx_in;
logic t6_idx_write_en;
logic t6_idx_clk;
logic t6_idx_reset;
logic [4:0] t6_idx_out;
logic t6_idx_done;
logic [4:0] t6_add_left;
logic [4:0] t6_add_right;
logic [4:0] t6_add_out;
logic [4:0] t7_idx_in;
logic t7_idx_write_en;
logic t7_idx_clk;
logic t7_idx_reset;
logic [4:0] t7_idx_out;
logic t7_idx_done;
logic [4:0] t7_add_left;
logic [4:0] t7_add_right;
logic [4:0] t7_add_out;
logic [4:0] t8_idx_in;
logic t8_idx_write_en;
logic t8_idx_clk;
logic t8_idx_reset;
logic [4:0] t8_idx_out;
logic t8_idx_done;
logic [4:0] t8_add_left;
logic [4:0] t8_add_right;
logic [4:0] t8_add_out;
logic [4:0] t9_idx_in;
logic t9_idx_write_en;
logic t9_idx_clk;
logic t9_idx_reset;
logic [4:0] t9_idx_out;
logic t9_idx_done;
logic [4:0] t9_add_left;
logic [4:0] t9_add_right;
logic [4:0] t9_add_out;
logic [4:0] t10_idx_in;
logic t10_idx_write_en;
logic t10_idx_clk;
logic t10_idx_reset;
logic [4:0] t10_idx_out;
logic t10_idx_done;
logic [4:0] t10_add_left;
logic [4:0] t10_add_right;
logic [4:0] t10_add_out;
logic [4:0] t11_idx_in;
logic t11_idx_write_en;
logic t11_idx_clk;
logic t11_idx_reset;
logic [4:0] t11_idx_out;
logic t11_idx_done;
logic [4:0] t11_add_left;
logic [4:0] t11_add_right;
logic [4:0] t11_add_out;
logic [4:0] t12_idx_in;
logic t12_idx_write_en;
logic t12_idx_clk;
logic t12_idx_reset;
logic [4:0] t12_idx_out;
logic t12_idx_done;
logic [4:0] t12_add_left;
logic [4:0] t12_add_right;
logic [4:0] t12_add_out;
logic [4:0] t13_idx_in;
logic t13_idx_write_en;
logic t13_idx_clk;
logic t13_idx_reset;
logic [4:0] t13_idx_out;
logic t13_idx_done;
logic [4:0] t13_add_left;
logic [4:0] t13_add_right;
logic [4:0] t13_add_out;
logic [4:0] t14_idx_in;
logic t14_idx_write_en;
logic t14_idx_clk;
logic t14_idx_reset;
logic [4:0] t14_idx_out;
logic t14_idx_done;
logic [4:0] t14_add_left;
logic [4:0] t14_add_right;
logic [4:0] t14_add_out;
logic [4:0] t15_idx_in;
logic t15_idx_write_en;
logic t15_idx_clk;
logic t15_idx_reset;
logic [4:0] t15_idx_out;
logic t15_idx_done;
logic [4:0] t15_add_left;
logic [4:0] t15_add_right;
logic [4:0] t15_add_out;
logic [4:0] l0_idx_in;
logic l0_idx_write_en;
logic l0_idx_clk;
logic l0_idx_reset;
logic [4:0] l0_idx_out;
logic l0_idx_done;
logic [4:0] l0_add_left;
logic [4:0] l0_add_right;
logic [4:0] l0_add_out;
logic [4:0] l1_idx_in;
logic l1_idx_write_en;
logic l1_idx_clk;
logic l1_idx_reset;
logic [4:0] l1_idx_out;
logic l1_idx_done;
logic [4:0] l1_add_left;
logic [4:0] l1_add_right;
logic [4:0] l1_add_out;
logic [4:0] l2_idx_in;
logic l2_idx_write_en;
logic l2_idx_clk;
logic l2_idx_reset;
logic [4:0] l2_idx_out;
logic l2_idx_done;
logic [4:0] l2_add_left;
logic [4:0] l2_add_right;
logic [4:0] l2_add_out;
logic [4:0] l3_idx_in;
logic l3_idx_write_en;
logic l3_idx_clk;
logic l3_idx_reset;
logic [4:0] l3_idx_out;
logic l3_idx_done;
logic [4:0] l3_add_left;
logic [4:0] l3_add_right;
logic [4:0] l3_add_out;
logic [4:0] l4_idx_in;
logic l4_idx_write_en;
logic l4_idx_clk;
logic l4_idx_reset;
logic [4:0] l4_idx_out;
logic l4_idx_done;
logic [4:0] l4_add_left;
logic [4:0] l4_add_right;
logic [4:0] l4_add_out;
logic [4:0] l5_idx_in;
logic l5_idx_write_en;
logic l5_idx_clk;
logic l5_idx_reset;
logic [4:0] l5_idx_out;
logic l5_idx_done;
logic [4:0] l5_add_left;
logic [4:0] l5_add_right;
logic [4:0] l5_add_out;
logic [4:0] l6_idx_in;
logic l6_idx_write_en;
logic l6_idx_clk;
logic l6_idx_reset;
logic [4:0] l6_idx_out;
logic l6_idx_done;
logic [4:0] l6_add_left;
logic [4:0] l6_add_right;
logic [4:0] l6_add_out;
logic [4:0] l7_idx_in;
logic l7_idx_write_en;
logic l7_idx_clk;
logic l7_idx_reset;
logic [4:0] l7_idx_out;
logic l7_idx_done;
logic [4:0] l7_add_left;
logic [4:0] l7_add_right;
logic [4:0] l7_add_out;
logic [4:0] l8_idx_in;
logic l8_idx_write_en;
logic l8_idx_clk;
logic l8_idx_reset;
logic [4:0] l8_idx_out;
logic l8_idx_done;
logic [4:0] l8_add_left;
logic [4:0] l8_add_right;
logic [4:0] l8_add_out;
logic [4:0] l9_idx_in;
logic l9_idx_write_en;
logic l9_idx_clk;
logic l9_idx_reset;
logic [4:0] l9_idx_out;
logic l9_idx_done;
logic [4:0] l9_add_left;
logic [4:0] l9_add_right;
logic [4:0] l9_add_out;
logic [4:0] l10_idx_in;
logic l10_idx_write_en;
logic l10_idx_clk;
logic l10_idx_reset;
logic [4:0] l10_idx_out;
logic l10_idx_done;
logic [4:0] l10_add_left;
logic [4:0] l10_add_right;
logic [4:0] l10_add_out;
logic [4:0] l11_idx_in;
logic l11_idx_write_en;
logic l11_idx_clk;
logic l11_idx_reset;
logic [4:0] l11_idx_out;
logic l11_idx_done;
logic [4:0] l11_add_left;
logic [4:0] l11_add_right;
logic [4:0] l11_add_out;
logic [4:0] l12_idx_in;
logic l12_idx_write_en;
logic l12_idx_clk;
logic l12_idx_reset;
logic [4:0] l12_idx_out;
logic l12_idx_done;
logic [4:0] l12_add_left;
logic [4:0] l12_add_right;
logic [4:0] l12_add_out;
logic [4:0] l13_idx_in;
logic l13_idx_write_en;
logic l13_idx_clk;
logic l13_idx_reset;
logic [4:0] l13_idx_out;
logic l13_idx_done;
logic [4:0] l13_add_left;
logic [4:0] l13_add_right;
logic [4:0] l13_add_out;
logic [4:0] l14_idx_in;
logic l14_idx_write_en;
logic l14_idx_clk;
logic l14_idx_reset;
logic [4:0] l14_idx_out;
logic l14_idx_done;
logic [4:0] l14_add_left;
logic [4:0] l14_add_right;
logic [4:0] l14_add_out;
logic [4:0] l15_idx_in;
logic l15_idx_write_en;
logic l15_idx_clk;
logic l15_idx_reset;
logic [4:0] l15_idx_out;
logic l15_idx_done;
logic [4:0] l15_add_left;
logic [4:0] l15_add_right;
logic [4:0] l15_add_out;
logic [5:0] idx_in;
logic idx_write_en;
logic idx_clk;
logic idx_reset;
logic [5:0] idx_out;
logic idx_done;
logic [5:0] idx_add_left;
logic [5:0] idx_add_right;
logic [5:0] idx_add_out;
logic idx_between_16_20_reg_in;
logic idx_between_16_20_reg_write_en;
logic idx_between_16_20_reg_clk;
logic idx_between_16_20_reg_reset;
logic idx_between_16_20_reg_out;
logic idx_between_16_20_reg_done;
logic [5:0] index_lt_20_left;
logic [5:0] index_lt_20_right;
logic index_lt_20_out;
logic [5:0] index_ge_16_left;
logic [5:0] index_ge_16_right;
logic index_ge_16_out;
logic idx_between_16_20_comb_left;
logic idx_between_16_20_comb_right;
logic idx_between_16_20_comb_out;
logic idx_between_26_30_reg_in;
logic idx_between_26_30_reg_write_en;
logic idx_between_26_30_reg_clk;
logic idx_between_26_30_reg_reset;
logic idx_between_26_30_reg_out;
logic idx_between_26_30_reg_done;
logic [5:0] index_lt_30_left;
logic [5:0] index_lt_30_right;
logic index_lt_30_out;
logic [5:0] index_ge_26_left;
logic [5:0] index_ge_26_right;
logic index_ge_26_out;
logic idx_between_26_30_comb_left;
logic idx_between_26_30_comb_right;
logic idx_between_26_30_comb_out;
logic idx_between_30_46_reg_in;
logic idx_between_30_46_reg_write_en;
logic idx_between_30_46_reg_clk;
logic idx_between_30_46_reg_reset;
logic idx_between_30_46_reg_out;
logic idx_between_30_46_reg_done;
logic [5:0] index_lt_46_left;
logic [5:0] index_lt_46_right;
logic index_lt_46_out;
logic [5:0] index_ge_30_left;
logic [5:0] index_ge_30_right;
logic index_ge_30_out;
logic idx_between_30_46_comb_left;
logic idx_between_30_46_comb_right;
logic idx_between_30_46_comb_out;
logic idx_between_44_45_reg_in;
logic idx_between_44_45_reg_write_en;
logic idx_between_44_45_reg_clk;
logic idx_between_44_45_reg_reset;
logic idx_between_44_45_reg_out;
logic idx_between_44_45_reg_done;
logic [5:0] index_lt_45_left;
logic [5:0] index_lt_45_right;
logic index_lt_45_out;
logic [5:0] index_ge_44_left;
logic [5:0] index_ge_44_right;
logic index_ge_44_out;
logic idx_between_44_45_comb_left;
logic idx_between_44_45_comb_right;
logic idx_between_44_45_comb_out;
logic idx_between_25_41_reg_in;
logic idx_between_25_41_reg_write_en;
logic idx_between_25_41_reg_clk;
logic idx_between_25_41_reg_reset;
logic idx_between_25_41_reg_out;
logic idx_between_25_41_reg_done;
logic [5:0] index_lt_41_left;
logic [5:0] index_lt_41_right;
logic index_lt_41_out;
logic [5:0] index_ge_25_left;
logic [5:0] index_ge_25_right;
logic index_ge_25_out;
logic idx_between_25_41_comb_left;
logic idx_between_25_41_comb_right;
logic idx_between_25_41_comb_out;
logic idx_between_35_51_reg_in;
logic idx_between_35_51_reg_write_en;
logic idx_between_35_51_reg_clk;
logic idx_between_35_51_reg_reset;
logic idx_between_35_51_reg_out;
logic idx_between_35_51_reg_done;
logic [5:0] index_lt_51_left;
logic [5:0] index_lt_51_right;
logic index_lt_51_out;
logic [5:0] index_ge_35_left;
logic [5:0] index_ge_35_right;
logic index_ge_35_out;
logic idx_between_35_51_comb_left;
logic idx_between_35_51_comb_right;
logic idx_between_35_51_comb_out;
logic idx_between_22_26_reg_in;
logic idx_between_22_26_reg_write_en;
logic idx_between_22_26_reg_clk;
logic idx_between_22_26_reg_reset;
logic idx_between_22_26_reg_out;
logic idx_between_22_26_reg_done;
logic [5:0] index_lt_26_left;
logic [5:0] index_lt_26_right;
logic index_lt_26_out;
logic [5:0] index_ge_22_left;
logic [5:0] index_ge_22_right;
logic index_ge_22_out;
logic idx_between_22_26_comb_left;
logic idx_between_22_26_comb_right;
logic idx_between_22_26_comb_out;
logic idx_between_40_41_reg_in;
logic idx_between_40_41_reg_write_en;
logic idx_between_40_41_reg_clk;
logic idx_between_40_41_reg_reset;
logic idx_between_40_41_reg_out;
logic idx_between_40_41_reg_done;
logic [5:0] index_ge_40_left;
logic [5:0] index_ge_40_right;
logic index_ge_40_out;
logic idx_between_40_41_comb_left;
logic idx_between_40_41_comb_right;
logic idx_between_40_41_comb_out;
logic idx_between_17_21_reg_in;
logic idx_between_17_21_reg_write_en;
logic idx_between_17_21_reg_clk;
logic idx_between_17_21_reg_reset;
logic idx_between_17_21_reg_out;
logic idx_between_17_21_reg_done;
logic [5:0] index_lt_21_left;
logic [5:0] index_lt_21_right;
logic index_lt_21_out;
logic [5:0] index_ge_17_left;
logic [5:0] index_ge_17_right;
logic index_ge_17_out;
logic idx_between_17_21_comb_left;
logic idx_between_17_21_comb_right;
logic idx_between_17_21_comb_out;
logic idx_between_21_37_reg_in;
logic idx_between_21_37_reg_write_en;
logic idx_between_21_37_reg_clk;
logic idx_between_21_37_reg_reset;
logic idx_between_21_37_reg_out;
logic idx_between_21_37_reg_done;
logic [5:0] index_lt_37_left;
logic [5:0] index_lt_37_right;
logic index_lt_37_out;
logic [5:0] index_ge_21_left;
logic [5:0] index_ge_21_right;
logic index_ge_21_out;
logic idx_between_21_37_comb_left;
logic idx_between_21_37_comb_right;
logic idx_between_21_37_comb_out;
logic idx_between_31_47_reg_in;
logic idx_between_31_47_reg_write_en;
logic idx_between_31_47_reg_clk;
logic idx_between_31_47_reg_reset;
logic idx_between_31_47_reg_out;
logic idx_between_31_47_reg_done;
logic [5:0] index_lt_47_left;
logic [5:0] index_lt_47_right;
logic index_lt_47_out;
logic [5:0] index_ge_31_left;
logic [5:0] index_ge_31_right;
logic index_ge_31_out;
logic idx_between_31_47_comb_left;
logic idx_between_31_47_comb_right;
logic idx_between_31_47_comb_out;
logic idx_between_13_17_reg_in;
logic idx_between_13_17_reg_write_en;
logic idx_between_13_17_reg_clk;
logic idx_between_13_17_reg_reset;
logic idx_between_13_17_reg_out;
logic idx_between_13_17_reg_done;
logic [5:0] index_lt_17_left;
logic [5:0] index_lt_17_right;
logic index_lt_17_out;
logic [5:0] index_ge_13_left;
logic [5:0] index_ge_13_right;
logic index_ge_13_out;
logic idx_between_13_17_comb_left;
logic idx_between_13_17_comb_right;
logic idx_between_13_17_comb_out;
logic idx_between_27_43_reg_in;
logic idx_between_27_43_reg_write_en;
logic idx_between_27_43_reg_clk;
logic idx_between_27_43_reg_reset;
logic idx_between_27_43_reg_out;
logic idx_between_27_43_reg_done;
logic [5:0] index_lt_43_left;
logic [5:0] index_lt_43_right;
logic index_lt_43_out;
logic [5:0] index_ge_27_left;
logic [5:0] index_ge_27_right;
logic index_ge_27_out;
logic idx_between_27_43_comb_left;
logic idx_between_27_43_comb_right;
logic idx_between_27_43_comb_out;
logic idx_between_41_42_reg_in;
logic idx_between_41_42_reg_write_en;
logic idx_between_41_42_reg_clk;
logic idx_between_41_42_reg_reset;
logic idx_between_41_42_reg_out;
logic idx_between_41_42_reg_done;
logic [5:0] index_lt_42_left;
logic [5:0] index_lt_42_right;
logic index_lt_42_out;
logic [5:0] index_ge_41_left;
logic [5:0] index_ge_41_right;
logic index_ge_41_out;
logic idx_between_41_42_comb_left;
logic idx_between_41_42_comb_right;
logic idx_between_41_42_comb_out;
logic idx_between_23_27_reg_in;
logic idx_between_23_27_reg_write_en;
logic idx_between_23_27_reg_clk;
logic idx_between_23_27_reg_reset;
logic idx_between_23_27_reg_out;
logic idx_between_23_27_reg_done;
logic [5:0] index_lt_27_left;
logic [5:0] index_lt_27_right;
logic index_lt_27_out;
logic [5:0] index_ge_23_left;
logic [5:0] index_ge_23_right;
logic index_ge_23_out;
logic idx_between_23_27_comb_left;
logic idx_between_23_27_comb_right;
logic idx_between_23_27_comb_out;
logic idx_between_5_21_reg_in;
logic idx_between_5_21_reg_write_en;
logic idx_between_5_21_reg_clk;
logic idx_between_5_21_reg_reset;
logic idx_between_5_21_reg_out;
logic idx_between_5_21_reg_done;
logic [5:0] index_ge_5_left;
logic [5:0] index_ge_5_right;
logic index_ge_5_out;
logic idx_between_5_21_comb_left;
logic idx_between_5_21_comb_right;
logic idx_between_5_21_comb_out;
logic idx_between_0_16_reg_in;
logic idx_between_0_16_reg_write_en;
logic idx_between_0_16_reg_clk;
logic idx_between_0_16_reg_reset;
logic idx_between_0_16_reg_out;
logic idx_between_0_16_reg_done;
logic [5:0] index_lt_16_left;
logic [5:0] index_lt_16_right;
logic index_lt_16_out;
logic idx_between_1_17_reg_in;
logic idx_between_1_17_reg_write_en;
logic idx_between_1_17_reg_clk;
logic idx_between_1_17_reg_reset;
logic idx_between_1_17_reg_out;
logic idx_between_1_17_reg_done;
logic [5:0] index_ge_1_left;
logic [5:0] index_ge_1_right;
logic index_ge_1_out;
logic idx_between_1_17_comb_left;
logic idx_between_1_17_comb_right;
logic idx_between_1_17_comb_out;
logic idx_between_47_48_reg_in;
logic idx_between_47_48_reg_write_en;
logic idx_between_47_48_reg_clk;
logic idx_between_47_48_reg_reset;
logic idx_between_47_48_reg_out;
logic idx_between_47_48_reg_done;
logic [5:0] index_lt_48_left;
logic [5:0] index_lt_48_right;
logic index_lt_48_out;
logic [5:0] index_ge_47_left;
logic [5:0] index_ge_47_right;
logic index_ge_47_out;
logic idx_between_47_48_comb_left;
logic idx_between_47_48_comb_right;
logic idx_between_47_48_comb_out;
logic idx_between_24_28_reg_in;
logic idx_between_24_28_reg_write_en;
logic idx_between_24_28_reg_clk;
logic idx_between_24_28_reg_reset;
logic idx_between_24_28_reg_out;
logic idx_between_24_28_reg_done;
logic [5:0] index_lt_28_left;
logic [5:0] index_lt_28_right;
logic index_lt_28_out;
logic [5:0] index_ge_24_left;
logic [5:0] index_ge_24_right;
logic index_ge_24_out;
logic idx_between_24_28_comb_left;
logic idx_between_24_28_comb_right;
logic idx_between_24_28_comb_out;
logic idx_between_42_43_reg_in;
logic idx_between_42_43_reg_write_en;
logic idx_between_42_43_reg_clk;
logic idx_between_42_43_reg_reset;
logic idx_between_42_43_reg_out;
logic idx_between_42_43_reg_done;
logic [5:0] index_ge_42_left;
logic [5:0] index_ge_42_right;
logic index_ge_42_out;
logic idx_between_42_43_comb_left;
logic idx_between_42_43_comb_right;
logic idx_between_42_43_comb_out;
logic idx_between_33_49_reg_in;
logic idx_between_33_49_reg_write_en;
logic idx_between_33_49_reg_clk;
logic idx_between_33_49_reg_reset;
logic idx_between_33_49_reg_out;
logic idx_between_33_49_reg_done;
logic [5:0] index_lt_49_left;
logic [5:0] index_lt_49_right;
logic index_lt_49_out;
logic [5:0] index_ge_33_left;
logic [5:0] index_ge_33_right;
logic index_ge_33_out;
logic idx_between_33_49_comb_left;
logic idx_between_33_49_comb_right;
logic idx_between_33_49_comb_out;
logic idx_between_20_24_reg_in;
logic idx_between_20_24_reg_write_en;
logic idx_between_20_24_reg_clk;
logic idx_between_20_24_reg_reset;
logic idx_between_20_24_reg_out;
logic idx_between_20_24_reg_done;
logic [5:0] index_lt_24_left;
logic [5:0] index_lt_24_right;
logic index_lt_24_out;
logic [5:0] index_ge_20_left;
logic [5:0] index_ge_20_right;
logic index_ge_20_out;
logic idx_between_20_24_comb_left;
logic idx_between_20_24_comb_right;
logic idx_between_20_24_comb_out;
logic idx_between_38_39_reg_in;
logic idx_between_38_39_reg_write_en;
logic idx_between_38_39_reg_clk;
logic idx_between_38_39_reg_reset;
logic idx_between_38_39_reg_out;
logic idx_between_38_39_reg_done;
logic [5:0] index_lt_39_left;
logic [5:0] index_lt_39_right;
logic index_lt_39_out;
logic [5:0] index_ge_38_left;
logic [5:0] index_ge_38_right;
logic index_ge_38_out;
logic idx_between_38_39_comb_left;
logic idx_between_38_39_comb_right;
logic idx_between_38_39_comb_out;
logic idx_between_48_49_reg_in;
logic idx_between_48_49_reg_write_en;
logic idx_between_48_49_reg_clk;
logic idx_between_48_49_reg_reset;
logic idx_between_48_49_reg_out;
logic idx_between_48_49_reg_done;
logic [5:0] index_ge_48_left;
logic [5:0] index_ge_48_right;
logic index_ge_48_out;
logic idx_between_48_49_comb_left;
logic idx_between_48_49_comb_right;
logic idx_between_48_49_comb_out;
logic idx_between_29_45_reg_in;
logic idx_between_29_45_reg_write_en;
logic idx_between_29_45_reg_clk;
logic idx_between_29_45_reg_reset;
logic idx_between_29_45_reg_out;
logic idx_between_29_45_reg_done;
logic [5:0] index_ge_29_left;
logic [5:0] index_ge_29_right;
logic index_ge_29_out;
logic idx_between_29_45_comb_left;
logic idx_between_29_45_comb_right;
logic idx_between_29_45_comb_out;
logic idx_between_30_34_reg_in;
logic idx_between_30_34_reg_write_en;
logic idx_between_30_34_reg_clk;
logic idx_between_30_34_reg_reset;
logic idx_between_30_34_reg_out;
logic idx_between_30_34_reg_done;
logic [5:0] index_lt_34_left;
logic [5:0] index_lt_34_right;
logic index_lt_34_out;
logic idx_between_30_34_comb_left;
logic idx_between_30_34_comb_right;
logic idx_between_30_34_comb_out;
logic idx_between_25_29_reg_in;
logic idx_between_25_29_reg_write_en;
logic idx_between_25_29_reg_clk;
logic idx_between_25_29_reg_reset;
logic idx_between_25_29_reg_out;
logic idx_between_25_29_reg_done;
logic [5:0] index_lt_29_left;
logic [5:0] index_lt_29_right;
logic index_lt_29_out;
logic idx_between_25_29_comb_left;
logic idx_between_25_29_comb_right;
logic idx_between_25_29_comb_out;
logic idx_between_7_23_reg_in;
logic idx_between_7_23_reg_write_en;
logic idx_between_7_23_reg_clk;
logic idx_between_7_23_reg_reset;
logic idx_between_7_23_reg_out;
logic idx_between_7_23_reg_done;
logic [5:0] index_lt_23_left;
logic [5:0] index_lt_23_right;
logic index_lt_23_out;
logic [5:0] index_ge_7_left;
logic [5:0] index_ge_7_right;
logic index_ge_7_out;
logic idx_between_7_23_comb_left;
logic idx_between_7_23_comb_right;
logic idx_between_7_23_comb_out;
logic idx_between_22_23_reg_in;
logic idx_between_22_23_reg_write_en;
logic idx_between_22_23_reg_clk;
logic idx_between_22_23_reg_reset;
logic idx_between_22_23_reg_out;
logic idx_between_22_23_reg_done;
logic idx_between_22_23_comb_left;
logic idx_between_22_23_comb_right;
logic idx_between_22_23_comb_out;
logic idx_between_21_25_reg_in;
logic idx_between_21_25_reg_write_en;
logic idx_between_21_25_reg_clk;
logic idx_between_21_25_reg_reset;
logic idx_between_21_25_reg_out;
logic idx_between_21_25_reg_done;
logic [5:0] index_lt_25_left;
logic [5:0] index_lt_25_right;
logic index_lt_25_out;
logic idx_between_21_25_comb_left;
logic idx_between_21_25_comb_right;
logic idx_between_21_25_comb_out;
logic idx_between_3_19_reg_in;
logic idx_between_3_19_reg_write_en;
logic idx_between_3_19_reg_clk;
logic idx_between_3_19_reg_reset;
logic idx_between_3_19_reg_out;
logic idx_between_3_19_reg_done;
logic [5:0] index_lt_19_left;
logic [5:0] index_lt_19_right;
logic index_lt_19_out;
logic [5:0] index_ge_3_left;
logic [5:0] index_ge_3_right;
logic index_ge_3_out;
logic idx_between_3_19_comb_left;
logic idx_between_3_19_comb_right;
logic idx_between_3_19_comb_out;
logic idx_between_31_35_reg_in;
logic idx_between_31_35_reg_write_en;
logic idx_between_31_35_reg_clk;
logic idx_between_31_35_reg_reset;
logic idx_between_31_35_reg_out;
logic idx_between_31_35_reg_done;
logic [5:0] index_lt_35_left;
logic [5:0] index_lt_35_right;
logic index_lt_35_out;
logic idx_between_31_35_comb_left;
logic idx_between_31_35_comb_right;
logic idx_between_31_35_comb_out;
logic idx_between_49_50_reg_in;
logic idx_between_49_50_reg_write_en;
logic idx_between_49_50_reg_clk;
logic idx_between_49_50_reg_reset;
logic idx_between_49_50_reg_out;
logic idx_between_49_50_reg_done;
logic [5:0] index_lt_50_left;
logic [5:0] index_lt_50_right;
logic index_lt_50_out;
logic [5:0] index_ge_49_left;
logic [5:0] index_ge_49_right;
logic index_ge_49_out;
logic idx_between_49_50_comb_left;
logic idx_between_49_50_comb_right;
logic idx_between_49_50_comb_out;
logic idx_between_27_31_reg_in;
logic idx_between_27_31_reg_write_en;
logic idx_between_27_31_reg_clk;
logic idx_between_27_31_reg_reset;
logic idx_between_27_31_reg_out;
logic idx_between_27_31_reg_done;
logic [5:0] index_lt_31_left;
logic [5:0] index_lt_31_right;
logic index_lt_31_out;
logic idx_between_27_31_comb_left;
logic idx_between_27_31_comb_right;
logic idx_between_27_31_comb_out;
logic idx_between_45_46_reg_in;
logic idx_between_45_46_reg_write_en;
logic idx_between_45_46_reg_clk;
logic idx_between_45_46_reg_reset;
logic idx_between_45_46_reg_out;
logic idx_between_45_46_reg_done;
logic [5:0] index_ge_45_left;
logic [5:0] index_ge_45_right;
logic index_ge_45_out;
logic idx_between_45_46_comb_left;
logic idx_between_45_46_comb_right;
logic idx_between_45_46_comb_out;
logic idx_between_50_51_reg_in;
logic idx_between_50_51_reg_write_en;
logic idx_between_50_51_reg_clk;
logic idx_between_50_51_reg_reset;
logic idx_between_50_51_reg_out;
logic idx_between_50_51_reg_done;
logic [5:0] index_ge_50_left;
logic [5:0] index_ge_50_right;
logic index_ge_50_out;
logic idx_between_50_51_comb_left;
logic idx_between_50_51_comb_right;
logic idx_between_50_51_comb_out;
logic idx_between_51_52_reg_in;
logic idx_between_51_52_reg_write_en;
logic idx_between_51_52_reg_clk;
logic idx_between_51_52_reg_reset;
logic idx_between_51_52_reg_out;
logic idx_between_51_52_reg_done;
logic [5:0] index_lt_52_left;
logic [5:0] index_lt_52_right;
logic index_lt_52_out;
logic [5:0] index_ge_51_left;
logic [5:0] index_ge_51_right;
logic index_ge_51_out;
logic idx_between_51_52_comb_left;
logic idx_between_51_52_comb_right;
logic idx_between_51_52_comb_out;
logic idx_between_32_48_reg_in;
logic idx_between_32_48_reg_write_en;
logic idx_between_32_48_reg_clk;
logic idx_between_32_48_reg_reset;
logic idx_between_32_48_reg_out;
logic idx_between_32_48_reg_done;
logic [5:0] index_ge_32_left;
logic [5:0] index_ge_32_right;
logic index_ge_32_out;
logic idx_between_32_48_comb_left;
logic idx_between_32_48_comb_right;
logic idx_between_32_48_comb_out;
logic idx_between_5_9_reg_in;
logic idx_between_5_9_reg_write_en;
logic idx_between_5_9_reg_clk;
logic idx_between_5_9_reg_reset;
logic idx_between_5_9_reg_out;
logic idx_between_5_9_reg_done;
logic [5:0] index_lt_9_left;
logic [5:0] index_lt_9_right;
logic index_lt_9_out;
logic idx_between_5_9_comb_left;
logic idx_between_5_9_comb_right;
logic idx_between_5_9_comb_out;
logic idx_between_46_47_reg_in;
logic idx_between_46_47_reg_write_en;
logic idx_between_46_47_reg_clk;
logic idx_between_46_47_reg_reset;
logic idx_between_46_47_reg_out;
logic idx_between_46_47_reg_done;
logic [5:0] index_ge_46_left;
logic [5:0] index_ge_46_right;
logic index_ge_46_out;
logic idx_between_46_47_comb_left;
logic idx_between_46_47_comb_right;
logic idx_between_46_47_comb_out;
logic idx_between_23_24_reg_in;
logic idx_between_23_24_reg_write_en;
logic idx_between_23_24_reg_clk;
logic idx_between_23_24_reg_reset;
logic idx_between_23_24_reg_out;
logic idx_between_23_24_reg_done;
logic idx_between_23_24_comb_left;
logic idx_between_23_24_comb_right;
logic idx_between_23_24_comb_out;
logic idx_between_4_20_reg_in;
logic idx_between_4_20_reg_write_en;
logic idx_between_4_20_reg_clk;
logic idx_between_4_20_reg_reset;
logic idx_between_4_20_reg_out;
logic idx_between_4_20_reg_done;
logic [5:0] index_ge_4_left;
logic [5:0] index_ge_4_right;
logic index_ge_4_out;
logic idx_between_4_20_comb_left;
logic idx_between_4_20_comb_right;
logic idx_between_4_20_comb_out;
logic idx_between_14_30_reg_in;
logic idx_between_14_30_reg_write_en;
logic idx_between_14_30_reg_clk;
logic idx_between_14_30_reg_reset;
logic idx_between_14_30_reg_out;
logic idx_between_14_30_reg_done;
logic [5:0] index_ge_14_left;
logic [5:0] index_ge_14_right;
logic index_ge_14_out;
logic idx_between_14_30_comb_left;
logic idx_between_14_30_comb_right;
logic idx_between_14_30_comb_out;
logic idx_between_1_5_reg_in;
logic idx_between_1_5_reg_write_en;
logic idx_between_1_5_reg_clk;
logic idx_between_1_5_reg_reset;
logic idx_between_1_5_reg_out;
logic idx_between_1_5_reg_done;
logic [5:0] index_lt_5_left;
logic [5:0] index_lt_5_right;
logic index_lt_5_out;
logic idx_between_1_5_comb_left;
logic idx_between_1_5_comb_right;
logic idx_between_1_5_comb_out;
logic idx_between_28_32_reg_in;
logic idx_between_28_32_reg_write_en;
logic idx_between_28_32_reg_clk;
logic idx_between_28_32_reg_reset;
logic idx_between_28_32_reg_out;
logic idx_between_28_32_reg_done;
logic [5:0] index_lt_32_left;
logic [5:0] index_lt_32_right;
logic index_lt_32_out;
logic [5:0] index_ge_28_left;
logic [5:0] index_ge_28_right;
logic index_ge_28_out;
logic idx_between_28_32_comb_left;
logic idx_between_28_32_comb_right;
logic idx_between_28_32_comb_out;
logic idx_between_10_26_reg_in;
logic idx_between_10_26_reg_write_en;
logic idx_between_10_26_reg_clk;
logic idx_between_10_26_reg_reset;
logic idx_between_10_26_reg_out;
logic idx_between_10_26_reg_done;
logic [5:0] index_ge_10_left;
logic [5:0] index_ge_10_right;
logic index_ge_10_out;
logic idx_between_10_26_comb_left;
logic idx_between_10_26_comb_right;
logic idx_between_10_26_comb_out;
logic idx_between_24_25_reg_in;
logic idx_between_24_25_reg_write_en;
logic idx_between_24_25_reg_clk;
logic idx_between_24_25_reg_reset;
logic idx_between_24_25_reg_out;
logic idx_between_24_25_reg_done;
logic idx_between_24_25_comb_left;
logic idx_between_24_25_comb_right;
logic idx_between_24_25_comb_out;
logic idx_between_6_22_reg_in;
logic idx_between_6_22_reg_write_en;
logic idx_between_6_22_reg_clk;
logic idx_between_6_22_reg_reset;
logic idx_between_6_22_reg_out;
logic idx_between_6_22_reg_done;
logic [5:0] index_lt_22_left;
logic [5:0] index_lt_22_right;
logic index_lt_22_out;
logic [5:0] index_ge_6_left;
logic [5:0] index_ge_6_right;
logic index_ge_6_out;
logic idx_between_6_22_comb_left;
logic idx_between_6_22_comb_right;
logic idx_between_6_22_comb_out;
logic idx_between_29_33_reg_in;
logic idx_between_29_33_reg_write_en;
logic idx_between_29_33_reg_clk;
logic idx_between_29_33_reg_reset;
logic idx_between_29_33_reg_out;
logic idx_between_29_33_reg_done;
logic [5:0] index_lt_33_left;
logic [5:0] index_lt_33_right;
logic index_lt_33_out;
logic idx_between_29_33_comb_left;
logic idx_between_29_33_comb_right;
logic idx_between_29_33_comb_out;
logic idx_between_2_6_reg_in;
logic idx_between_2_6_reg_write_en;
logic idx_between_2_6_reg_clk;
logic idx_between_2_6_reg_reset;
logic idx_between_2_6_reg_out;
logic idx_between_2_6_reg_done;
logic [5:0] index_lt_6_left;
logic [5:0] index_lt_6_right;
logic index_lt_6_out;
logic [5:0] index_ge_2_left;
logic [5:0] index_ge_2_right;
logic index_ge_2_out;
logic idx_between_2_6_comb_left;
logic idx_between_2_6_comb_right;
logic idx_between_2_6_comb_out;
logic idx_between_30_31_reg_in;
logic idx_between_30_31_reg_write_en;
logic idx_between_30_31_reg_clk;
logic idx_between_30_31_reg_reset;
logic idx_between_30_31_reg_out;
logic idx_between_30_31_reg_done;
logic idx_between_30_31_comb_left;
logic idx_between_30_31_comb_right;
logic idx_between_30_31_comb_out;
logic idx_between_34_50_reg_in;
logic idx_between_34_50_reg_write_en;
logic idx_between_34_50_reg_clk;
logic idx_between_34_50_reg_reset;
logic idx_between_34_50_reg_out;
logic idx_between_34_50_reg_done;
logic [5:0] index_ge_34_left;
logic [5:0] index_ge_34_right;
logic index_ge_34_out;
logic idx_between_34_50_comb_left;
logic idx_between_34_50_comb_right;
logic idx_between_34_50_comb_out;
logic idx_between_7_11_reg_in;
logic idx_between_7_11_reg_write_en;
logic idx_between_7_11_reg_clk;
logic idx_between_7_11_reg_reset;
logic idx_between_7_11_reg_out;
logic idx_between_7_11_reg_done;
logic [5:0] index_lt_11_left;
logic [5:0] index_lt_11_right;
logic index_lt_11_out;
logic idx_between_7_11_comb_left;
logic idx_between_7_11_comb_right;
logic idx_between_7_11_comb_out;
logic idx_between_11_27_reg_in;
logic idx_between_11_27_reg_write_en;
logic idx_between_11_27_reg_clk;
logic idx_between_11_27_reg_reset;
logic idx_between_11_27_reg_out;
logic idx_between_11_27_reg_done;
logic [5:0] index_ge_11_left;
logic [5:0] index_ge_11_right;
logic index_ge_11_out;
logic idx_between_11_27_comb_left;
logic idx_between_11_27_comb_right;
logic idx_between_11_27_comb_out;
logic idx_between_25_26_reg_in;
logic idx_between_25_26_reg_write_en;
logic idx_between_25_26_reg_clk;
logic idx_between_25_26_reg_reset;
logic idx_between_25_26_reg_out;
logic idx_between_25_26_reg_done;
logic idx_between_25_26_comb_left;
logic idx_between_25_26_comb_right;
logic idx_between_25_26_comb_out;
logic idx_between_26_27_reg_in;
logic idx_between_26_27_reg_write_en;
logic idx_between_26_27_reg_clk;
logic idx_between_26_27_reg_reset;
logic idx_between_26_27_reg_out;
logic idx_between_26_27_reg_done;
logic idx_between_26_27_comb_left;
logic idx_between_26_27_comb_right;
logic idx_between_26_27_comb_out;
logic idx_between_3_7_reg_in;
logic idx_between_3_7_reg_write_en;
logic idx_between_3_7_reg_clk;
logic idx_between_3_7_reg_reset;
logic idx_between_3_7_reg_out;
logic idx_between_3_7_reg_done;
logic [5:0] index_lt_7_left;
logic [5:0] index_lt_7_right;
logic index_lt_7_out;
logic idx_between_3_7_comb_left;
logic idx_between_3_7_comb_right;
logic idx_between_3_7_comb_out;
logic idx_between_21_22_reg_in;
logic idx_between_21_22_reg_write_en;
logic idx_between_21_22_reg_clk;
logic idx_between_21_22_reg_reset;
logic idx_between_21_22_reg_out;
logic idx_between_21_22_reg_done;
logic idx_between_21_22_comb_left;
logic idx_between_21_22_comb_right;
logic idx_between_21_22_comb_out;
logic idx_between_31_32_reg_in;
logic idx_between_31_32_reg_write_en;
logic idx_between_31_32_reg_clk;
logic idx_between_31_32_reg_reset;
logic idx_between_31_32_reg_out;
logic idx_between_31_32_reg_done;
logic idx_between_31_32_comb_left;
logic idx_between_31_32_comb_right;
logic idx_between_31_32_comb_out;
logic idx_between_12_28_reg_in;
logic idx_between_12_28_reg_write_en;
logic idx_between_12_28_reg_clk;
logic idx_between_12_28_reg_reset;
logic idx_between_12_28_reg_out;
logic idx_between_12_28_reg_done;
logic [5:0] index_ge_12_left;
logic [5:0] index_ge_12_right;
logic index_ge_12_out;
logic idx_between_12_28_comb_left;
logic idx_between_12_28_comb_right;
logic idx_between_12_28_comb_out;
logic idx_between_27_28_reg_in;
logic idx_between_27_28_reg_write_en;
logic idx_between_27_28_reg_clk;
logic idx_between_27_28_reg_reset;
logic idx_between_27_28_reg_out;
logic idx_between_27_28_reg_done;
logic idx_between_27_28_comb_left;
logic idx_between_27_28_comb_right;
logic idx_between_27_28_comb_out;
logic idx_between_8_24_reg_in;
logic idx_between_8_24_reg_write_en;
logic idx_between_8_24_reg_clk;
logic idx_between_8_24_reg_reset;
logic idx_between_8_24_reg_out;
logic idx_between_8_24_reg_done;
logic [5:0] index_ge_8_left;
logic [5:0] index_ge_8_right;
logic index_ge_8_out;
logic idx_between_8_24_comb_left;
logic idx_between_8_24_comb_right;
logic idx_between_8_24_comb_out;
logic idx_between_4_8_reg_in;
logic idx_between_4_8_reg_write_en;
logic idx_between_4_8_reg_clk;
logic idx_between_4_8_reg_reset;
logic idx_between_4_8_reg_out;
logic idx_between_4_8_reg_done;
logic [5:0] index_lt_8_left;
logic [5:0] index_lt_8_right;
logic index_lt_8_out;
logic idx_between_4_8_comb_left;
logic idx_between_4_8_comb_right;
logic idx_between_4_8_comb_out;
logic idx_between_14_18_reg_in;
logic idx_between_14_18_reg_write_en;
logic idx_between_14_18_reg_clk;
logic idx_between_14_18_reg_reset;
logic idx_between_14_18_reg_out;
logic idx_between_14_18_reg_done;
logic [5:0] index_lt_18_left;
logic [5:0] index_lt_18_right;
logic index_lt_18_out;
logic idx_between_14_18_comb_left;
logic idx_between_14_18_comb_right;
logic idx_between_14_18_comb_out;
logic idx_between_18_34_reg_in;
logic idx_between_18_34_reg_write_en;
logic idx_between_18_34_reg_clk;
logic idx_between_18_34_reg_reset;
logic idx_between_18_34_reg_out;
logic idx_between_18_34_reg_done;
logic [5:0] index_ge_18_left;
logic [5:0] index_ge_18_right;
logic index_ge_18_out;
logic idx_between_18_34_comb_left;
logic idx_between_18_34_comb_right;
logic idx_between_18_34_comb_out;
logic idx_between_10_14_reg_in;
logic idx_between_10_14_reg_write_en;
logic idx_between_10_14_reg_clk;
logic idx_between_10_14_reg_reset;
logic idx_between_10_14_reg_out;
logic idx_between_10_14_reg_done;
logic [5:0] index_lt_14_left;
logic [5:0] index_lt_14_right;
logic index_lt_14_out;
logic idx_between_10_14_comb_left;
logic idx_between_10_14_comb_right;
logic idx_between_10_14_comb_out;
logic idx_between_28_29_reg_in;
logic idx_between_28_29_reg_write_en;
logic idx_between_28_29_reg_clk;
logic idx_between_28_29_reg_reset;
logic idx_between_28_29_reg_out;
logic idx_between_28_29_reg_done;
logic idx_between_28_29_comb_left;
logic idx_between_28_29_comb_right;
logic idx_between_28_29_comb_out;
logic idx_between_9_25_reg_in;
logic idx_between_9_25_reg_write_en;
logic idx_between_9_25_reg_clk;
logic idx_between_9_25_reg_reset;
logic idx_between_9_25_reg_out;
logic idx_between_9_25_reg_done;
logic [5:0] index_ge_9_left;
logic [5:0] index_ge_9_right;
logic index_ge_9_out;
logic idx_between_9_25_comb_left;
logic idx_between_9_25_comb_right;
logic idx_between_9_25_comb_out;
logic idx_between_19_35_reg_in;
logic idx_between_19_35_reg_write_en;
logic idx_between_19_35_reg_clk;
logic idx_between_19_35_reg_reset;
logic idx_between_19_35_reg_out;
logic idx_between_19_35_reg_done;
logic [5:0] index_ge_19_left;
logic [5:0] index_ge_19_right;
logic index_ge_19_out;
logic idx_between_19_35_comb_left;
logic idx_between_19_35_comb_right;
logic idx_between_19_35_comb_out;
logic idx_between_6_10_reg_in;
logic idx_between_6_10_reg_write_en;
logic idx_between_6_10_reg_clk;
logic idx_between_6_10_reg_reset;
logic idx_between_6_10_reg_out;
logic idx_between_6_10_reg_done;
logic [5:0] index_lt_10_left;
logic [5:0] index_lt_10_right;
logic index_lt_10_out;
logic idx_between_6_10_comb_left;
logic idx_between_6_10_comb_right;
logic idx_between_6_10_comb_out;
logic idx_between_15_31_reg_in;
logic idx_between_15_31_reg_write_en;
logic idx_between_15_31_reg_clk;
logic idx_between_15_31_reg_reset;
logic idx_between_15_31_reg_out;
logic idx_between_15_31_reg_done;
logic [5:0] index_ge_15_left;
logic [5:0] index_ge_15_right;
logic index_ge_15_out;
logic idx_between_15_31_comb_left;
logic idx_between_15_31_comb_right;
logic idx_between_15_31_comb_out;
logic idx_between_29_30_reg_in;
logic idx_between_29_30_reg_write_en;
logic idx_between_29_30_reg_clk;
logic idx_between_29_30_reg_reset;
logic idx_between_29_30_reg_out;
logic idx_between_29_30_reg_done;
logic idx_between_29_30_comb_left;
logic idx_between_29_30_comb_right;
logic idx_between_29_30_comb_out;
logic idx_between_11_15_reg_in;
logic idx_between_11_15_reg_write_en;
logic idx_between_11_15_reg_clk;
logic idx_between_11_15_reg_reset;
logic idx_between_11_15_reg_out;
logic idx_between_11_15_reg_done;
logic [5:0] index_lt_15_left;
logic [5:0] index_lt_15_right;
logic index_lt_15_out;
logic idx_between_11_15_comb_left;
logic idx_between_11_15_comb_right;
logic idx_between_11_15_comb_out;
logic idx_between_35_36_reg_in;
logic idx_between_35_36_reg_write_en;
logic idx_between_35_36_reg_clk;
logic idx_between_35_36_reg_reset;
logic idx_between_35_36_reg_out;
logic idx_between_35_36_reg_done;
logic [5:0] index_lt_36_left;
logic [5:0] index_lt_36_right;
logic index_lt_36_out;
logic idx_between_35_36_comb_left;
logic idx_between_35_36_comb_right;
logic idx_between_35_36_comb_out;
logic idx_between_12_16_reg_in;
logic idx_between_12_16_reg_write_en;
logic idx_between_12_16_reg_clk;
logic idx_between_12_16_reg_reset;
logic idx_between_12_16_reg_out;
logic idx_between_12_16_reg_done;
logic idx_between_12_16_comb_left;
logic idx_between_12_16_comb_right;
logic idx_between_12_16_comb_out;
logic idx_between_16_32_reg_in;
logic idx_between_16_32_reg_write_en;
logic idx_between_16_32_reg_clk;
logic idx_between_16_32_reg_reset;
logic idx_between_16_32_reg_out;
logic idx_between_16_32_reg_done;
logic idx_between_16_32_comb_left;
logic idx_between_16_32_comb_right;
logic idx_between_16_32_comb_out;
logic idx_between_26_42_reg_in;
logic idx_between_26_42_reg_write_en;
logic idx_between_26_42_reg_clk;
logic idx_between_26_42_reg_reset;
logic idx_between_26_42_reg_out;
logic idx_between_26_42_reg_done;
logic idx_between_26_42_comb_left;
logic idx_between_26_42_comb_right;
logic idx_between_26_42_comb_out;
logic idx_between_8_12_reg_in;
logic idx_between_8_12_reg_write_en;
logic idx_between_8_12_reg_clk;
logic idx_between_8_12_reg_reset;
logic idx_between_8_12_reg_out;
logic idx_between_8_12_reg_done;
logic [5:0] index_lt_12_left;
logic [5:0] index_lt_12_right;
logic index_lt_12_out;
logic idx_between_8_12_comb_left;
logic idx_between_8_12_comb_right;
logic idx_between_8_12_comb_out;
logic idx_between_22_38_reg_in;
logic idx_between_22_38_reg_write_en;
logic idx_between_22_38_reg_clk;
logic idx_between_22_38_reg_reset;
logic idx_between_22_38_reg_out;
logic idx_between_22_38_reg_done;
logic [5:0] index_lt_38_left;
logic [5:0] index_lt_38_right;
logic index_lt_38_out;
logic idx_between_22_38_comb_left;
logic idx_between_22_38_comb_right;
logic idx_between_22_38_comb_out;
logic idx_between_36_37_reg_in;
logic idx_between_36_37_reg_write_en;
logic idx_between_36_37_reg_clk;
logic idx_between_36_37_reg_reset;
logic idx_between_36_37_reg_out;
logic idx_between_36_37_reg_done;
logic [5:0] index_ge_36_left;
logic [5:0] index_ge_36_right;
logic index_ge_36_out;
logic idx_between_36_37_comb_left;
logic idx_between_36_37_comb_right;
logic idx_between_36_37_comb_out;
logic idx_between_17_33_reg_in;
logic idx_between_17_33_reg_write_en;
logic idx_between_17_33_reg_clk;
logic idx_between_17_33_reg_reset;
logic idx_between_17_33_reg_out;
logic idx_between_17_33_reg_done;
logic idx_between_17_33_comb_left;
logic idx_between_17_33_comb_right;
logic idx_between_17_33_comb_out;
logic idx_between_32_33_reg_in;
logic idx_between_32_33_reg_write_en;
logic idx_between_32_33_reg_clk;
logic idx_between_32_33_reg_reset;
logic idx_between_32_33_reg_out;
logic idx_between_32_33_reg_done;
logic idx_between_32_33_comb_left;
logic idx_between_32_33_comb_right;
logic idx_between_32_33_comb_out;
logic idx_between_13_29_reg_in;
logic idx_between_13_29_reg_write_en;
logic idx_between_13_29_reg_clk;
logic idx_between_13_29_reg_reset;
logic idx_between_13_29_reg_out;
logic idx_between_13_29_reg_done;
logic idx_between_13_29_comb_left;
logic idx_between_13_29_comb_right;
logic idx_between_13_29_comb_out;
logic idx_between_18_22_reg_in;
logic idx_between_18_22_reg_write_en;
logic idx_between_18_22_reg_clk;
logic idx_between_18_22_reg_reset;
logic idx_between_18_22_reg_out;
logic idx_between_18_22_reg_done;
logic idx_between_18_22_comb_left;
logic idx_between_18_22_comb_right;
logic idx_between_18_22_comb_out;
logic idx_between_9_13_reg_in;
logic idx_between_9_13_reg_write_en;
logic idx_between_9_13_reg_clk;
logic idx_between_9_13_reg_reset;
logic idx_between_9_13_reg_out;
logic idx_between_9_13_reg_done;
logic [5:0] index_lt_13_left;
logic [5:0] index_lt_13_right;
logic index_lt_13_out;
logic idx_between_9_13_comb_left;
logic idx_between_9_13_comb_right;
logic idx_between_9_13_comb_out;
logic idx_between_19_23_reg_in;
logic idx_between_19_23_reg_write_en;
logic idx_between_19_23_reg_clk;
logic idx_between_19_23_reg_reset;
logic idx_between_19_23_reg_out;
logic idx_between_19_23_reg_done;
logic idx_between_19_23_comb_left;
logic idx_between_19_23_comb_right;
logic idx_between_19_23_comb_out;
logic idx_between_23_39_reg_in;
logic idx_between_23_39_reg_write_en;
logic idx_between_23_39_reg_clk;
logic idx_between_23_39_reg_reset;
logic idx_between_23_39_reg_out;
logic idx_between_23_39_reg_done;
logic idx_between_23_39_comb_left;
logic idx_between_23_39_comb_right;
logic idx_between_23_39_comb_out;
logic idx_between_37_38_reg_in;
logic idx_between_37_38_reg_write_en;
logic idx_between_37_38_reg_clk;
logic idx_between_37_38_reg_reset;
logic idx_between_37_38_reg_out;
logic idx_between_37_38_reg_done;
logic [5:0] index_ge_37_left;
logic [5:0] index_ge_37_right;
logic index_ge_37_out;
logic idx_between_37_38_comb_left;
logic idx_between_37_38_comb_right;
logic idx_between_37_38_comb_out;
logic idx_between_28_44_reg_in;
logic idx_between_28_44_reg_write_en;
logic idx_between_28_44_reg_clk;
logic idx_between_28_44_reg_reset;
logic idx_between_28_44_reg_out;
logic idx_between_28_44_reg_done;
logic [5:0] index_lt_44_left;
logic [5:0] index_lt_44_right;
logic index_lt_44_out;
logic idx_between_28_44_comb_left;
logic idx_between_28_44_comb_right;
logic idx_between_28_44_comb_out;
logic idx_between_15_19_reg_in;
logic idx_between_15_19_reg_write_en;
logic idx_between_15_19_reg_clk;
logic idx_between_15_19_reg_reset;
logic idx_between_15_19_reg_out;
logic idx_between_15_19_reg_done;
logic idx_between_15_19_comb_left;
logic idx_between_15_19_comb_right;
logic idx_between_15_19_comb_out;
logic idx_between_33_34_reg_in;
logic idx_between_33_34_reg_write_en;
logic idx_between_33_34_reg_clk;
logic idx_between_33_34_reg_reset;
logic idx_between_33_34_reg_out;
logic idx_between_33_34_reg_done;
logic idx_between_33_34_comb_left;
logic idx_between_33_34_comb_right;
logic idx_between_33_34_comb_out;
logic idx_between_43_44_reg_in;
logic idx_between_43_44_reg_write_en;
logic idx_between_43_44_reg_clk;
logic idx_between_43_44_reg_reset;
logic idx_between_43_44_reg_out;
logic idx_between_43_44_reg_done;
logic [5:0] index_ge_43_left;
logic [5:0] index_ge_43_right;
logic index_ge_43_out;
logic idx_between_43_44_comb_left;
logic idx_between_43_44_comb_right;
logic idx_between_43_44_comb_out;
logic idx_between_24_40_reg_in;
logic idx_between_24_40_reg_write_en;
logic idx_between_24_40_reg_clk;
logic idx_between_24_40_reg_reset;
logic idx_between_24_40_reg_out;
logic idx_between_24_40_reg_done;
logic [5:0] index_lt_40_left;
logic [5:0] index_lt_40_right;
logic index_lt_40_out;
logic idx_between_24_40_comb_left;
logic idx_between_24_40_comb_right;
logic idx_between_24_40_comb_out;
logic idx_between_39_40_reg_in;
logic idx_between_39_40_reg_write_en;
logic idx_between_39_40_reg_clk;
logic idx_between_39_40_reg_reset;
logic idx_between_39_40_reg_out;
logic idx_between_39_40_reg_done;
logic [5:0] index_ge_39_left;
logic [5:0] index_ge_39_right;
logic index_ge_39_out;
logic idx_between_39_40_comb_left;
logic idx_between_39_40_comb_right;
logic idx_between_39_40_comb_out;
logic idx_between_20_36_reg_in;
logic idx_between_20_36_reg_write_en;
logic idx_between_20_36_reg_clk;
logic idx_between_20_36_reg_reset;
logic idx_between_20_36_reg_out;
logic idx_between_20_36_reg_done;
logic idx_between_20_36_comb_left;
logic idx_between_20_36_comb_right;
logic idx_between_20_36_comb_out;
logic idx_between_34_35_reg_in;
logic idx_between_34_35_reg_write_en;
logic idx_between_34_35_reg_clk;
logic idx_between_34_35_reg_reset;
logic idx_between_34_35_reg_out;
logic idx_between_34_35_reg_done;
logic idx_between_34_35_comb_left;
logic idx_between_34_35_comb_right;
logic idx_between_34_35_comb_out;
logic idx_between_2_18_reg_in;
logic idx_between_2_18_reg_write_en;
logic idx_between_2_18_reg_clk;
logic idx_between_2_18_reg_reset;
logic idx_between_2_18_reg_out;
logic idx_between_2_18_reg_done;
logic idx_between_2_18_comb_left;
logic idx_between_2_18_comb_right;
logic idx_between_2_18_comb_out;
logic cond_in;
logic cond_write_en;
logic cond_clk;
logic cond_reset;
logic cond_out;
logic cond_done;
logic cond_wire_in;
logic cond_wire_out;
logic cond0_in;
logic cond0_write_en;
logic cond0_clk;
logic cond0_reset;
logic cond0_out;
logic cond0_done;
logic cond_wire0_in;
logic cond_wire0_out;
logic cond1_in;
logic cond1_write_en;
logic cond1_clk;
logic cond1_reset;
logic cond1_out;
logic cond1_done;
logic cond_wire1_in;
logic cond_wire1_out;
logic cond2_in;
logic cond2_write_en;
logic cond2_clk;
logic cond2_reset;
logic cond2_out;
logic cond2_done;
logic cond_wire2_in;
logic cond_wire2_out;
logic cond3_in;
logic cond3_write_en;
logic cond3_clk;
logic cond3_reset;
logic cond3_out;
logic cond3_done;
logic cond_wire3_in;
logic cond_wire3_out;
logic cond4_in;
logic cond4_write_en;
logic cond4_clk;
logic cond4_reset;
logic cond4_out;
logic cond4_done;
logic cond_wire4_in;
logic cond_wire4_out;
logic cond5_in;
logic cond5_write_en;
logic cond5_clk;
logic cond5_reset;
logic cond5_out;
logic cond5_done;
logic cond_wire5_in;
logic cond_wire5_out;
logic cond6_in;
logic cond6_write_en;
logic cond6_clk;
logic cond6_reset;
logic cond6_out;
logic cond6_done;
logic cond_wire6_in;
logic cond_wire6_out;
logic cond7_in;
logic cond7_write_en;
logic cond7_clk;
logic cond7_reset;
logic cond7_out;
logic cond7_done;
logic cond_wire7_in;
logic cond_wire7_out;
logic cond8_in;
logic cond8_write_en;
logic cond8_clk;
logic cond8_reset;
logic cond8_out;
logic cond8_done;
logic cond_wire8_in;
logic cond_wire8_out;
logic cond9_in;
logic cond9_write_en;
logic cond9_clk;
logic cond9_reset;
logic cond9_out;
logic cond9_done;
logic cond_wire9_in;
logic cond_wire9_out;
logic cond10_in;
logic cond10_write_en;
logic cond10_clk;
logic cond10_reset;
logic cond10_out;
logic cond10_done;
logic cond_wire10_in;
logic cond_wire10_out;
logic cond11_in;
logic cond11_write_en;
logic cond11_clk;
logic cond11_reset;
logic cond11_out;
logic cond11_done;
logic cond_wire11_in;
logic cond_wire11_out;
logic cond12_in;
logic cond12_write_en;
logic cond12_clk;
logic cond12_reset;
logic cond12_out;
logic cond12_done;
logic cond_wire12_in;
logic cond_wire12_out;
logic cond13_in;
logic cond13_write_en;
logic cond13_clk;
logic cond13_reset;
logic cond13_out;
logic cond13_done;
logic cond_wire13_in;
logic cond_wire13_out;
logic cond14_in;
logic cond14_write_en;
logic cond14_clk;
logic cond14_reset;
logic cond14_out;
logic cond14_done;
logic cond_wire14_in;
logic cond_wire14_out;
logic cond15_in;
logic cond15_write_en;
logic cond15_clk;
logic cond15_reset;
logic cond15_out;
logic cond15_done;
logic cond_wire15_in;
logic cond_wire15_out;
logic cond16_in;
logic cond16_write_en;
logic cond16_clk;
logic cond16_reset;
logic cond16_out;
logic cond16_done;
logic cond_wire16_in;
logic cond_wire16_out;
logic cond17_in;
logic cond17_write_en;
logic cond17_clk;
logic cond17_reset;
logic cond17_out;
logic cond17_done;
logic cond_wire17_in;
logic cond_wire17_out;
logic cond18_in;
logic cond18_write_en;
logic cond18_clk;
logic cond18_reset;
logic cond18_out;
logic cond18_done;
logic cond_wire18_in;
logic cond_wire18_out;
logic cond19_in;
logic cond19_write_en;
logic cond19_clk;
logic cond19_reset;
logic cond19_out;
logic cond19_done;
logic cond_wire19_in;
logic cond_wire19_out;
logic cond20_in;
logic cond20_write_en;
logic cond20_clk;
logic cond20_reset;
logic cond20_out;
logic cond20_done;
logic cond_wire20_in;
logic cond_wire20_out;
logic cond21_in;
logic cond21_write_en;
logic cond21_clk;
logic cond21_reset;
logic cond21_out;
logic cond21_done;
logic cond_wire21_in;
logic cond_wire21_out;
logic cond22_in;
logic cond22_write_en;
logic cond22_clk;
logic cond22_reset;
logic cond22_out;
logic cond22_done;
logic cond_wire22_in;
logic cond_wire22_out;
logic cond23_in;
logic cond23_write_en;
logic cond23_clk;
logic cond23_reset;
logic cond23_out;
logic cond23_done;
logic cond_wire23_in;
logic cond_wire23_out;
logic cond24_in;
logic cond24_write_en;
logic cond24_clk;
logic cond24_reset;
logic cond24_out;
logic cond24_done;
logic cond_wire24_in;
logic cond_wire24_out;
logic cond25_in;
logic cond25_write_en;
logic cond25_clk;
logic cond25_reset;
logic cond25_out;
logic cond25_done;
logic cond_wire25_in;
logic cond_wire25_out;
logic cond26_in;
logic cond26_write_en;
logic cond26_clk;
logic cond26_reset;
logic cond26_out;
logic cond26_done;
logic cond_wire26_in;
logic cond_wire26_out;
logic cond27_in;
logic cond27_write_en;
logic cond27_clk;
logic cond27_reset;
logic cond27_out;
logic cond27_done;
logic cond_wire27_in;
logic cond_wire27_out;
logic cond28_in;
logic cond28_write_en;
logic cond28_clk;
logic cond28_reset;
logic cond28_out;
logic cond28_done;
logic cond_wire28_in;
logic cond_wire28_out;
logic cond29_in;
logic cond29_write_en;
logic cond29_clk;
logic cond29_reset;
logic cond29_out;
logic cond29_done;
logic cond_wire29_in;
logic cond_wire29_out;
logic cond30_in;
logic cond30_write_en;
logic cond30_clk;
logic cond30_reset;
logic cond30_out;
logic cond30_done;
logic cond_wire30_in;
logic cond_wire30_out;
logic cond31_in;
logic cond31_write_en;
logic cond31_clk;
logic cond31_reset;
logic cond31_out;
logic cond31_done;
logic cond_wire31_in;
logic cond_wire31_out;
logic cond32_in;
logic cond32_write_en;
logic cond32_clk;
logic cond32_reset;
logic cond32_out;
logic cond32_done;
logic cond_wire32_in;
logic cond_wire32_out;
logic cond33_in;
logic cond33_write_en;
logic cond33_clk;
logic cond33_reset;
logic cond33_out;
logic cond33_done;
logic cond_wire33_in;
logic cond_wire33_out;
logic cond34_in;
logic cond34_write_en;
logic cond34_clk;
logic cond34_reset;
logic cond34_out;
logic cond34_done;
logic cond_wire34_in;
logic cond_wire34_out;
logic cond35_in;
logic cond35_write_en;
logic cond35_clk;
logic cond35_reset;
logic cond35_out;
logic cond35_done;
logic cond_wire35_in;
logic cond_wire35_out;
logic cond36_in;
logic cond36_write_en;
logic cond36_clk;
logic cond36_reset;
logic cond36_out;
logic cond36_done;
logic cond_wire36_in;
logic cond_wire36_out;
logic cond37_in;
logic cond37_write_en;
logic cond37_clk;
logic cond37_reset;
logic cond37_out;
logic cond37_done;
logic cond_wire37_in;
logic cond_wire37_out;
logic cond38_in;
logic cond38_write_en;
logic cond38_clk;
logic cond38_reset;
logic cond38_out;
logic cond38_done;
logic cond_wire38_in;
logic cond_wire38_out;
logic cond39_in;
logic cond39_write_en;
logic cond39_clk;
logic cond39_reset;
logic cond39_out;
logic cond39_done;
logic cond_wire39_in;
logic cond_wire39_out;
logic cond40_in;
logic cond40_write_en;
logic cond40_clk;
logic cond40_reset;
logic cond40_out;
logic cond40_done;
logic cond_wire40_in;
logic cond_wire40_out;
logic cond41_in;
logic cond41_write_en;
logic cond41_clk;
logic cond41_reset;
logic cond41_out;
logic cond41_done;
logic cond_wire41_in;
logic cond_wire41_out;
logic cond42_in;
logic cond42_write_en;
logic cond42_clk;
logic cond42_reset;
logic cond42_out;
logic cond42_done;
logic cond_wire42_in;
logic cond_wire42_out;
logic cond43_in;
logic cond43_write_en;
logic cond43_clk;
logic cond43_reset;
logic cond43_out;
logic cond43_done;
logic cond_wire43_in;
logic cond_wire43_out;
logic cond44_in;
logic cond44_write_en;
logic cond44_clk;
logic cond44_reset;
logic cond44_out;
logic cond44_done;
logic cond_wire44_in;
logic cond_wire44_out;
logic cond45_in;
logic cond45_write_en;
logic cond45_clk;
logic cond45_reset;
logic cond45_out;
logic cond45_done;
logic cond_wire45_in;
logic cond_wire45_out;
logic cond46_in;
logic cond46_write_en;
logic cond46_clk;
logic cond46_reset;
logic cond46_out;
logic cond46_done;
logic cond_wire46_in;
logic cond_wire46_out;
logic cond47_in;
logic cond47_write_en;
logic cond47_clk;
logic cond47_reset;
logic cond47_out;
logic cond47_done;
logic cond_wire47_in;
logic cond_wire47_out;
logic cond48_in;
logic cond48_write_en;
logic cond48_clk;
logic cond48_reset;
logic cond48_out;
logic cond48_done;
logic cond_wire48_in;
logic cond_wire48_out;
logic cond49_in;
logic cond49_write_en;
logic cond49_clk;
logic cond49_reset;
logic cond49_out;
logic cond49_done;
logic cond_wire49_in;
logic cond_wire49_out;
logic cond50_in;
logic cond50_write_en;
logic cond50_clk;
logic cond50_reset;
logic cond50_out;
logic cond50_done;
logic cond_wire50_in;
logic cond_wire50_out;
logic cond51_in;
logic cond51_write_en;
logic cond51_clk;
logic cond51_reset;
logic cond51_out;
logic cond51_done;
logic cond_wire51_in;
logic cond_wire51_out;
logic cond52_in;
logic cond52_write_en;
logic cond52_clk;
logic cond52_reset;
logic cond52_out;
logic cond52_done;
logic cond_wire52_in;
logic cond_wire52_out;
logic cond53_in;
logic cond53_write_en;
logic cond53_clk;
logic cond53_reset;
logic cond53_out;
logic cond53_done;
logic cond_wire53_in;
logic cond_wire53_out;
logic cond54_in;
logic cond54_write_en;
logic cond54_clk;
logic cond54_reset;
logic cond54_out;
logic cond54_done;
logic cond_wire54_in;
logic cond_wire54_out;
logic cond55_in;
logic cond55_write_en;
logic cond55_clk;
logic cond55_reset;
logic cond55_out;
logic cond55_done;
logic cond_wire55_in;
logic cond_wire55_out;
logic cond56_in;
logic cond56_write_en;
logic cond56_clk;
logic cond56_reset;
logic cond56_out;
logic cond56_done;
logic cond_wire56_in;
logic cond_wire56_out;
logic cond57_in;
logic cond57_write_en;
logic cond57_clk;
logic cond57_reset;
logic cond57_out;
logic cond57_done;
logic cond_wire57_in;
logic cond_wire57_out;
logic cond58_in;
logic cond58_write_en;
logic cond58_clk;
logic cond58_reset;
logic cond58_out;
logic cond58_done;
logic cond_wire58_in;
logic cond_wire58_out;
logic cond59_in;
logic cond59_write_en;
logic cond59_clk;
logic cond59_reset;
logic cond59_out;
logic cond59_done;
logic cond_wire59_in;
logic cond_wire59_out;
logic cond60_in;
logic cond60_write_en;
logic cond60_clk;
logic cond60_reset;
logic cond60_out;
logic cond60_done;
logic cond_wire60_in;
logic cond_wire60_out;
logic cond61_in;
logic cond61_write_en;
logic cond61_clk;
logic cond61_reset;
logic cond61_out;
logic cond61_done;
logic cond_wire61_in;
logic cond_wire61_out;
logic cond62_in;
logic cond62_write_en;
logic cond62_clk;
logic cond62_reset;
logic cond62_out;
logic cond62_done;
logic cond_wire62_in;
logic cond_wire62_out;
logic cond63_in;
logic cond63_write_en;
logic cond63_clk;
logic cond63_reset;
logic cond63_out;
logic cond63_done;
logic cond_wire63_in;
logic cond_wire63_out;
logic cond64_in;
logic cond64_write_en;
logic cond64_clk;
logic cond64_reset;
logic cond64_out;
logic cond64_done;
logic cond_wire64_in;
logic cond_wire64_out;
logic cond65_in;
logic cond65_write_en;
logic cond65_clk;
logic cond65_reset;
logic cond65_out;
logic cond65_done;
logic cond_wire65_in;
logic cond_wire65_out;
logic cond66_in;
logic cond66_write_en;
logic cond66_clk;
logic cond66_reset;
logic cond66_out;
logic cond66_done;
logic cond_wire66_in;
logic cond_wire66_out;
logic cond67_in;
logic cond67_write_en;
logic cond67_clk;
logic cond67_reset;
logic cond67_out;
logic cond67_done;
logic cond_wire67_in;
logic cond_wire67_out;
logic cond68_in;
logic cond68_write_en;
logic cond68_clk;
logic cond68_reset;
logic cond68_out;
logic cond68_done;
logic cond_wire68_in;
logic cond_wire68_out;
logic cond69_in;
logic cond69_write_en;
logic cond69_clk;
logic cond69_reset;
logic cond69_out;
logic cond69_done;
logic cond_wire69_in;
logic cond_wire69_out;
logic cond70_in;
logic cond70_write_en;
logic cond70_clk;
logic cond70_reset;
logic cond70_out;
logic cond70_done;
logic cond_wire70_in;
logic cond_wire70_out;
logic cond71_in;
logic cond71_write_en;
logic cond71_clk;
logic cond71_reset;
logic cond71_out;
logic cond71_done;
logic cond_wire71_in;
logic cond_wire71_out;
logic cond72_in;
logic cond72_write_en;
logic cond72_clk;
logic cond72_reset;
logic cond72_out;
logic cond72_done;
logic cond_wire72_in;
logic cond_wire72_out;
logic cond73_in;
logic cond73_write_en;
logic cond73_clk;
logic cond73_reset;
logic cond73_out;
logic cond73_done;
logic cond_wire73_in;
logic cond_wire73_out;
logic cond74_in;
logic cond74_write_en;
logic cond74_clk;
logic cond74_reset;
logic cond74_out;
logic cond74_done;
logic cond_wire74_in;
logic cond_wire74_out;
logic cond75_in;
logic cond75_write_en;
logic cond75_clk;
logic cond75_reset;
logic cond75_out;
logic cond75_done;
logic cond_wire75_in;
logic cond_wire75_out;
logic cond76_in;
logic cond76_write_en;
logic cond76_clk;
logic cond76_reset;
logic cond76_out;
logic cond76_done;
logic cond_wire76_in;
logic cond_wire76_out;
logic cond77_in;
logic cond77_write_en;
logic cond77_clk;
logic cond77_reset;
logic cond77_out;
logic cond77_done;
logic cond_wire77_in;
logic cond_wire77_out;
logic cond78_in;
logic cond78_write_en;
logic cond78_clk;
logic cond78_reset;
logic cond78_out;
logic cond78_done;
logic cond_wire78_in;
logic cond_wire78_out;
logic cond79_in;
logic cond79_write_en;
logic cond79_clk;
logic cond79_reset;
logic cond79_out;
logic cond79_done;
logic cond_wire79_in;
logic cond_wire79_out;
logic cond80_in;
logic cond80_write_en;
logic cond80_clk;
logic cond80_reset;
logic cond80_out;
logic cond80_done;
logic cond_wire80_in;
logic cond_wire80_out;
logic cond81_in;
logic cond81_write_en;
logic cond81_clk;
logic cond81_reset;
logic cond81_out;
logic cond81_done;
logic cond_wire81_in;
logic cond_wire81_out;
logic cond82_in;
logic cond82_write_en;
logic cond82_clk;
logic cond82_reset;
logic cond82_out;
logic cond82_done;
logic cond_wire82_in;
logic cond_wire82_out;
logic cond83_in;
logic cond83_write_en;
logic cond83_clk;
logic cond83_reset;
logic cond83_out;
logic cond83_done;
logic cond_wire83_in;
logic cond_wire83_out;
logic cond84_in;
logic cond84_write_en;
logic cond84_clk;
logic cond84_reset;
logic cond84_out;
logic cond84_done;
logic cond_wire84_in;
logic cond_wire84_out;
logic cond85_in;
logic cond85_write_en;
logic cond85_clk;
logic cond85_reset;
logic cond85_out;
logic cond85_done;
logic cond_wire85_in;
logic cond_wire85_out;
logic cond86_in;
logic cond86_write_en;
logic cond86_clk;
logic cond86_reset;
logic cond86_out;
logic cond86_done;
logic cond_wire86_in;
logic cond_wire86_out;
logic cond87_in;
logic cond87_write_en;
logic cond87_clk;
logic cond87_reset;
logic cond87_out;
logic cond87_done;
logic cond_wire87_in;
logic cond_wire87_out;
logic cond88_in;
logic cond88_write_en;
logic cond88_clk;
logic cond88_reset;
logic cond88_out;
logic cond88_done;
logic cond_wire88_in;
logic cond_wire88_out;
logic cond89_in;
logic cond89_write_en;
logic cond89_clk;
logic cond89_reset;
logic cond89_out;
logic cond89_done;
logic cond_wire89_in;
logic cond_wire89_out;
logic cond90_in;
logic cond90_write_en;
logic cond90_clk;
logic cond90_reset;
logic cond90_out;
logic cond90_done;
logic cond_wire90_in;
logic cond_wire90_out;
logic cond91_in;
logic cond91_write_en;
logic cond91_clk;
logic cond91_reset;
logic cond91_out;
logic cond91_done;
logic cond_wire91_in;
logic cond_wire91_out;
logic cond92_in;
logic cond92_write_en;
logic cond92_clk;
logic cond92_reset;
logic cond92_out;
logic cond92_done;
logic cond_wire92_in;
logic cond_wire92_out;
logic cond93_in;
logic cond93_write_en;
logic cond93_clk;
logic cond93_reset;
logic cond93_out;
logic cond93_done;
logic cond_wire93_in;
logic cond_wire93_out;
logic cond94_in;
logic cond94_write_en;
logic cond94_clk;
logic cond94_reset;
logic cond94_out;
logic cond94_done;
logic cond_wire94_in;
logic cond_wire94_out;
logic cond95_in;
logic cond95_write_en;
logic cond95_clk;
logic cond95_reset;
logic cond95_out;
logic cond95_done;
logic cond_wire95_in;
logic cond_wire95_out;
logic cond96_in;
logic cond96_write_en;
logic cond96_clk;
logic cond96_reset;
logic cond96_out;
logic cond96_done;
logic cond_wire96_in;
logic cond_wire96_out;
logic cond97_in;
logic cond97_write_en;
logic cond97_clk;
logic cond97_reset;
logic cond97_out;
logic cond97_done;
logic cond_wire97_in;
logic cond_wire97_out;
logic cond98_in;
logic cond98_write_en;
logic cond98_clk;
logic cond98_reset;
logic cond98_out;
logic cond98_done;
logic cond_wire98_in;
logic cond_wire98_out;
logic cond99_in;
logic cond99_write_en;
logic cond99_clk;
logic cond99_reset;
logic cond99_out;
logic cond99_done;
logic cond_wire99_in;
logic cond_wire99_out;
logic cond100_in;
logic cond100_write_en;
logic cond100_clk;
logic cond100_reset;
logic cond100_out;
logic cond100_done;
logic cond_wire100_in;
logic cond_wire100_out;
logic cond101_in;
logic cond101_write_en;
logic cond101_clk;
logic cond101_reset;
logic cond101_out;
logic cond101_done;
logic cond_wire101_in;
logic cond_wire101_out;
logic cond102_in;
logic cond102_write_en;
logic cond102_clk;
logic cond102_reset;
logic cond102_out;
logic cond102_done;
logic cond_wire102_in;
logic cond_wire102_out;
logic cond103_in;
logic cond103_write_en;
logic cond103_clk;
logic cond103_reset;
logic cond103_out;
logic cond103_done;
logic cond_wire103_in;
logic cond_wire103_out;
logic cond104_in;
logic cond104_write_en;
logic cond104_clk;
logic cond104_reset;
logic cond104_out;
logic cond104_done;
logic cond_wire104_in;
logic cond_wire104_out;
logic cond105_in;
logic cond105_write_en;
logic cond105_clk;
logic cond105_reset;
logic cond105_out;
logic cond105_done;
logic cond_wire105_in;
logic cond_wire105_out;
logic cond106_in;
logic cond106_write_en;
logic cond106_clk;
logic cond106_reset;
logic cond106_out;
logic cond106_done;
logic cond_wire106_in;
logic cond_wire106_out;
logic cond107_in;
logic cond107_write_en;
logic cond107_clk;
logic cond107_reset;
logic cond107_out;
logic cond107_done;
logic cond_wire107_in;
logic cond_wire107_out;
logic cond108_in;
logic cond108_write_en;
logic cond108_clk;
logic cond108_reset;
logic cond108_out;
logic cond108_done;
logic cond_wire108_in;
logic cond_wire108_out;
logic cond109_in;
logic cond109_write_en;
logic cond109_clk;
logic cond109_reset;
logic cond109_out;
logic cond109_done;
logic cond_wire109_in;
logic cond_wire109_out;
logic cond110_in;
logic cond110_write_en;
logic cond110_clk;
logic cond110_reset;
logic cond110_out;
logic cond110_done;
logic cond_wire110_in;
logic cond_wire110_out;
logic cond111_in;
logic cond111_write_en;
logic cond111_clk;
logic cond111_reset;
logic cond111_out;
logic cond111_done;
logic cond_wire111_in;
logic cond_wire111_out;
logic cond112_in;
logic cond112_write_en;
logic cond112_clk;
logic cond112_reset;
logic cond112_out;
logic cond112_done;
logic cond_wire112_in;
logic cond_wire112_out;
logic cond113_in;
logic cond113_write_en;
logic cond113_clk;
logic cond113_reset;
logic cond113_out;
logic cond113_done;
logic cond_wire113_in;
logic cond_wire113_out;
logic cond114_in;
logic cond114_write_en;
logic cond114_clk;
logic cond114_reset;
logic cond114_out;
logic cond114_done;
logic cond_wire114_in;
logic cond_wire114_out;
logic cond115_in;
logic cond115_write_en;
logic cond115_clk;
logic cond115_reset;
logic cond115_out;
logic cond115_done;
logic cond_wire115_in;
logic cond_wire115_out;
logic cond116_in;
logic cond116_write_en;
logic cond116_clk;
logic cond116_reset;
logic cond116_out;
logic cond116_done;
logic cond_wire116_in;
logic cond_wire116_out;
logic cond117_in;
logic cond117_write_en;
logic cond117_clk;
logic cond117_reset;
logic cond117_out;
logic cond117_done;
logic cond_wire117_in;
logic cond_wire117_out;
logic cond118_in;
logic cond118_write_en;
logic cond118_clk;
logic cond118_reset;
logic cond118_out;
logic cond118_done;
logic cond_wire118_in;
logic cond_wire118_out;
logic cond119_in;
logic cond119_write_en;
logic cond119_clk;
logic cond119_reset;
logic cond119_out;
logic cond119_done;
logic cond_wire119_in;
logic cond_wire119_out;
logic cond120_in;
logic cond120_write_en;
logic cond120_clk;
logic cond120_reset;
logic cond120_out;
logic cond120_done;
logic cond_wire120_in;
logic cond_wire120_out;
logic cond121_in;
logic cond121_write_en;
logic cond121_clk;
logic cond121_reset;
logic cond121_out;
logic cond121_done;
logic cond_wire121_in;
logic cond_wire121_out;
logic cond122_in;
logic cond122_write_en;
logic cond122_clk;
logic cond122_reset;
logic cond122_out;
logic cond122_done;
logic cond_wire122_in;
logic cond_wire122_out;
logic cond123_in;
logic cond123_write_en;
logic cond123_clk;
logic cond123_reset;
logic cond123_out;
logic cond123_done;
logic cond_wire123_in;
logic cond_wire123_out;
logic cond124_in;
logic cond124_write_en;
logic cond124_clk;
logic cond124_reset;
logic cond124_out;
logic cond124_done;
logic cond_wire124_in;
logic cond_wire124_out;
logic cond125_in;
logic cond125_write_en;
logic cond125_clk;
logic cond125_reset;
logic cond125_out;
logic cond125_done;
logic cond_wire125_in;
logic cond_wire125_out;
logic cond126_in;
logic cond126_write_en;
logic cond126_clk;
logic cond126_reset;
logic cond126_out;
logic cond126_done;
logic cond_wire126_in;
logic cond_wire126_out;
logic cond127_in;
logic cond127_write_en;
logic cond127_clk;
logic cond127_reset;
logic cond127_out;
logic cond127_done;
logic cond_wire127_in;
logic cond_wire127_out;
logic cond128_in;
logic cond128_write_en;
logic cond128_clk;
logic cond128_reset;
logic cond128_out;
logic cond128_done;
logic cond_wire128_in;
logic cond_wire128_out;
logic cond129_in;
logic cond129_write_en;
logic cond129_clk;
logic cond129_reset;
logic cond129_out;
logic cond129_done;
logic cond_wire129_in;
logic cond_wire129_out;
logic cond130_in;
logic cond130_write_en;
logic cond130_clk;
logic cond130_reset;
logic cond130_out;
logic cond130_done;
logic cond_wire130_in;
logic cond_wire130_out;
logic cond131_in;
logic cond131_write_en;
logic cond131_clk;
logic cond131_reset;
logic cond131_out;
logic cond131_done;
logic cond_wire131_in;
logic cond_wire131_out;
logic cond132_in;
logic cond132_write_en;
logic cond132_clk;
logic cond132_reset;
logic cond132_out;
logic cond132_done;
logic cond_wire132_in;
logic cond_wire132_out;
logic cond133_in;
logic cond133_write_en;
logic cond133_clk;
logic cond133_reset;
logic cond133_out;
logic cond133_done;
logic cond_wire133_in;
logic cond_wire133_out;
logic cond134_in;
logic cond134_write_en;
logic cond134_clk;
logic cond134_reset;
logic cond134_out;
logic cond134_done;
logic cond_wire134_in;
logic cond_wire134_out;
logic cond135_in;
logic cond135_write_en;
logic cond135_clk;
logic cond135_reset;
logic cond135_out;
logic cond135_done;
logic cond_wire135_in;
logic cond_wire135_out;
logic cond136_in;
logic cond136_write_en;
logic cond136_clk;
logic cond136_reset;
logic cond136_out;
logic cond136_done;
logic cond_wire136_in;
logic cond_wire136_out;
logic cond137_in;
logic cond137_write_en;
logic cond137_clk;
logic cond137_reset;
logic cond137_out;
logic cond137_done;
logic cond_wire137_in;
logic cond_wire137_out;
logic cond138_in;
logic cond138_write_en;
logic cond138_clk;
logic cond138_reset;
logic cond138_out;
logic cond138_done;
logic cond_wire138_in;
logic cond_wire138_out;
logic cond139_in;
logic cond139_write_en;
logic cond139_clk;
logic cond139_reset;
logic cond139_out;
logic cond139_done;
logic cond_wire139_in;
logic cond_wire139_out;
logic cond140_in;
logic cond140_write_en;
logic cond140_clk;
logic cond140_reset;
logic cond140_out;
logic cond140_done;
logic cond_wire140_in;
logic cond_wire140_out;
logic cond141_in;
logic cond141_write_en;
logic cond141_clk;
logic cond141_reset;
logic cond141_out;
logic cond141_done;
logic cond_wire141_in;
logic cond_wire141_out;
logic cond142_in;
logic cond142_write_en;
logic cond142_clk;
logic cond142_reset;
logic cond142_out;
logic cond142_done;
logic cond_wire142_in;
logic cond_wire142_out;
logic cond143_in;
logic cond143_write_en;
logic cond143_clk;
logic cond143_reset;
logic cond143_out;
logic cond143_done;
logic cond_wire143_in;
logic cond_wire143_out;
logic cond144_in;
logic cond144_write_en;
logic cond144_clk;
logic cond144_reset;
logic cond144_out;
logic cond144_done;
logic cond_wire144_in;
logic cond_wire144_out;
logic cond145_in;
logic cond145_write_en;
logic cond145_clk;
logic cond145_reset;
logic cond145_out;
logic cond145_done;
logic cond_wire145_in;
logic cond_wire145_out;
logic cond146_in;
logic cond146_write_en;
logic cond146_clk;
logic cond146_reset;
logic cond146_out;
logic cond146_done;
logic cond_wire146_in;
logic cond_wire146_out;
logic cond147_in;
logic cond147_write_en;
logic cond147_clk;
logic cond147_reset;
logic cond147_out;
logic cond147_done;
logic cond_wire147_in;
logic cond_wire147_out;
logic cond148_in;
logic cond148_write_en;
logic cond148_clk;
logic cond148_reset;
logic cond148_out;
logic cond148_done;
logic cond_wire148_in;
logic cond_wire148_out;
logic cond149_in;
logic cond149_write_en;
logic cond149_clk;
logic cond149_reset;
logic cond149_out;
logic cond149_done;
logic cond_wire149_in;
logic cond_wire149_out;
logic cond150_in;
logic cond150_write_en;
logic cond150_clk;
logic cond150_reset;
logic cond150_out;
logic cond150_done;
logic cond_wire150_in;
logic cond_wire150_out;
logic cond151_in;
logic cond151_write_en;
logic cond151_clk;
logic cond151_reset;
logic cond151_out;
logic cond151_done;
logic cond_wire151_in;
logic cond_wire151_out;
logic cond152_in;
logic cond152_write_en;
logic cond152_clk;
logic cond152_reset;
logic cond152_out;
logic cond152_done;
logic cond_wire152_in;
logic cond_wire152_out;
logic cond153_in;
logic cond153_write_en;
logic cond153_clk;
logic cond153_reset;
logic cond153_out;
logic cond153_done;
logic cond_wire153_in;
logic cond_wire153_out;
logic cond154_in;
logic cond154_write_en;
logic cond154_clk;
logic cond154_reset;
logic cond154_out;
logic cond154_done;
logic cond_wire154_in;
logic cond_wire154_out;
logic cond155_in;
logic cond155_write_en;
logic cond155_clk;
logic cond155_reset;
logic cond155_out;
logic cond155_done;
logic cond_wire155_in;
logic cond_wire155_out;
logic cond156_in;
logic cond156_write_en;
logic cond156_clk;
logic cond156_reset;
logic cond156_out;
logic cond156_done;
logic cond_wire156_in;
logic cond_wire156_out;
logic cond157_in;
logic cond157_write_en;
logic cond157_clk;
logic cond157_reset;
logic cond157_out;
logic cond157_done;
logic cond_wire157_in;
logic cond_wire157_out;
logic cond158_in;
logic cond158_write_en;
logic cond158_clk;
logic cond158_reset;
logic cond158_out;
logic cond158_done;
logic cond_wire158_in;
logic cond_wire158_out;
logic cond159_in;
logic cond159_write_en;
logic cond159_clk;
logic cond159_reset;
logic cond159_out;
logic cond159_done;
logic cond_wire159_in;
logic cond_wire159_out;
logic cond160_in;
logic cond160_write_en;
logic cond160_clk;
logic cond160_reset;
logic cond160_out;
logic cond160_done;
logic cond_wire160_in;
logic cond_wire160_out;
logic cond161_in;
logic cond161_write_en;
logic cond161_clk;
logic cond161_reset;
logic cond161_out;
logic cond161_done;
logic cond_wire161_in;
logic cond_wire161_out;
logic cond162_in;
logic cond162_write_en;
logic cond162_clk;
logic cond162_reset;
logic cond162_out;
logic cond162_done;
logic cond_wire162_in;
logic cond_wire162_out;
logic cond163_in;
logic cond163_write_en;
logic cond163_clk;
logic cond163_reset;
logic cond163_out;
logic cond163_done;
logic cond_wire163_in;
logic cond_wire163_out;
logic cond164_in;
logic cond164_write_en;
logic cond164_clk;
logic cond164_reset;
logic cond164_out;
logic cond164_done;
logic cond_wire164_in;
logic cond_wire164_out;
logic cond165_in;
logic cond165_write_en;
logic cond165_clk;
logic cond165_reset;
logic cond165_out;
logic cond165_done;
logic cond_wire165_in;
logic cond_wire165_out;
logic cond166_in;
logic cond166_write_en;
logic cond166_clk;
logic cond166_reset;
logic cond166_out;
logic cond166_done;
logic cond_wire166_in;
logic cond_wire166_out;
logic cond167_in;
logic cond167_write_en;
logic cond167_clk;
logic cond167_reset;
logic cond167_out;
logic cond167_done;
logic cond_wire167_in;
logic cond_wire167_out;
logic cond168_in;
logic cond168_write_en;
logic cond168_clk;
logic cond168_reset;
logic cond168_out;
logic cond168_done;
logic cond_wire168_in;
logic cond_wire168_out;
logic cond169_in;
logic cond169_write_en;
logic cond169_clk;
logic cond169_reset;
logic cond169_out;
logic cond169_done;
logic cond_wire169_in;
logic cond_wire169_out;
logic cond170_in;
logic cond170_write_en;
logic cond170_clk;
logic cond170_reset;
logic cond170_out;
logic cond170_done;
logic cond_wire170_in;
logic cond_wire170_out;
logic cond171_in;
logic cond171_write_en;
logic cond171_clk;
logic cond171_reset;
logic cond171_out;
logic cond171_done;
logic cond_wire171_in;
logic cond_wire171_out;
logic cond172_in;
logic cond172_write_en;
logic cond172_clk;
logic cond172_reset;
logic cond172_out;
logic cond172_done;
logic cond_wire172_in;
logic cond_wire172_out;
logic cond173_in;
logic cond173_write_en;
logic cond173_clk;
logic cond173_reset;
logic cond173_out;
logic cond173_done;
logic cond_wire173_in;
logic cond_wire173_out;
logic cond174_in;
logic cond174_write_en;
logic cond174_clk;
logic cond174_reset;
logic cond174_out;
logic cond174_done;
logic cond_wire174_in;
logic cond_wire174_out;
logic cond175_in;
logic cond175_write_en;
logic cond175_clk;
logic cond175_reset;
logic cond175_out;
logic cond175_done;
logic cond_wire175_in;
logic cond_wire175_out;
logic cond176_in;
logic cond176_write_en;
logic cond176_clk;
logic cond176_reset;
logic cond176_out;
logic cond176_done;
logic cond_wire176_in;
logic cond_wire176_out;
logic cond177_in;
logic cond177_write_en;
logic cond177_clk;
logic cond177_reset;
logic cond177_out;
logic cond177_done;
logic cond_wire177_in;
logic cond_wire177_out;
logic cond178_in;
logic cond178_write_en;
logic cond178_clk;
logic cond178_reset;
logic cond178_out;
logic cond178_done;
logic cond_wire178_in;
logic cond_wire178_out;
logic cond179_in;
logic cond179_write_en;
logic cond179_clk;
logic cond179_reset;
logic cond179_out;
logic cond179_done;
logic cond_wire179_in;
logic cond_wire179_out;
logic cond180_in;
logic cond180_write_en;
logic cond180_clk;
logic cond180_reset;
logic cond180_out;
logic cond180_done;
logic cond_wire180_in;
logic cond_wire180_out;
logic cond181_in;
logic cond181_write_en;
logic cond181_clk;
logic cond181_reset;
logic cond181_out;
logic cond181_done;
logic cond_wire181_in;
logic cond_wire181_out;
logic cond182_in;
logic cond182_write_en;
logic cond182_clk;
logic cond182_reset;
logic cond182_out;
logic cond182_done;
logic cond_wire182_in;
logic cond_wire182_out;
logic cond183_in;
logic cond183_write_en;
logic cond183_clk;
logic cond183_reset;
logic cond183_out;
logic cond183_done;
logic cond_wire183_in;
logic cond_wire183_out;
logic cond184_in;
logic cond184_write_en;
logic cond184_clk;
logic cond184_reset;
logic cond184_out;
logic cond184_done;
logic cond_wire184_in;
logic cond_wire184_out;
logic cond185_in;
logic cond185_write_en;
logic cond185_clk;
logic cond185_reset;
logic cond185_out;
logic cond185_done;
logic cond_wire185_in;
logic cond_wire185_out;
logic cond186_in;
logic cond186_write_en;
logic cond186_clk;
logic cond186_reset;
logic cond186_out;
logic cond186_done;
logic cond_wire186_in;
logic cond_wire186_out;
logic cond187_in;
logic cond187_write_en;
logic cond187_clk;
logic cond187_reset;
logic cond187_out;
logic cond187_done;
logic cond_wire187_in;
logic cond_wire187_out;
logic cond188_in;
logic cond188_write_en;
logic cond188_clk;
logic cond188_reset;
logic cond188_out;
logic cond188_done;
logic cond_wire188_in;
logic cond_wire188_out;
logic cond189_in;
logic cond189_write_en;
logic cond189_clk;
logic cond189_reset;
logic cond189_out;
logic cond189_done;
logic cond_wire189_in;
logic cond_wire189_out;
logic cond190_in;
logic cond190_write_en;
logic cond190_clk;
logic cond190_reset;
logic cond190_out;
logic cond190_done;
logic cond_wire190_in;
logic cond_wire190_out;
logic cond191_in;
logic cond191_write_en;
logic cond191_clk;
logic cond191_reset;
logic cond191_out;
logic cond191_done;
logic cond_wire191_in;
logic cond_wire191_out;
logic cond192_in;
logic cond192_write_en;
logic cond192_clk;
logic cond192_reset;
logic cond192_out;
logic cond192_done;
logic cond_wire192_in;
logic cond_wire192_out;
logic cond193_in;
logic cond193_write_en;
logic cond193_clk;
logic cond193_reset;
logic cond193_out;
logic cond193_done;
logic cond_wire193_in;
logic cond_wire193_out;
logic cond194_in;
logic cond194_write_en;
logic cond194_clk;
logic cond194_reset;
logic cond194_out;
logic cond194_done;
logic cond_wire194_in;
logic cond_wire194_out;
logic cond195_in;
logic cond195_write_en;
logic cond195_clk;
logic cond195_reset;
logic cond195_out;
logic cond195_done;
logic cond_wire195_in;
logic cond_wire195_out;
logic cond196_in;
logic cond196_write_en;
logic cond196_clk;
logic cond196_reset;
logic cond196_out;
logic cond196_done;
logic cond_wire196_in;
logic cond_wire196_out;
logic cond197_in;
logic cond197_write_en;
logic cond197_clk;
logic cond197_reset;
logic cond197_out;
logic cond197_done;
logic cond_wire197_in;
logic cond_wire197_out;
logic cond198_in;
logic cond198_write_en;
logic cond198_clk;
logic cond198_reset;
logic cond198_out;
logic cond198_done;
logic cond_wire198_in;
logic cond_wire198_out;
logic cond199_in;
logic cond199_write_en;
logic cond199_clk;
logic cond199_reset;
logic cond199_out;
logic cond199_done;
logic cond_wire199_in;
logic cond_wire199_out;
logic cond200_in;
logic cond200_write_en;
logic cond200_clk;
logic cond200_reset;
logic cond200_out;
logic cond200_done;
logic cond_wire200_in;
logic cond_wire200_out;
logic cond201_in;
logic cond201_write_en;
logic cond201_clk;
logic cond201_reset;
logic cond201_out;
logic cond201_done;
logic cond_wire201_in;
logic cond_wire201_out;
logic cond202_in;
logic cond202_write_en;
logic cond202_clk;
logic cond202_reset;
logic cond202_out;
logic cond202_done;
logic cond_wire202_in;
logic cond_wire202_out;
logic cond203_in;
logic cond203_write_en;
logic cond203_clk;
logic cond203_reset;
logic cond203_out;
logic cond203_done;
logic cond_wire203_in;
logic cond_wire203_out;
logic cond204_in;
logic cond204_write_en;
logic cond204_clk;
logic cond204_reset;
logic cond204_out;
logic cond204_done;
logic cond_wire204_in;
logic cond_wire204_out;
logic cond205_in;
logic cond205_write_en;
logic cond205_clk;
logic cond205_reset;
logic cond205_out;
logic cond205_done;
logic cond_wire205_in;
logic cond_wire205_out;
logic cond206_in;
logic cond206_write_en;
logic cond206_clk;
logic cond206_reset;
logic cond206_out;
logic cond206_done;
logic cond_wire206_in;
logic cond_wire206_out;
logic cond207_in;
logic cond207_write_en;
logic cond207_clk;
logic cond207_reset;
logic cond207_out;
logic cond207_done;
logic cond_wire207_in;
logic cond_wire207_out;
logic cond208_in;
logic cond208_write_en;
logic cond208_clk;
logic cond208_reset;
logic cond208_out;
logic cond208_done;
logic cond_wire208_in;
logic cond_wire208_out;
logic cond209_in;
logic cond209_write_en;
logic cond209_clk;
logic cond209_reset;
logic cond209_out;
logic cond209_done;
logic cond_wire209_in;
logic cond_wire209_out;
logic cond210_in;
logic cond210_write_en;
logic cond210_clk;
logic cond210_reset;
logic cond210_out;
logic cond210_done;
logic cond_wire210_in;
logic cond_wire210_out;
logic cond211_in;
logic cond211_write_en;
logic cond211_clk;
logic cond211_reset;
logic cond211_out;
logic cond211_done;
logic cond_wire211_in;
logic cond_wire211_out;
logic cond212_in;
logic cond212_write_en;
logic cond212_clk;
logic cond212_reset;
logic cond212_out;
logic cond212_done;
logic cond_wire212_in;
logic cond_wire212_out;
logic cond213_in;
logic cond213_write_en;
logic cond213_clk;
logic cond213_reset;
logic cond213_out;
logic cond213_done;
logic cond_wire213_in;
logic cond_wire213_out;
logic cond214_in;
logic cond214_write_en;
logic cond214_clk;
logic cond214_reset;
logic cond214_out;
logic cond214_done;
logic cond_wire214_in;
logic cond_wire214_out;
logic cond215_in;
logic cond215_write_en;
logic cond215_clk;
logic cond215_reset;
logic cond215_out;
logic cond215_done;
logic cond_wire215_in;
logic cond_wire215_out;
logic cond216_in;
logic cond216_write_en;
logic cond216_clk;
logic cond216_reset;
logic cond216_out;
logic cond216_done;
logic cond_wire216_in;
logic cond_wire216_out;
logic cond217_in;
logic cond217_write_en;
logic cond217_clk;
logic cond217_reset;
logic cond217_out;
logic cond217_done;
logic cond_wire217_in;
logic cond_wire217_out;
logic cond218_in;
logic cond218_write_en;
logic cond218_clk;
logic cond218_reset;
logic cond218_out;
logic cond218_done;
logic cond_wire218_in;
logic cond_wire218_out;
logic cond219_in;
logic cond219_write_en;
logic cond219_clk;
logic cond219_reset;
logic cond219_out;
logic cond219_done;
logic cond_wire219_in;
logic cond_wire219_out;
logic cond220_in;
logic cond220_write_en;
logic cond220_clk;
logic cond220_reset;
logic cond220_out;
logic cond220_done;
logic cond_wire220_in;
logic cond_wire220_out;
logic cond221_in;
logic cond221_write_en;
logic cond221_clk;
logic cond221_reset;
logic cond221_out;
logic cond221_done;
logic cond_wire221_in;
logic cond_wire221_out;
logic cond222_in;
logic cond222_write_en;
logic cond222_clk;
logic cond222_reset;
logic cond222_out;
logic cond222_done;
logic cond_wire222_in;
logic cond_wire222_out;
logic cond223_in;
logic cond223_write_en;
logic cond223_clk;
logic cond223_reset;
logic cond223_out;
logic cond223_done;
logic cond_wire223_in;
logic cond_wire223_out;
logic cond224_in;
logic cond224_write_en;
logic cond224_clk;
logic cond224_reset;
logic cond224_out;
logic cond224_done;
logic cond_wire224_in;
logic cond_wire224_out;
logic cond225_in;
logic cond225_write_en;
logic cond225_clk;
logic cond225_reset;
logic cond225_out;
logic cond225_done;
logic cond_wire225_in;
logic cond_wire225_out;
logic cond226_in;
logic cond226_write_en;
logic cond226_clk;
logic cond226_reset;
logic cond226_out;
logic cond226_done;
logic cond_wire226_in;
logic cond_wire226_out;
logic cond227_in;
logic cond227_write_en;
logic cond227_clk;
logic cond227_reset;
logic cond227_out;
logic cond227_done;
logic cond_wire227_in;
logic cond_wire227_out;
logic cond228_in;
logic cond228_write_en;
logic cond228_clk;
logic cond228_reset;
logic cond228_out;
logic cond228_done;
logic cond_wire228_in;
logic cond_wire228_out;
logic cond229_in;
logic cond229_write_en;
logic cond229_clk;
logic cond229_reset;
logic cond229_out;
logic cond229_done;
logic cond_wire229_in;
logic cond_wire229_out;
logic cond230_in;
logic cond230_write_en;
logic cond230_clk;
logic cond230_reset;
logic cond230_out;
logic cond230_done;
logic cond_wire230_in;
logic cond_wire230_out;
logic cond231_in;
logic cond231_write_en;
logic cond231_clk;
logic cond231_reset;
logic cond231_out;
logic cond231_done;
logic cond_wire231_in;
logic cond_wire231_out;
logic cond232_in;
logic cond232_write_en;
logic cond232_clk;
logic cond232_reset;
logic cond232_out;
logic cond232_done;
logic cond_wire232_in;
logic cond_wire232_out;
logic cond233_in;
logic cond233_write_en;
logic cond233_clk;
logic cond233_reset;
logic cond233_out;
logic cond233_done;
logic cond_wire233_in;
logic cond_wire233_out;
logic cond234_in;
logic cond234_write_en;
logic cond234_clk;
logic cond234_reset;
logic cond234_out;
logic cond234_done;
logic cond_wire234_in;
logic cond_wire234_out;
logic cond235_in;
logic cond235_write_en;
logic cond235_clk;
logic cond235_reset;
logic cond235_out;
logic cond235_done;
logic cond_wire235_in;
logic cond_wire235_out;
logic cond236_in;
logic cond236_write_en;
logic cond236_clk;
logic cond236_reset;
logic cond236_out;
logic cond236_done;
logic cond_wire236_in;
logic cond_wire236_out;
logic cond237_in;
logic cond237_write_en;
logic cond237_clk;
logic cond237_reset;
logic cond237_out;
logic cond237_done;
logic cond_wire237_in;
logic cond_wire237_out;
logic cond238_in;
logic cond238_write_en;
logic cond238_clk;
logic cond238_reset;
logic cond238_out;
logic cond238_done;
logic cond_wire238_in;
logic cond_wire238_out;
logic cond239_in;
logic cond239_write_en;
logic cond239_clk;
logic cond239_reset;
logic cond239_out;
logic cond239_done;
logic cond_wire239_in;
logic cond_wire239_out;
logic cond240_in;
logic cond240_write_en;
logic cond240_clk;
logic cond240_reset;
logic cond240_out;
logic cond240_done;
logic cond_wire240_in;
logic cond_wire240_out;
logic cond241_in;
logic cond241_write_en;
logic cond241_clk;
logic cond241_reset;
logic cond241_out;
logic cond241_done;
logic cond_wire241_in;
logic cond_wire241_out;
logic cond242_in;
logic cond242_write_en;
logic cond242_clk;
logic cond242_reset;
logic cond242_out;
logic cond242_done;
logic cond_wire242_in;
logic cond_wire242_out;
logic cond243_in;
logic cond243_write_en;
logic cond243_clk;
logic cond243_reset;
logic cond243_out;
logic cond243_done;
logic cond_wire243_in;
logic cond_wire243_out;
logic cond244_in;
logic cond244_write_en;
logic cond244_clk;
logic cond244_reset;
logic cond244_out;
logic cond244_done;
logic cond_wire244_in;
logic cond_wire244_out;
logic cond245_in;
logic cond245_write_en;
logic cond245_clk;
logic cond245_reset;
logic cond245_out;
logic cond245_done;
logic cond_wire245_in;
logic cond_wire245_out;
logic cond246_in;
logic cond246_write_en;
logic cond246_clk;
logic cond246_reset;
logic cond246_out;
logic cond246_done;
logic cond_wire246_in;
logic cond_wire246_out;
logic cond247_in;
logic cond247_write_en;
logic cond247_clk;
logic cond247_reset;
logic cond247_out;
logic cond247_done;
logic cond_wire247_in;
logic cond_wire247_out;
logic cond248_in;
logic cond248_write_en;
logic cond248_clk;
logic cond248_reset;
logic cond248_out;
logic cond248_done;
logic cond_wire248_in;
logic cond_wire248_out;
logic cond249_in;
logic cond249_write_en;
logic cond249_clk;
logic cond249_reset;
logic cond249_out;
logic cond249_done;
logic cond_wire249_in;
logic cond_wire249_out;
logic cond250_in;
logic cond250_write_en;
logic cond250_clk;
logic cond250_reset;
logic cond250_out;
logic cond250_done;
logic cond_wire250_in;
logic cond_wire250_out;
logic cond251_in;
logic cond251_write_en;
logic cond251_clk;
logic cond251_reset;
logic cond251_out;
logic cond251_done;
logic cond_wire251_in;
logic cond_wire251_out;
logic cond252_in;
logic cond252_write_en;
logic cond252_clk;
logic cond252_reset;
logic cond252_out;
logic cond252_done;
logic cond_wire252_in;
logic cond_wire252_out;
logic cond253_in;
logic cond253_write_en;
logic cond253_clk;
logic cond253_reset;
logic cond253_out;
logic cond253_done;
logic cond_wire253_in;
logic cond_wire253_out;
logic cond254_in;
logic cond254_write_en;
logic cond254_clk;
logic cond254_reset;
logic cond254_out;
logic cond254_done;
logic cond_wire254_in;
logic cond_wire254_out;
logic cond255_in;
logic cond255_write_en;
logic cond255_clk;
logic cond255_reset;
logic cond255_out;
logic cond255_done;
logic cond_wire255_in;
logic cond_wire255_out;
logic cond256_in;
logic cond256_write_en;
logic cond256_clk;
logic cond256_reset;
logic cond256_out;
logic cond256_done;
logic cond_wire256_in;
logic cond_wire256_out;
logic cond257_in;
logic cond257_write_en;
logic cond257_clk;
logic cond257_reset;
logic cond257_out;
logic cond257_done;
logic cond_wire257_in;
logic cond_wire257_out;
logic cond258_in;
logic cond258_write_en;
logic cond258_clk;
logic cond258_reset;
logic cond258_out;
logic cond258_done;
logic cond_wire258_in;
logic cond_wire258_out;
logic cond259_in;
logic cond259_write_en;
logic cond259_clk;
logic cond259_reset;
logic cond259_out;
logic cond259_done;
logic cond_wire259_in;
logic cond_wire259_out;
logic cond260_in;
logic cond260_write_en;
logic cond260_clk;
logic cond260_reset;
logic cond260_out;
logic cond260_done;
logic cond_wire260_in;
logic cond_wire260_out;
logic cond261_in;
logic cond261_write_en;
logic cond261_clk;
logic cond261_reset;
logic cond261_out;
logic cond261_done;
logic cond_wire261_in;
logic cond_wire261_out;
logic cond262_in;
logic cond262_write_en;
logic cond262_clk;
logic cond262_reset;
logic cond262_out;
logic cond262_done;
logic cond_wire262_in;
logic cond_wire262_out;
logic cond263_in;
logic cond263_write_en;
logic cond263_clk;
logic cond263_reset;
logic cond263_out;
logic cond263_done;
logic cond_wire263_in;
logic cond_wire263_out;
logic cond264_in;
logic cond264_write_en;
logic cond264_clk;
logic cond264_reset;
logic cond264_out;
logic cond264_done;
logic cond_wire264_in;
logic cond_wire264_out;
logic cond265_in;
logic cond265_write_en;
logic cond265_clk;
logic cond265_reset;
logic cond265_out;
logic cond265_done;
logic cond_wire265_in;
logic cond_wire265_out;
logic cond266_in;
logic cond266_write_en;
logic cond266_clk;
logic cond266_reset;
logic cond266_out;
logic cond266_done;
logic cond_wire266_in;
logic cond_wire266_out;
logic cond267_in;
logic cond267_write_en;
logic cond267_clk;
logic cond267_reset;
logic cond267_out;
logic cond267_done;
logic cond_wire267_in;
logic cond_wire267_out;
logic cond268_in;
logic cond268_write_en;
logic cond268_clk;
logic cond268_reset;
logic cond268_out;
logic cond268_done;
logic cond_wire268_in;
logic cond_wire268_out;
logic cond269_in;
logic cond269_write_en;
logic cond269_clk;
logic cond269_reset;
logic cond269_out;
logic cond269_done;
logic cond_wire269_in;
logic cond_wire269_out;
logic cond270_in;
logic cond270_write_en;
logic cond270_clk;
logic cond270_reset;
logic cond270_out;
logic cond270_done;
logic cond_wire270_in;
logic cond_wire270_out;
logic cond271_in;
logic cond271_write_en;
logic cond271_clk;
logic cond271_reset;
logic cond271_out;
logic cond271_done;
logic cond_wire271_in;
logic cond_wire271_out;
logic cond272_in;
logic cond272_write_en;
logic cond272_clk;
logic cond272_reset;
logic cond272_out;
logic cond272_done;
logic cond_wire272_in;
logic cond_wire272_out;
logic cond273_in;
logic cond273_write_en;
logic cond273_clk;
logic cond273_reset;
logic cond273_out;
logic cond273_done;
logic cond_wire273_in;
logic cond_wire273_out;
logic cond274_in;
logic cond274_write_en;
logic cond274_clk;
logic cond274_reset;
logic cond274_out;
logic cond274_done;
logic cond_wire274_in;
logic cond_wire274_out;
logic cond275_in;
logic cond275_write_en;
logic cond275_clk;
logic cond275_reset;
logic cond275_out;
logic cond275_done;
logic cond_wire275_in;
logic cond_wire275_out;
logic cond276_in;
logic cond276_write_en;
logic cond276_clk;
logic cond276_reset;
logic cond276_out;
logic cond276_done;
logic cond_wire276_in;
logic cond_wire276_out;
logic cond277_in;
logic cond277_write_en;
logic cond277_clk;
logic cond277_reset;
logic cond277_out;
logic cond277_done;
logic cond_wire277_in;
logic cond_wire277_out;
logic cond278_in;
logic cond278_write_en;
logic cond278_clk;
logic cond278_reset;
logic cond278_out;
logic cond278_done;
logic cond_wire278_in;
logic cond_wire278_out;
logic cond279_in;
logic cond279_write_en;
logic cond279_clk;
logic cond279_reset;
logic cond279_out;
logic cond279_done;
logic cond_wire279_in;
logic cond_wire279_out;
logic cond280_in;
logic cond280_write_en;
logic cond280_clk;
logic cond280_reset;
logic cond280_out;
logic cond280_done;
logic cond_wire280_in;
logic cond_wire280_out;
logic cond281_in;
logic cond281_write_en;
logic cond281_clk;
logic cond281_reset;
logic cond281_out;
logic cond281_done;
logic cond_wire281_in;
logic cond_wire281_out;
logic cond282_in;
logic cond282_write_en;
logic cond282_clk;
logic cond282_reset;
logic cond282_out;
logic cond282_done;
logic cond_wire282_in;
logic cond_wire282_out;
logic cond283_in;
logic cond283_write_en;
logic cond283_clk;
logic cond283_reset;
logic cond283_out;
logic cond283_done;
logic cond_wire283_in;
logic cond_wire283_out;
logic cond284_in;
logic cond284_write_en;
logic cond284_clk;
logic cond284_reset;
logic cond284_out;
logic cond284_done;
logic cond_wire284_in;
logic cond_wire284_out;
logic cond285_in;
logic cond285_write_en;
logic cond285_clk;
logic cond285_reset;
logic cond285_out;
logic cond285_done;
logic cond_wire285_in;
logic cond_wire285_out;
logic cond286_in;
logic cond286_write_en;
logic cond286_clk;
logic cond286_reset;
logic cond286_out;
logic cond286_done;
logic cond_wire286_in;
logic cond_wire286_out;
logic cond287_in;
logic cond287_write_en;
logic cond287_clk;
logic cond287_reset;
logic cond287_out;
logic cond287_done;
logic cond_wire287_in;
logic cond_wire287_out;
logic cond288_in;
logic cond288_write_en;
logic cond288_clk;
logic cond288_reset;
logic cond288_out;
logic cond288_done;
logic cond_wire288_in;
logic cond_wire288_out;
logic cond289_in;
logic cond289_write_en;
logic cond289_clk;
logic cond289_reset;
logic cond289_out;
logic cond289_done;
logic cond_wire289_in;
logic cond_wire289_out;
logic cond290_in;
logic cond290_write_en;
logic cond290_clk;
logic cond290_reset;
logic cond290_out;
logic cond290_done;
logic cond_wire290_in;
logic cond_wire290_out;
logic cond291_in;
logic cond291_write_en;
logic cond291_clk;
logic cond291_reset;
logic cond291_out;
logic cond291_done;
logic cond_wire291_in;
logic cond_wire291_out;
logic cond292_in;
logic cond292_write_en;
logic cond292_clk;
logic cond292_reset;
logic cond292_out;
logic cond292_done;
logic cond_wire292_in;
logic cond_wire292_out;
logic cond293_in;
logic cond293_write_en;
logic cond293_clk;
logic cond293_reset;
logic cond293_out;
logic cond293_done;
logic cond_wire293_in;
logic cond_wire293_out;
logic cond294_in;
logic cond294_write_en;
logic cond294_clk;
logic cond294_reset;
logic cond294_out;
logic cond294_done;
logic cond_wire294_in;
logic cond_wire294_out;
logic cond295_in;
logic cond295_write_en;
logic cond295_clk;
logic cond295_reset;
logic cond295_out;
logic cond295_done;
logic cond_wire295_in;
logic cond_wire295_out;
logic cond296_in;
logic cond296_write_en;
logic cond296_clk;
logic cond296_reset;
logic cond296_out;
logic cond296_done;
logic cond_wire296_in;
logic cond_wire296_out;
logic cond297_in;
logic cond297_write_en;
logic cond297_clk;
logic cond297_reset;
logic cond297_out;
logic cond297_done;
logic cond_wire297_in;
logic cond_wire297_out;
logic cond298_in;
logic cond298_write_en;
logic cond298_clk;
logic cond298_reset;
logic cond298_out;
logic cond298_done;
logic cond_wire298_in;
logic cond_wire298_out;
logic cond299_in;
logic cond299_write_en;
logic cond299_clk;
logic cond299_reset;
logic cond299_out;
logic cond299_done;
logic cond_wire299_in;
logic cond_wire299_out;
logic cond300_in;
logic cond300_write_en;
logic cond300_clk;
logic cond300_reset;
logic cond300_out;
logic cond300_done;
logic cond_wire300_in;
logic cond_wire300_out;
logic cond301_in;
logic cond301_write_en;
logic cond301_clk;
logic cond301_reset;
logic cond301_out;
logic cond301_done;
logic cond_wire301_in;
logic cond_wire301_out;
logic cond302_in;
logic cond302_write_en;
logic cond302_clk;
logic cond302_reset;
logic cond302_out;
logic cond302_done;
logic cond_wire302_in;
logic cond_wire302_out;
logic cond303_in;
logic cond303_write_en;
logic cond303_clk;
logic cond303_reset;
logic cond303_out;
logic cond303_done;
logic cond_wire303_in;
logic cond_wire303_out;
logic cond304_in;
logic cond304_write_en;
logic cond304_clk;
logic cond304_reset;
logic cond304_out;
logic cond304_done;
logic cond_wire304_in;
logic cond_wire304_out;
logic cond305_in;
logic cond305_write_en;
logic cond305_clk;
logic cond305_reset;
logic cond305_out;
logic cond305_done;
logic cond_wire305_in;
logic cond_wire305_out;
logic cond306_in;
logic cond306_write_en;
logic cond306_clk;
logic cond306_reset;
logic cond306_out;
logic cond306_done;
logic cond_wire306_in;
logic cond_wire306_out;
logic cond307_in;
logic cond307_write_en;
logic cond307_clk;
logic cond307_reset;
logic cond307_out;
logic cond307_done;
logic cond_wire307_in;
logic cond_wire307_out;
logic cond308_in;
logic cond308_write_en;
logic cond308_clk;
logic cond308_reset;
logic cond308_out;
logic cond308_done;
logic cond_wire308_in;
logic cond_wire308_out;
logic cond309_in;
logic cond309_write_en;
logic cond309_clk;
logic cond309_reset;
logic cond309_out;
logic cond309_done;
logic cond_wire309_in;
logic cond_wire309_out;
logic cond310_in;
logic cond310_write_en;
logic cond310_clk;
logic cond310_reset;
logic cond310_out;
logic cond310_done;
logic cond_wire310_in;
logic cond_wire310_out;
logic cond311_in;
logic cond311_write_en;
logic cond311_clk;
logic cond311_reset;
logic cond311_out;
logic cond311_done;
logic cond_wire311_in;
logic cond_wire311_out;
logic cond312_in;
logic cond312_write_en;
logic cond312_clk;
logic cond312_reset;
logic cond312_out;
logic cond312_done;
logic cond_wire312_in;
logic cond_wire312_out;
logic cond313_in;
logic cond313_write_en;
logic cond313_clk;
logic cond313_reset;
logic cond313_out;
logic cond313_done;
logic cond_wire313_in;
logic cond_wire313_out;
logic cond314_in;
logic cond314_write_en;
logic cond314_clk;
logic cond314_reset;
logic cond314_out;
logic cond314_done;
logic cond_wire314_in;
logic cond_wire314_out;
logic cond315_in;
logic cond315_write_en;
logic cond315_clk;
logic cond315_reset;
logic cond315_out;
logic cond315_done;
logic cond_wire315_in;
logic cond_wire315_out;
logic cond316_in;
logic cond316_write_en;
logic cond316_clk;
logic cond316_reset;
logic cond316_out;
logic cond316_done;
logic cond_wire316_in;
logic cond_wire316_out;
logic cond317_in;
logic cond317_write_en;
logic cond317_clk;
logic cond317_reset;
logic cond317_out;
logic cond317_done;
logic cond_wire317_in;
logic cond_wire317_out;
logic cond318_in;
logic cond318_write_en;
logic cond318_clk;
logic cond318_reset;
logic cond318_out;
logic cond318_done;
logic cond_wire318_in;
logic cond_wire318_out;
logic cond319_in;
logic cond319_write_en;
logic cond319_clk;
logic cond319_reset;
logic cond319_out;
logic cond319_done;
logic cond_wire319_in;
logic cond_wire319_out;
logic cond320_in;
logic cond320_write_en;
logic cond320_clk;
logic cond320_reset;
logic cond320_out;
logic cond320_done;
logic cond_wire320_in;
logic cond_wire320_out;
logic cond321_in;
logic cond321_write_en;
logic cond321_clk;
logic cond321_reset;
logic cond321_out;
logic cond321_done;
logic cond_wire321_in;
logic cond_wire321_out;
logic cond322_in;
logic cond322_write_en;
logic cond322_clk;
logic cond322_reset;
logic cond322_out;
logic cond322_done;
logic cond_wire322_in;
logic cond_wire322_out;
logic cond323_in;
logic cond323_write_en;
logic cond323_clk;
logic cond323_reset;
logic cond323_out;
logic cond323_done;
logic cond_wire323_in;
logic cond_wire323_out;
logic cond324_in;
logic cond324_write_en;
logic cond324_clk;
logic cond324_reset;
logic cond324_out;
logic cond324_done;
logic cond_wire324_in;
logic cond_wire324_out;
logic cond325_in;
logic cond325_write_en;
logic cond325_clk;
logic cond325_reset;
logic cond325_out;
logic cond325_done;
logic cond_wire325_in;
logic cond_wire325_out;
logic cond326_in;
logic cond326_write_en;
logic cond326_clk;
logic cond326_reset;
logic cond326_out;
logic cond326_done;
logic cond_wire326_in;
logic cond_wire326_out;
logic cond327_in;
logic cond327_write_en;
logic cond327_clk;
logic cond327_reset;
logic cond327_out;
logic cond327_done;
logic cond_wire327_in;
logic cond_wire327_out;
logic cond328_in;
logic cond328_write_en;
logic cond328_clk;
logic cond328_reset;
logic cond328_out;
logic cond328_done;
logic cond_wire328_in;
logic cond_wire328_out;
logic cond329_in;
logic cond329_write_en;
logic cond329_clk;
logic cond329_reset;
logic cond329_out;
logic cond329_done;
logic cond_wire329_in;
logic cond_wire329_out;
logic cond330_in;
logic cond330_write_en;
logic cond330_clk;
logic cond330_reset;
logic cond330_out;
logic cond330_done;
logic cond_wire330_in;
logic cond_wire330_out;
logic cond331_in;
logic cond331_write_en;
logic cond331_clk;
logic cond331_reset;
logic cond331_out;
logic cond331_done;
logic cond_wire331_in;
logic cond_wire331_out;
logic cond332_in;
logic cond332_write_en;
logic cond332_clk;
logic cond332_reset;
logic cond332_out;
logic cond332_done;
logic cond_wire332_in;
logic cond_wire332_out;
logic cond333_in;
logic cond333_write_en;
logic cond333_clk;
logic cond333_reset;
logic cond333_out;
logic cond333_done;
logic cond_wire333_in;
logic cond_wire333_out;
logic cond334_in;
logic cond334_write_en;
logic cond334_clk;
logic cond334_reset;
logic cond334_out;
logic cond334_done;
logic cond_wire334_in;
logic cond_wire334_out;
logic cond335_in;
logic cond335_write_en;
logic cond335_clk;
logic cond335_reset;
logic cond335_out;
logic cond335_done;
logic cond_wire335_in;
logic cond_wire335_out;
logic cond336_in;
logic cond336_write_en;
logic cond336_clk;
logic cond336_reset;
logic cond336_out;
logic cond336_done;
logic cond_wire336_in;
logic cond_wire336_out;
logic cond337_in;
logic cond337_write_en;
logic cond337_clk;
logic cond337_reset;
logic cond337_out;
logic cond337_done;
logic cond_wire337_in;
logic cond_wire337_out;
logic cond338_in;
logic cond338_write_en;
logic cond338_clk;
logic cond338_reset;
logic cond338_out;
logic cond338_done;
logic cond_wire338_in;
logic cond_wire338_out;
logic cond339_in;
logic cond339_write_en;
logic cond339_clk;
logic cond339_reset;
logic cond339_out;
logic cond339_done;
logic cond_wire339_in;
logic cond_wire339_out;
logic cond340_in;
logic cond340_write_en;
logic cond340_clk;
logic cond340_reset;
logic cond340_out;
logic cond340_done;
logic cond_wire340_in;
logic cond_wire340_out;
logic cond341_in;
logic cond341_write_en;
logic cond341_clk;
logic cond341_reset;
logic cond341_out;
logic cond341_done;
logic cond_wire341_in;
logic cond_wire341_out;
logic cond342_in;
logic cond342_write_en;
logic cond342_clk;
logic cond342_reset;
logic cond342_out;
logic cond342_done;
logic cond_wire342_in;
logic cond_wire342_out;
logic cond343_in;
logic cond343_write_en;
logic cond343_clk;
logic cond343_reset;
logic cond343_out;
logic cond343_done;
logic cond_wire343_in;
logic cond_wire343_out;
logic cond344_in;
logic cond344_write_en;
logic cond344_clk;
logic cond344_reset;
logic cond344_out;
logic cond344_done;
logic cond_wire344_in;
logic cond_wire344_out;
logic cond345_in;
logic cond345_write_en;
logic cond345_clk;
logic cond345_reset;
logic cond345_out;
logic cond345_done;
logic cond_wire345_in;
logic cond_wire345_out;
logic cond346_in;
logic cond346_write_en;
logic cond346_clk;
logic cond346_reset;
logic cond346_out;
logic cond346_done;
logic cond_wire346_in;
logic cond_wire346_out;
logic cond347_in;
logic cond347_write_en;
logic cond347_clk;
logic cond347_reset;
logic cond347_out;
logic cond347_done;
logic cond_wire347_in;
logic cond_wire347_out;
logic cond348_in;
logic cond348_write_en;
logic cond348_clk;
logic cond348_reset;
logic cond348_out;
logic cond348_done;
logic cond_wire348_in;
logic cond_wire348_out;
logic cond349_in;
logic cond349_write_en;
logic cond349_clk;
logic cond349_reset;
logic cond349_out;
logic cond349_done;
logic cond_wire349_in;
logic cond_wire349_out;
logic cond350_in;
logic cond350_write_en;
logic cond350_clk;
logic cond350_reset;
logic cond350_out;
logic cond350_done;
logic cond_wire350_in;
logic cond_wire350_out;
logic cond351_in;
logic cond351_write_en;
logic cond351_clk;
logic cond351_reset;
logic cond351_out;
logic cond351_done;
logic cond_wire351_in;
logic cond_wire351_out;
logic cond352_in;
logic cond352_write_en;
logic cond352_clk;
logic cond352_reset;
logic cond352_out;
logic cond352_done;
logic cond_wire352_in;
logic cond_wire352_out;
logic cond353_in;
logic cond353_write_en;
logic cond353_clk;
logic cond353_reset;
logic cond353_out;
logic cond353_done;
logic cond_wire353_in;
logic cond_wire353_out;
logic cond354_in;
logic cond354_write_en;
logic cond354_clk;
logic cond354_reset;
logic cond354_out;
logic cond354_done;
logic cond_wire354_in;
logic cond_wire354_out;
logic cond355_in;
logic cond355_write_en;
logic cond355_clk;
logic cond355_reset;
logic cond355_out;
logic cond355_done;
logic cond_wire355_in;
logic cond_wire355_out;
logic cond356_in;
logic cond356_write_en;
logic cond356_clk;
logic cond356_reset;
logic cond356_out;
logic cond356_done;
logic cond_wire356_in;
logic cond_wire356_out;
logic cond357_in;
logic cond357_write_en;
logic cond357_clk;
logic cond357_reset;
logic cond357_out;
logic cond357_done;
logic cond_wire357_in;
logic cond_wire357_out;
logic cond358_in;
logic cond358_write_en;
logic cond358_clk;
logic cond358_reset;
logic cond358_out;
logic cond358_done;
logic cond_wire358_in;
logic cond_wire358_out;
logic cond359_in;
logic cond359_write_en;
logic cond359_clk;
logic cond359_reset;
logic cond359_out;
logic cond359_done;
logic cond_wire359_in;
logic cond_wire359_out;
logic cond360_in;
logic cond360_write_en;
logic cond360_clk;
logic cond360_reset;
logic cond360_out;
logic cond360_done;
logic cond_wire360_in;
logic cond_wire360_out;
logic cond361_in;
logic cond361_write_en;
logic cond361_clk;
logic cond361_reset;
logic cond361_out;
logic cond361_done;
logic cond_wire361_in;
logic cond_wire361_out;
logic cond362_in;
logic cond362_write_en;
logic cond362_clk;
logic cond362_reset;
logic cond362_out;
logic cond362_done;
logic cond_wire362_in;
logic cond_wire362_out;
logic cond363_in;
logic cond363_write_en;
logic cond363_clk;
logic cond363_reset;
logic cond363_out;
logic cond363_done;
logic cond_wire363_in;
logic cond_wire363_out;
logic cond364_in;
logic cond364_write_en;
logic cond364_clk;
logic cond364_reset;
logic cond364_out;
logic cond364_done;
logic cond_wire364_in;
logic cond_wire364_out;
logic cond365_in;
logic cond365_write_en;
logic cond365_clk;
logic cond365_reset;
logic cond365_out;
logic cond365_done;
logic cond_wire365_in;
logic cond_wire365_out;
logic cond366_in;
logic cond366_write_en;
logic cond366_clk;
logic cond366_reset;
logic cond366_out;
logic cond366_done;
logic cond_wire366_in;
logic cond_wire366_out;
logic cond367_in;
logic cond367_write_en;
logic cond367_clk;
logic cond367_reset;
logic cond367_out;
logic cond367_done;
logic cond_wire367_in;
logic cond_wire367_out;
logic cond368_in;
logic cond368_write_en;
logic cond368_clk;
logic cond368_reset;
logic cond368_out;
logic cond368_done;
logic cond_wire368_in;
logic cond_wire368_out;
logic cond369_in;
logic cond369_write_en;
logic cond369_clk;
logic cond369_reset;
logic cond369_out;
logic cond369_done;
logic cond_wire369_in;
logic cond_wire369_out;
logic cond370_in;
logic cond370_write_en;
logic cond370_clk;
logic cond370_reset;
logic cond370_out;
logic cond370_done;
logic cond_wire370_in;
logic cond_wire370_out;
logic cond371_in;
logic cond371_write_en;
logic cond371_clk;
logic cond371_reset;
logic cond371_out;
logic cond371_done;
logic cond_wire371_in;
logic cond_wire371_out;
logic cond372_in;
logic cond372_write_en;
logic cond372_clk;
logic cond372_reset;
logic cond372_out;
logic cond372_done;
logic cond_wire372_in;
logic cond_wire372_out;
logic cond373_in;
logic cond373_write_en;
logic cond373_clk;
logic cond373_reset;
logic cond373_out;
logic cond373_done;
logic cond_wire373_in;
logic cond_wire373_out;
logic cond374_in;
logic cond374_write_en;
logic cond374_clk;
logic cond374_reset;
logic cond374_out;
logic cond374_done;
logic cond_wire374_in;
logic cond_wire374_out;
logic cond375_in;
logic cond375_write_en;
logic cond375_clk;
logic cond375_reset;
logic cond375_out;
logic cond375_done;
logic cond_wire375_in;
logic cond_wire375_out;
logic cond376_in;
logic cond376_write_en;
logic cond376_clk;
logic cond376_reset;
logic cond376_out;
logic cond376_done;
logic cond_wire376_in;
logic cond_wire376_out;
logic cond377_in;
logic cond377_write_en;
logic cond377_clk;
logic cond377_reset;
logic cond377_out;
logic cond377_done;
logic cond_wire377_in;
logic cond_wire377_out;
logic cond378_in;
logic cond378_write_en;
logic cond378_clk;
logic cond378_reset;
logic cond378_out;
logic cond378_done;
logic cond_wire378_in;
logic cond_wire378_out;
logic cond379_in;
logic cond379_write_en;
logic cond379_clk;
logic cond379_reset;
logic cond379_out;
logic cond379_done;
logic cond_wire379_in;
logic cond_wire379_out;
logic cond380_in;
logic cond380_write_en;
logic cond380_clk;
logic cond380_reset;
logic cond380_out;
logic cond380_done;
logic cond_wire380_in;
logic cond_wire380_out;
logic cond381_in;
logic cond381_write_en;
logic cond381_clk;
logic cond381_reset;
logic cond381_out;
logic cond381_done;
logic cond_wire381_in;
logic cond_wire381_out;
logic cond382_in;
logic cond382_write_en;
logic cond382_clk;
logic cond382_reset;
logic cond382_out;
logic cond382_done;
logic cond_wire382_in;
logic cond_wire382_out;
logic cond383_in;
logic cond383_write_en;
logic cond383_clk;
logic cond383_reset;
logic cond383_out;
logic cond383_done;
logic cond_wire383_in;
logic cond_wire383_out;
logic cond384_in;
logic cond384_write_en;
logic cond384_clk;
logic cond384_reset;
logic cond384_out;
logic cond384_done;
logic cond_wire384_in;
logic cond_wire384_out;
logic cond385_in;
logic cond385_write_en;
logic cond385_clk;
logic cond385_reset;
logic cond385_out;
logic cond385_done;
logic cond_wire385_in;
logic cond_wire385_out;
logic cond386_in;
logic cond386_write_en;
logic cond386_clk;
logic cond386_reset;
logic cond386_out;
logic cond386_done;
logic cond_wire386_in;
logic cond_wire386_out;
logic cond387_in;
logic cond387_write_en;
logic cond387_clk;
logic cond387_reset;
logic cond387_out;
logic cond387_done;
logic cond_wire387_in;
logic cond_wire387_out;
logic cond388_in;
logic cond388_write_en;
logic cond388_clk;
logic cond388_reset;
logic cond388_out;
logic cond388_done;
logic cond_wire388_in;
logic cond_wire388_out;
logic cond389_in;
logic cond389_write_en;
logic cond389_clk;
logic cond389_reset;
logic cond389_out;
logic cond389_done;
logic cond_wire389_in;
logic cond_wire389_out;
logic cond390_in;
logic cond390_write_en;
logic cond390_clk;
logic cond390_reset;
logic cond390_out;
logic cond390_done;
logic cond_wire390_in;
logic cond_wire390_out;
logic cond391_in;
logic cond391_write_en;
logic cond391_clk;
logic cond391_reset;
logic cond391_out;
logic cond391_done;
logic cond_wire391_in;
logic cond_wire391_out;
logic cond392_in;
logic cond392_write_en;
logic cond392_clk;
logic cond392_reset;
logic cond392_out;
logic cond392_done;
logic cond_wire392_in;
logic cond_wire392_out;
logic cond393_in;
logic cond393_write_en;
logic cond393_clk;
logic cond393_reset;
logic cond393_out;
logic cond393_done;
logic cond_wire393_in;
logic cond_wire393_out;
logic cond394_in;
logic cond394_write_en;
logic cond394_clk;
logic cond394_reset;
logic cond394_out;
logic cond394_done;
logic cond_wire394_in;
logic cond_wire394_out;
logic cond395_in;
logic cond395_write_en;
logic cond395_clk;
logic cond395_reset;
logic cond395_out;
logic cond395_done;
logic cond_wire395_in;
logic cond_wire395_out;
logic cond396_in;
logic cond396_write_en;
logic cond396_clk;
logic cond396_reset;
logic cond396_out;
logic cond396_done;
logic cond_wire396_in;
logic cond_wire396_out;
logic cond397_in;
logic cond397_write_en;
logic cond397_clk;
logic cond397_reset;
logic cond397_out;
logic cond397_done;
logic cond_wire397_in;
logic cond_wire397_out;
logic cond398_in;
logic cond398_write_en;
logic cond398_clk;
logic cond398_reset;
logic cond398_out;
logic cond398_done;
logic cond_wire398_in;
logic cond_wire398_out;
logic cond399_in;
logic cond399_write_en;
logic cond399_clk;
logic cond399_reset;
logic cond399_out;
logic cond399_done;
logic cond_wire399_in;
logic cond_wire399_out;
logic cond400_in;
logic cond400_write_en;
logic cond400_clk;
logic cond400_reset;
logic cond400_out;
logic cond400_done;
logic cond_wire400_in;
logic cond_wire400_out;
logic cond401_in;
logic cond401_write_en;
logic cond401_clk;
logic cond401_reset;
logic cond401_out;
logic cond401_done;
logic cond_wire401_in;
logic cond_wire401_out;
logic cond402_in;
logic cond402_write_en;
logic cond402_clk;
logic cond402_reset;
logic cond402_out;
logic cond402_done;
logic cond_wire402_in;
logic cond_wire402_out;
logic cond403_in;
logic cond403_write_en;
logic cond403_clk;
logic cond403_reset;
logic cond403_out;
logic cond403_done;
logic cond_wire403_in;
logic cond_wire403_out;
logic cond404_in;
logic cond404_write_en;
logic cond404_clk;
logic cond404_reset;
logic cond404_out;
logic cond404_done;
logic cond_wire404_in;
logic cond_wire404_out;
logic cond405_in;
logic cond405_write_en;
logic cond405_clk;
logic cond405_reset;
logic cond405_out;
logic cond405_done;
logic cond_wire405_in;
logic cond_wire405_out;
logic cond406_in;
logic cond406_write_en;
logic cond406_clk;
logic cond406_reset;
logic cond406_out;
logic cond406_done;
logic cond_wire406_in;
logic cond_wire406_out;
logic cond407_in;
logic cond407_write_en;
logic cond407_clk;
logic cond407_reset;
logic cond407_out;
logic cond407_done;
logic cond_wire407_in;
logic cond_wire407_out;
logic cond408_in;
logic cond408_write_en;
logic cond408_clk;
logic cond408_reset;
logic cond408_out;
logic cond408_done;
logic cond_wire408_in;
logic cond_wire408_out;
logic cond409_in;
logic cond409_write_en;
logic cond409_clk;
logic cond409_reset;
logic cond409_out;
logic cond409_done;
logic cond_wire409_in;
logic cond_wire409_out;
logic cond410_in;
logic cond410_write_en;
logic cond410_clk;
logic cond410_reset;
logic cond410_out;
logic cond410_done;
logic cond_wire410_in;
logic cond_wire410_out;
logic cond411_in;
logic cond411_write_en;
logic cond411_clk;
logic cond411_reset;
logic cond411_out;
logic cond411_done;
logic cond_wire411_in;
logic cond_wire411_out;
logic cond412_in;
logic cond412_write_en;
logic cond412_clk;
logic cond412_reset;
logic cond412_out;
logic cond412_done;
logic cond_wire412_in;
logic cond_wire412_out;
logic cond413_in;
logic cond413_write_en;
logic cond413_clk;
logic cond413_reset;
logic cond413_out;
logic cond413_done;
logic cond_wire413_in;
logic cond_wire413_out;
logic cond414_in;
logic cond414_write_en;
logic cond414_clk;
logic cond414_reset;
logic cond414_out;
logic cond414_done;
logic cond_wire414_in;
logic cond_wire414_out;
logic cond415_in;
logic cond415_write_en;
logic cond415_clk;
logic cond415_reset;
logic cond415_out;
logic cond415_done;
logic cond_wire415_in;
logic cond_wire415_out;
logic cond416_in;
logic cond416_write_en;
logic cond416_clk;
logic cond416_reset;
logic cond416_out;
logic cond416_done;
logic cond_wire416_in;
logic cond_wire416_out;
logic cond417_in;
logic cond417_write_en;
logic cond417_clk;
logic cond417_reset;
logic cond417_out;
logic cond417_done;
logic cond_wire417_in;
logic cond_wire417_out;
logic cond418_in;
logic cond418_write_en;
logic cond418_clk;
logic cond418_reset;
logic cond418_out;
logic cond418_done;
logic cond_wire418_in;
logic cond_wire418_out;
logic cond419_in;
logic cond419_write_en;
logic cond419_clk;
logic cond419_reset;
logic cond419_out;
logic cond419_done;
logic cond_wire419_in;
logic cond_wire419_out;
logic cond420_in;
logic cond420_write_en;
logic cond420_clk;
logic cond420_reset;
logic cond420_out;
logic cond420_done;
logic cond_wire420_in;
logic cond_wire420_out;
logic cond421_in;
logic cond421_write_en;
logic cond421_clk;
logic cond421_reset;
logic cond421_out;
logic cond421_done;
logic cond_wire421_in;
logic cond_wire421_out;
logic cond422_in;
logic cond422_write_en;
logic cond422_clk;
logic cond422_reset;
logic cond422_out;
logic cond422_done;
logic cond_wire422_in;
logic cond_wire422_out;
logic cond423_in;
logic cond423_write_en;
logic cond423_clk;
logic cond423_reset;
logic cond423_out;
logic cond423_done;
logic cond_wire423_in;
logic cond_wire423_out;
logic cond424_in;
logic cond424_write_en;
logic cond424_clk;
logic cond424_reset;
logic cond424_out;
logic cond424_done;
logic cond_wire424_in;
logic cond_wire424_out;
logic cond425_in;
logic cond425_write_en;
logic cond425_clk;
logic cond425_reset;
logic cond425_out;
logic cond425_done;
logic cond_wire425_in;
logic cond_wire425_out;
logic cond426_in;
logic cond426_write_en;
logic cond426_clk;
logic cond426_reset;
logic cond426_out;
logic cond426_done;
logic cond_wire426_in;
logic cond_wire426_out;
logic cond427_in;
logic cond427_write_en;
logic cond427_clk;
logic cond427_reset;
logic cond427_out;
logic cond427_done;
logic cond_wire427_in;
logic cond_wire427_out;
logic cond428_in;
logic cond428_write_en;
logic cond428_clk;
logic cond428_reset;
logic cond428_out;
logic cond428_done;
logic cond_wire428_in;
logic cond_wire428_out;
logic cond429_in;
logic cond429_write_en;
logic cond429_clk;
logic cond429_reset;
logic cond429_out;
logic cond429_done;
logic cond_wire429_in;
logic cond_wire429_out;
logic cond430_in;
logic cond430_write_en;
logic cond430_clk;
logic cond430_reset;
logic cond430_out;
logic cond430_done;
logic cond_wire430_in;
logic cond_wire430_out;
logic cond431_in;
logic cond431_write_en;
logic cond431_clk;
logic cond431_reset;
logic cond431_out;
logic cond431_done;
logic cond_wire431_in;
logic cond_wire431_out;
logic cond432_in;
logic cond432_write_en;
logic cond432_clk;
logic cond432_reset;
logic cond432_out;
logic cond432_done;
logic cond_wire432_in;
logic cond_wire432_out;
logic cond433_in;
logic cond433_write_en;
logic cond433_clk;
logic cond433_reset;
logic cond433_out;
logic cond433_done;
logic cond_wire433_in;
logic cond_wire433_out;
logic cond434_in;
logic cond434_write_en;
logic cond434_clk;
logic cond434_reset;
logic cond434_out;
logic cond434_done;
logic cond_wire434_in;
logic cond_wire434_out;
logic cond435_in;
logic cond435_write_en;
logic cond435_clk;
logic cond435_reset;
logic cond435_out;
logic cond435_done;
logic cond_wire435_in;
logic cond_wire435_out;
logic cond436_in;
logic cond436_write_en;
logic cond436_clk;
logic cond436_reset;
logic cond436_out;
logic cond436_done;
logic cond_wire436_in;
logic cond_wire436_out;
logic cond437_in;
logic cond437_write_en;
logic cond437_clk;
logic cond437_reset;
logic cond437_out;
logic cond437_done;
logic cond_wire437_in;
logic cond_wire437_out;
logic cond438_in;
logic cond438_write_en;
logic cond438_clk;
logic cond438_reset;
logic cond438_out;
logic cond438_done;
logic cond_wire438_in;
logic cond_wire438_out;
logic cond439_in;
logic cond439_write_en;
logic cond439_clk;
logic cond439_reset;
logic cond439_out;
logic cond439_done;
logic cond_wire439_in;
logic cond_wire439_out;
logic cond440_in;
logic cond440_write_en;
logic cond440_clk;
logic cond440_reset;
logic cond440_out;
logic cond440_done;
logic cond_wire440_in;
logic cond_wire440_out;
logic cond441_in;
logic cond441_write_en;
logic cond441_clk;
logic cond441_reset;
logic cond441_out;
logic cond441_done;
logic cond_wire441_in;
logic cond_wire441_out;
logic cond442_in;
logic cond442_write_en;
logic cond442_clk;
logic cond442_reset;
logic cond442_out;
logic cond442_done;
logic cond_wire442_in;
logic cond_wire442_out;
logic cond443_in;
logic cond443_write_en;
logic cond443_clk;
logic cond443_reset;
logic cond443_out;
logic cond443_done;
logic cond_wire443_in;
logic cond_wire443_out;
logic cond444_in;
logic cond444_write_en;
logic cond444_clk;
logic cond444_reset;
logic cond444_out;
logic cond444_done;
logic cond_wire444_in;
logic cond_wire444_out;
logic cond445_in;
logic cond445_write_en;
logic cond445_clk;
logic cond445_reset;
logic cond445_out;
logic cond445_done;
logic cond_wire445_in;
logic cond_wire445_out;
logic cond446_in;
logic cond446_write_en;
logic cond446_clk;
logic cond446_reset;
logic cond446_out;
logic cond446_done;
logic cond_wire446_in;
logic cond_wire446_out;
logic cond447_in;
logic cond447_write_en;
logic cond447_clk;
logic cond447_reset;
logic cond447_out;
logic cond447_done;
logic cond_wire447_in;
logic cond_wire447_out;
logic cond448_in;
logic cond448_write_en;
logic cond448_clk;
logic cond448_reset;
logic cond448_out;
logic cond448_done;
logic cond_wire448_in;
logic cond_wire448_out;
logic cond449_in;
logic cond449_write_en;
logic cond449_clk;
logic cond449_reset;
logic cond449_out;
logic cond449_done;
logic cond_wire449_in;
logic cond_wire449_out;
logic cond450_in;
logic cond450_write_en;
logic cond450_clk;
logic cond450_reset;
logic cond450_out;
logic cond450_done;
logic cond_wire450_in;
logic cond_wire450_out;
logic cond451_in;
logic cond451_write_en;
logic cond451_clk;
logic cond451_reset;
logic cond451_out;
logic cond451_done;
logic cond_wire451_in;
logic cond_wire451_out;
logic cond452_in;
logic cond452_write_en;
logic cond452_clk;
logic cond452_reset;
logic cond452_out;
logic cond452_done;
logic cond_wire452_in;
logic cond_wire452_out;
logic cond453_in;
logic cond453_write_en;
logic cond453_clk;
logic cond453_reset;
logic cond453_out;
logic cond453_done;
logic cond_wire453_in;
logic cond_wire453_out;
logic cond454_in;
logic cond454_write_en;
logic cond454_clk;
logic cond454_reset;
logic cond454_out;
logic cond454_done;
logic cond_wire454_in;
logic cond_wire454_out;
logic cond455_in;
logic cond455_write_en;
logic cond455_clk;
logic cond455_reset;
logic cond455_out;
logic cond455_done;
logic cond_wire455_in;
logic cond_wire455_out;
logic cond456_in;
logic cond456_write_en;
logic cond456_clk;
logic cond456_reset;
logic cond456_out;
logic cond456_done;
logic cond_wire456_in;
logic cond_wire456_out;
logic cond457_in;
logic cond457_write_en;
logic cond457_clk;
logic cond457_reset;
logic cond457_out;
logic cond457_done;
logic cond_wire457_in;
logic cond_wire457_out;
logic cond458_in;
logic cond458_write_en;
logic cond458_clk;
logic cond458_reset;
logic cond458_out;
logic cond458_done;
logic cond_wire458_in;
logic cond_wire458_out;
logic cond459_in;
logic cond459_write_en;
logic cond459_clk;
logic cond459_reset;
logic cond459_out;
logic cond459_done;
logic cond_wire459_in;
logic cond_wire459_out;
logic cond460_in;
logic cond460_write_en;
logic cond460_clk;
logic cond460_reset;
logic cond460_out;
logic cond460_done;
logic cond_wire460_in;
logic cond_wire460_out;
logic cond461_in;
logic cond461_write_en;
logic cond461_clk;
logic cond461_reset;
logic cond461_out;
logic cond461_done;
logic cond_wire461_in;
logic cond_wire461_out;
logic cond462_in;
logic cond462_write_en;
logic cond462_clk;
logic cond462_reset;
logic cond462_out;
logic cond462_done;
logic cond_wire462_in;
logic cond_wire462_out;
logic cond463_in;
logic cond463_write_en;
logic cond463_clk;
logic cond463_reset;
logic cond463_out;
logic cond463_done;
logic cond_wire463_in;
logic cond_wire463_out;
logic cond464_in;
logic cond464_write_en;
logic cond464_clk;
logic cond464_reset;
logic cond464_out;
logic cond464_done;
logic cond_wire464_in;
logic cond_wire464_out;
logic cond465_in;
logic cond465_write_en;
logic cond465_clk;
logic cond465_reset;
logic cond465_out;
logic cond465_done;
logic cond_wire465_in;
logic cond_wire465_out;
logic cond466_in;
logic cond466_write_en;
logic cond466_clk;
logic cond466_reset;
logic cond466_out;
logic cond466_done;
logic cond_wire466_in;
logic cond_wire466_out;
logic cond467_in;
logic cond467_write_en;
logic cond467_clk;
logic cond467_reset;
logic cond467_out;
logic cond467_done;
logic cond_wire467_in;
logic cond_wire467_out;
logic cond468_in;
logic cond468_write_en;
logic cond468_clk;
logic cond468_reset;
logic cond468_out;
logic cond468_done;
logic cond_wire468_in;
logic cond_wire468_out;
logic cond469_in;
logic cond469_write_en;
logic cond469_clk;
logic cond469_reset;
logic cond469_out;
logic cond469_done;
logic cond_wire469_in;
logic cond_wire469_out;
logic cond470_in;
logic cond470_write_en;
logic cond470_clk;
logic cond470_reset;
logic cond470_out;
logic cond470_done;
logic cond_wire470_in;
logic cond_wire470_out;
logic cond471_in;
logic cond471_write_en;
logic cond471_clk;
logic cond471_reset;
logic cond471_out;
logic cond471_done;
logic cond_wire471_in;
logic cond_wire471_out;
logic cond472_in;
logic cond472_write_en;
logic cond472_clk;
logic cond472_reset;
logic cond472_out;
logic cond472_done;
logic cond_wire472_in;
logic cond_wire472_out;
logic cond473_in;
logic cond473_write_en;
logic cond473_clk;
logic cond473_reset;
logic cond473_out;
logic cond473_done;
logic cond_wire473_in;
logic cond_wire473_out;
logic cond474_in;
logic cond474_write_en;
logic cond474_clk;
logic cond474_reset;
logic cond474_out;
logic cond474_done;
logic cond_wire474_in;
logic cond_wire474_out;
logic cond475_in;
logic cond475_write_en;
logic cond475_clk;
logic cond475_reset;
logic cond475_out;
logic cond475_done;
logic cond_wire475_in;
logic cond_wire475_out;
logic cond476_in;
logic cond476_write_en;
logic cond476_clk;
logic cond476_reset;
logic cond476_out;
logic cond476_done;
logic cond_wire476_in;
logic cond_wire476_out;
logic cond477_in;
logic cond477_write_en;
logic cond477_clk;
logic cond477_reset;
logic cond477_out;
logic cond477_done;
logic cond_wire477_in;
logic cond_wire477_out;
logic cond478_in;
logic cond478_write_en;
logic cond478_clk;
logic cond478_reset;
logic cond478_out;
logic cond478_done;
logic cond_wire478_in;
logic cond_wire478_out;
logic cond479_in;
logic cond479_write_en;
logic cond479_clk;
logic cond479_reset;
logic cond479_out;
logic cond479_done;
logic cond_wire479_in;
logic cond_wire479_out;
logic cond480_in;
logic cond480_write_en;
logic cond480_clk;
logic cond480_reset;
logic cond480_out;
logic cond480_done;
logic cond_wire480_in;
logic cond_wire480_out;
logic cond481_in;
logic cond481_write_en;
logic cond481_clk;
logic cond481_reset;
logic cond481_out;
logic cond481_done;
logic cond_wire481_in;
logic cond_wire481_out;
logic cond482_in;
logic cond482_write_en;
logic cond482_clk;
logic cond482_reset;
logic cond482_out;
logic cond482_done;
logic cond_wire482_in;
logic cond_wire482_out;
logic cond483_in;
logic cond483_write_en;
logic cond483_clk;
logic cond483_reset;
logic cond483_out;
logic cond483_done;
logic cond_wire483_in;
logic cond_wire483_out;
logic cond484_in;
logic cond484_write_en;
logic cond484_clk;
logic cond484_reset;
logic cond484_out;
logic cond484_done;
logic cond_wire484_in;
logic cond_wire484_out;
logic cond485_in;
logic cond485_write_en;
logic cond485_clk;
logic cond485_reset;
logic cond485_out;
logic cond485_done;
logic cond_wire485_in;
logic cond_wire485_out;
logic cond486_in;
logic cond486_write_en;
logic cond486_clk;
logic cond486_reset;
logic cond486_out;
logic cond486_done;
logic cond_wire486_in;
logic cond_wire486_out;
logic cond487_in;
logic cond487_write_en;
logic cond487_clk;
logic cond487_reset;
logic cond487_out;
logic cond487_done;
logic cond_wire487_in;
logic cond_wire487_out;
logic cond488_in;
logic cond488_write_en;
logic cond488_clk;
logic cond488_reset;
logic cond488_out;
logic cond488_done;
logic cond_wire488_in;
logic cond_wire488_out;
logic cond489_in;
logic cond489_write_en;
logic cond489_clk;
logic cond489_reset;
logic cond489_out;
logic cond489_done;
logic cond_wire489_in;
logic cond_wire489_out;
logic cond490_in;
logic cond490_write_en;
logic cond490_clk;
logic cond490_reset;
logic cond490_out;
logic cond490_done;
logic cond_wire490_in;
logic cond_wire490_out;
logic cond491_in;
logic cond491_write_en;
logic cond491_clk;
logic cond491_reset;
logic cond491_out;
logic cond491_done;
logic cond_wire491_in;
logic cond_wire491_out;
logic cond492_in;
logic cond492_write_en;
logic cond492_clk;
logic cond492_reset;
logic cond492_out;
logic cond492_done;
logic cond_wire492_in;
logic cond_wire492_out;
logic cond493_in;
logic cond493_write_en;
logic cond493_clk;
logic cond493_reset;
logic cond493_out;
logic cond493_done;
logic cond_wire493_in;
logic cond_wire493_out;
logic cond494_in;
logic cond494_write_en;
logic cond494_clk;
logic cond494_reset;
logic cond494_out;
logic cond494_done;
logic cond_wire494_in;
logic cond_wire494_out;
logic cond495_in;
logic cond495_write_en;
logic cond495_clk;
logic cond495_reset;
logic cond495_out;
logic cond495_done;
logic cond_wire495_in;
logic cond_wire495_out;
logic cond496_in;
logic cond496_write_en;
logic cond496_clk;
logic cond496_reset;
logic cond496_out;
logic cond496_done;
logic cond_wire496_in;
logic cond_wire496_out;
logic cond497_in;
logic cond497_write_en;
logic cond497_clk;
logic cond497_reset;
logic cond497_out;
logic cond497_done;
logic cond_wire497_in;
logic cond_wire497_out;
logic cond498_in;
logic cond498_write_en;
logic cond498_clk;
logic cond498_reset;
logic cond498_out;
logic cond498_done;
logic cond_wire498_in;
logic cond_wire498_out;
logic cond499_in;
logic cond499_write_en;
logic cond499_clk;
logic cond499_reset;
logic cond499_out;
logic cond499_done;
logic cond_wire499_in;
logic cond_wire499_out;
logic cond500_in;
logic cond500_write_en;
logic cond500_clk;
logic cond500_reset;
logic cond500_out;
logic cond500_done;
logic cond_wire500_in;
logic cond_wire500_out;
logic cond501_in;
logic cond501_write_en;
logic cond501_clk;
logic cond501_reset;
logic cond501_out;
logic cond501_done;
logic cond_wire501_in;
logic cond_wire501_out;
logic cond502_in;
logic cond502_write_en;
logic cond502_clk;
logic cond502_reset;
logic cond502_out;
logic cond502_done;
logic cond_wire502_in;
logic cond_wire502_out;
logic cond503_in;
logic cond503_write_en;
logic cond503_clk;
logic cond503_reset;
logic cond503_out;
logic cond503_done;
logic cond_wire503_in;
logic cond_wire503_out;
logic cond504_in;
logic cond504_write_en;
logic cond504_clk;
logic cond504_reset;
logic cond504_out;
logic cond504_done;
logic cond_wire504_in;
logic cond_wire504_out;
logic cond505_in;
logic cond505_write_en;
logic cond505_clk;
logic cond505_reset;
logic cond505_out;
logic cond505_done;
logic cond_wire505_in;
logic cond_wire505_out;
logic cond506_in;
logic cond506_write_en;
logic cond506_clk;
logic cond506_reset;
logic cond506_out;
logic cond506_done;
logic cond_wire506_in;
logic cond_wire506_out;
logic cond507_in;
logic cond507_write_en;
logic cond507_clk;
logic cond507_reset;
logic cond507_out;
logic cond507_done;
logic cond_wire507_in;
logic cond_wire507_out;
logic cond508_in;
logic cond508_write_en;
logic cond508_clk;
logic cond508_reset;
logic cond508_out;
logic cond508_done;
logic cond_wire508_in;
logic cond_wire508_out;
logic cond509_in;
logic cond509_write_en;
logic cond509_clk;
logic cond509_reset;
logic cond509_out;
logic cond509_done;
logic cond_wire509_in;
logic cond_wire509_out;
logic cond510_in;
logic cond510_write_en;
logic cond510_clk;
logic cond510_reset;
logic cond510_out;
logic cond510_done;
logic cond_wire510_in;
logic cond_wire510_out;
logic cond511_in;
logic cond511_write_en;
logic cond511_clk;
logic cond511_reset;
logic cond511_out;
logic cond511_done;
logic cond_wire511_in;
logic cond_wire511_out;
logic cond512_in;
logic cond512_write_en;
logic cond512_clk;
logic cond512_reset;
logic cond512_out;
logic cond512_done;
logic cond_wire512_in;
logic cond_wire512_out;
logic cond513_in;
logic cond513_write_en;
logic cond513_clk;
logic cond513_reset;
logic cond513_out;
logic cond513_done;
logic cond_wire513_in;
logic cond_wire513_out;
logic cond514_in;
logic cond514_write_en;
logic cond514_clk;
logic cond514_reset;
logic cond514_out;
logic cond514_done;
logic cond_wire514_in;
logic cond_wire514_out;
logic cond515_in;
logic cond515_write_en;
logic cond515_clk;
logic cond515_reset;
logic cond515_out;
logic cond515_done;
logic cond_wire515_in;
logic cond_wire515_out;
logic cond516_in;
logic cond516_write_en;
logic cond516_clk;
logic cond516_reset;
logic cond516_out;
logic cond516_done;
logic cond_wire516_in;
logic cond_wire516_out;
logic cond517_in;
logic cond517_write_en;
logic cond517_clk;
logic cond517_reset;
logic cond517_out;
logic cond517_done;
logic cond_wire517_in;
logic cond_wire517_out;
logic cond518_in;
logic cond518_write_en;
logic cond518_clk;
logic cond518_reset;
logic cond518_out;
logic cond518_done;
logic cond_wire518_in;
logic cond_wire518_out;
logic cond519_in;
logic cond519_write_en;
logic cond519_clk;
logic cond519_reset;
logic cond519_out;
logic cond519_done;
logic cond_wire519_in;
logic cond_wire519_out;
logic cond520_in;
logic cond520_write_en;
logic cond520_clk;
logic cond520_reset;
logic cond520_out;
logic cond520_done;
logic cond_wire520_in;
logic cond_wire520_out;
logic cond521_in;
logic cond521_write_en;
logic cond521_clk;
logic cond521_reset;
logic cond521_out;
logic cond521_done;
logic cond_wire521_in;
logic cond_wire521_out;
logic cond522_in;
logic cond522_write_en;
logic cond522_clk;
logic cond522_reset;
logic cond522_out;
logic cond522_done;
logic cond_wire522_in;
logic cond_wire522_out;
logic cond523_in;
logic cond523_write_en;
logic cond523_clk;
logic cond523_reset;
logic cond523_out;
logic cond523_done;
logic cond_wire523_in;
logic cond_wire523_out;
logic cond524_in;
logic cond524_write_en;
logic cond524_clk;
logic cond524_reset;
logic cond524_out;
logic cond524_done;
logic cond_wire524_in;
logic cond_wire524_out;
logic cond525_in;
logic cond525_write_en;
logic cond525_clk;
logic cond525_reset;
logic cond525_out;
logic cond525_done;
logic cond_wire525_in;
logic cond_wire525_out;
logic cond526_in;
logic cond526_write_en;
logic cond526_clk;
logic cond526_reset;
logic cond526_out;
logic cond526_done;
logic cond_wire526_in;
logic cond_wire526_out;
logic cond527_in;
logic cond527_write_en;
logic cond527_clk;
logic cond527_reset;
logic cond527_out;
logic cond527_done;
logic cond_wire527_in;
logic cond_wire527_out;
logic cond528_in;
logic cond528_write_en;
logic cond528_clk;
logic cond528_reset;
logic cond528_out;
logic cond528_done;
logic cond_wire528_in;
logic cond_wire528_out;
logic cond529_in;
logic cond529_write_en;
logic cond529_clk;
logic cond529_reset;
logic cond529_out;
logic cond529_done;
logic cond_wire529_in;
logic cond_wire529_out;
logic cond530_in;
logic cond530_write_en;
logic cond530_clk;
logic cond530_reset;
logic cond530_out;
logic cond530_done;
logic cond_wire530_in;
logic cond_wire530_out;
logic cond531_in;
logic cond531_write_en;
logic cond531_clk;
logic cond531_reset;
logic cond531_out;
logic cond531_done;
logic cond_wire531_in;
logic cond_wire531_out;
logic cond532_in;
logic cond532_write_en;
logic cond532_clk;
logic cond532_reset;
logic cond532_out;
logic cond532_done;
logic cond_wire532_in;
logic cond_wire532_out;
logic cond533_in;
logic cond533_write_en;
logic cond533_clk;
logic cond533_reset;
logic cond533_out;
logic cond533_done;
logic cond_wire533_in;
logic cond_wire533_out;
logic cond534_in;
logic cond534_write_en;
logic cond534_clk;
logic cond534_reset;
logic cond534_out;
logic cond534_done;
logic cond_wire534_in;
logic cond_wire534_out;
logic cond535_in;
logic cond535_write_en;
logic cond535_clk;
logic cond535_reset;
logic cond535_out;
logic cond535_done;
logic cond_wire535_in;
logic cond_wire535_out;
logic cond536_in;
logic cond536_write_en;
logic cond536_clk;
logic cond536_reset;
logic cond536_out;
logic cond536_done;
logic cond_wire536_in;
logic cond_wire536_out;
logic cond537_in;
logic cond537_write_en;
logic cond537_clk;
logic cond537_reset;
logic cond537_out;
logic cond537_done;
logic cond_wire537_in;
logic cond_wire537_out;
logic cond538_in;
logic cond538_write_en;
logic cond538_clk;
logic cond538_reset;
logic cond538_out;
logic cond538_done;
logic cond_wire538_in;
logic cond_wire538_out;
logic cond539_in;
logic cond539_write_en;
logic cond539_clk;
logic cond539_reset;
logic cond539_out;
logic cond539_done;
logic cond_wire539_in;
logic cond_wire539_out;
logic cond540_in;
logic cond540_write_en;
logic cond540_clk;
logic cond540_reset;
logic cond540_out;
logic cond540_done;
logic cond_wire540_in;
logic cond_wire540_out;
logic cond541_in;
logic cond541_write_en;
logic cond541_clk;
logic cond541_reset;
logic cond541_out;
logic cond541_done;
logic cond_wire541_in;
logic cond_wire541_out;
logic cond542_in;
logic cond542_write_en;
logic cond542_clk;
logic cond542_reset;
logic cond542_out;
logic cond542_done;
logic cond_wire542_in;
logic cond_wire542_out;
logic cond543_in;
logic cond543_write_en;
logic cond543_clk;
logic cond543_reset;
logic cond543_out;
logic cond543_done;
logic cond_wire543_in;
logic cond_wire543_out;
logic cond544_in;
logic cond544_write_en;
logic cond544_clk;
logic cond544_reset;
logic cond544_out;
logic cond544_done;
logic cond_wire544_in;
logic cond_wire544_out;
logic cond545_in;
logic cond545_write_en;
logic cond545_clk;
logic cond545_reset;
logic cond545_out;
logic cond545_done;
logic cond_wire545_in;
logic cond_wire545_out;
logic cond546_in;
logic cond546_write_en;
logic cond546_clk;
logic cond546_reset;
logic cond546_out;
logic cond546_done;
logic cond_wire546_in;
logic cond_wire546_out;
logic cond547_in;
logic cond547_write_en;
logic cond547_clk;
logic cond547_reset;
logic cond547_out;
logic cond547_done;
logic cond_wire547_in;
logic cond_wire547_out;
logic cond548_in;
logic cond548_write_en;
logic cond548_clk;
logic cond548_reset;
logic cond548_out;
logic cond548_done;
logic cond_wire548_in;
logic cond_wire548_out;
logic cond549_in;
logic cond549_write_en;
logic cond549_clk;
logic cond549_reset;
logic cond549_out;
logic cond549_done;
logic cond_wire549_in;
logic cond_wire549_out;
logic cond550_in;
logic cond550_write_en;
logic cond550_clk;
logic cond550_reset;
logic cond550_out;
logic cond550_done;
logic cond_wire550_in;
logic cond_wire550_out;
logic cond551_in;
logic cond551_write_en;
logic cond551_clk;
logic cond551_reset;
logic cond551_out;
logic cond551_done;
logic cond_wire551_in;
logic cond_wire551_out;
logic cond552_in;
logic cond552_write_en;
logic cond552_clk;
logic cond552_reset;
logic cond552_out;
logic cond552_done;
logic cond_wire552_in;
logic cond_wire552_out;
logic cond553_in;
logic cond553_write_en;
logic cond553_clk;
logic cond553_reset;
logic cond553_out;
logic cond553_done;
logic cond_wire553_in;
logic cond_wire553_out;
logic cond554_in;
logic cond554_write_en;
logic cond554_clk;
logic cond554_reset;
logic cond554_out;
logic cond554_done;
logic cond_wire554_in;
logic cond_wire554_out;
logic cond555_in;
logic cond555_write_en;
logic cond555_clk;
logic cond555_reset;
logic cond555_out;
logic cond555_done;
logic cond_wire555_in;
logic cond_wire555_out;
logic cond556_in;
logic cond556_write_en;
logic cond556_clk;
logic cond556_reset;
logic cond556_out;
logic cond556_done;
logic cond_wire556_in;
logic cond_wire556_out;
logic cond557_in;
logic cond557_write_en;
logic cond557_clk;
logic cond557_reset;
logic cond557_out;
logic cond557_done;
logic cond_wire557_in;
logic cond_wire557_out;
logic cond558_in;
logic cond558_write_en;
logic cond558_clk;
logic cond558_reset;
logic cond558_out;
logic cond558_done;
logic cond_wire558_in;
logic cond_wire558_out;
logic cond559_in;
logic cond559_write_en;
logic cond559_clk;
logic cond559_reset;
logic cond559_out;
logic cond559_done;
logic cond_wire559_in;
logic cond_wire559_out;
logic cond560_in;
logic cond560_write_en;
logic cond560_clk;
logic cond560_reset;
logic cond560_out;
logic cond560_done;
logic cond_wire560_in;
logic cond_wire560_out;
logic cond561_in;
logic cond561_write_en;
logic cond561_clk;
logic cond561_reset;
logic cond561_out;
logic cond561_done;
logic cond_wire561_in;
logic cond_wire561_out;
logic cond562_in;
logic cond562_write_en;
logic cond562_clk;
logic cond562_reset;
logic cond562_out;
logic cond562_done;
logic cond_wire562_in;
logic cond_wire562_out;
logic cond563_in;
logic cond563_write_en;
logic cond563_clk;
logic cond563_reset;
logic cond563_out;
logic cond563_done;
logic cond_wire563_in;
logic cond_wire563_out;
logic cond564_in;
logic cond564_write_en;
logic cond564_clk;
logic cond564_reset;
logic cond564_out;
logic cond564_done;
logic cond_wire564_in;
logic cond_wire564_out;
logic cond565_in;
logic cond565_write_en;
logic cond565_clk;
logic cond565_reset;
logic cond565_out;
logic cond565_done;
logic cond_wire565_in;
logic cond_wire565_out;
logic cond566_in;
logic cond566_write_en;
logic cond566_clk;
logic cond566_reset;
logic cond566_out;
logic cond566_done;
logic cond_wire566_in;
logic cond_wire566_out;
logic cond567_in;
logic cond567_write_en;
logic cond567_clk;
logic cond567_reset;
logic cond567_out;
logic cond567_done;
logic cond_wire567_in;
logic cond_wire567_out;
logic cond568_in;
logic cond568_write_en;
logic cond568_clk;
logic cond568_reset;
logic cond568_out;
logic cond568_done;
logic cond_wire568_in;
logic cond_wire568_out;
logic cond569_in;
logic cond569_write_en;
logic cond569_clk;
logic cond569_reset;
logic cond569_out;
logic cond569_done;
logic cond_wire569_in;
logic cond_wire569_out;
logic cond570_in;
logic cond570_write_en;
logic cond570_clk;
logic cond570_reset;
logic cond570_out;
logic cond570_done;
logic cond_wire570_in;
logic cond_wire570_out;
logic cond571_in;
logic cond571_write_en;
logic cond571_clk;
logic cond571_reset;
logic cond571_out;
logic cond571_done;
logic cond_wire571_in;
logic cond_wire571_out;
logic cond572_in;
logic cond572_write_en;
logic cond572_clk;
logic cond572_reset;
logic cond572_out;
logic cond572_done;
logic cond_wire572_in;
logic cond_wire572_out;
logic cond573_in;
logic cond573_write_en;
logic cond573_clk;
logic cond573_reset;
logic cond573_out;
logic cond573_done;
logic cond_wire573_in;
logic cond_wire573_out;
logic cond574_in;
logic cond574_write_en;
logic cond574_clk;
logic cond574_reset;
logic cond574_out;
logic cond574_done;
logic cond_wire574_in;
logic cond_wire574_out;
logic cond575_in;
logic cond575_write_en;
logic cond575_clk;
logic cond575_reset;
logic cond575_out;
logic cond575_done;
logic cond_wire575_in;
logic cond_wire575_out;
logic cond576_in;
logic cond576_write_en;
logic cond576_clk;
logic cond576_reset;
logic cond576_out;
logic cond576_done;
logic cond_wire576_in;
logic cond_wire576_out;
logic cond577_in;
logic cond577_write_en;
logic cond577_clk;
logic cond577_reset;
logic cond577_out;
logic cond577_done;
logic cond_wire577_in;
logic cond_wire577_out;
logic cond578_in;
logic cond578_write_en;
logic cond578_clk;
logic cond578_reset;
logic cond578_out;
logic cond578_done;
logic cond_wire578_in;
logic cond_wire578_out;
logic cond579_in;
logic cond579_write_en;
logic cond579_clk;
logic cond579_reset;
logic cond579_out;
logic cond579_done;
logic cond_wire579_in;
logic cond_wire579_out;
logic cond580_in;
logic cond580_write_en;
logic cond580_clk;
logic cond580_reset;
logic cond580_out;
logic cond580_done;
logic cond_wire580_in;
logic cond_wire580_out;
logic cond581_in;
logic cond581_write_en;
logic cond581_clk;
logic cond581_reset;
logic cond581_out;
logic cond581_done;
logic cond_wire581_in;
logic cond_wire581_out;
logic cond582_in;
logic cond582_write_en;
logic cond582_clk;
logic cond582_reset;
logic cond582_out;
logic cond582_done;
logic cond_wire582_in;
logic cond_wire582_out;
logic cond583_in;
logic cond583_write_en;
logic cond583_clk;
logic cond583_reset;
logic cond583_out;
logic cond583_done;
logic cond_wire583_in;
logic cond_wire583_out;
logic cond584_in;
logic cond584_write_en;
logic cond584_clk;
logic cond584_reset;
logic cond584_out;
logic cond584_done;
logic cond_wire584_in;
logic cond_wire584_out;
logic cond585_in;
logic cond585_write_en;
logic cond585_clk;
logic cond585_reset;
logic cond585_out;
logic cond585_done;
logic cond_wire585_in;
logic cond_wire585_out;
logic cond586_in;
logic cond586_write_en;
logic cond586_clk;
logic cond586_reset;
logic cond586_out;
logic cond586_done;
logic cond_wire586_in;
logic cond_wire586_out;
logic cond587_in;
logic cond587_write_en;
logic cond587_clk;
logic cond587_reset;
logic cond587_out;
logic cond587_done;
logic cond_wire587_in;
logic cond_wire587_out;
logic cond588_in;
logic cond588_write_en;
logic cond588_clk;
logic cond588_reset;
logic cond588_out;
logic cond588_done;
logic cond_wire588_in;
logic cond_wire588_out;
logic cond589_in;
logic cond589_write_en;
logic cond589_clk;
logic cond589_reset;
logic cond589_out;
logic cond589_done;
logic cond_wire589_in;
logic cond_wire589_out;
logic cond590_in;
logic cond590_write_en;
logic cond590_clk;
logic cond590_reset;
logic cond590_out;
logic cond590_done;
logic cond_wire590_in;
logic cond_wire590_out;
logic cond591_in;
logic cond591_write_en;
logic cond591_clk;
logic cond591_reset;
logic cond591_out;
logic cond591_done;
logic cond_wire591_in;
logic cond_wire591_out;
logic cond592_in;
logic cond592_write_en;
logic cond592_clk;
logic cond592_reset;
logic cond592_out;
logic cond592_done;
logic cond_wire592_in;
logic cond_wire592_out;
logic cond593_in;
logic cond593_write_en;
logic cond593_clk;
logic cond593_reset;
logic cond593_out;
logic cond593_done;
logic cond_wire593_in;
logic cond_wire593_out;
logic cond594_in;
logic cond594_write_en;
logic cond594_clk;
logic cond594_reset;
logic cond594_out;
logic cond594_done;
logic cond_wire594_in;
logic cond_wire594_out;
logic cond595_in;
logic cond595_write_en;
logic cond595_clk;
logic cond595_reset;
logic cond595_out;
logic cond595_done;
logic cond_wire595_in;
logic cond_wire595_out;
logic cond596_in;
logic cond596_write_en;
logic cond596_clk;
logic cond596_reset;
logic cond596_out;
logic cond596_done;
logic cond_wire596_in;
logic cond_wire596_out;
logic cond597_in;
logic cond597_write_en;
logic cond597_clk;
logic cond597_reset;
logic cond597_out;
logic cond597_done;
logic cond_wire597_in;
logic cond_wire597_out;
logic cond598_in;
logic cond598_write_en;
logic cond598_clk;
logic cond598_reset;
logic cond598_out;
logic cond598_done;
logic cond_wire598_in;
logic cond_wire598_out;
logic cond599_in;
logic cond599_write_en;
logic cond599_clk;
logic cond599_reset;
logic cond599_out;
logic cond599_done;
logic cond_wire599_in;
logic cond_wire599_out;
logic cond600_in;
logic cond600_write_en;
logic cond600_clk;
logic cond600_reset;
logic cond600_out;
logic cond600_done;
logic cond_wire600_in;
logic cond_wire600_out;
logic cond601_in;
logic cond601_write_en;
logic cond601_clk;
logic cond601_reset;
logic cond601_out;
logic cond601_done;
logic cond_wire601_in;
logic cond_wire601_out;
logic cond602_in;
logic cond602_write_en;
logic cond602_clk;
logic cond602_reset;
logic cond602_out;
logic cond602_done;
logic cond_wire602_in;
logic cond_wire602_out;
logic cond603_in;
logic cond603_write_en;
logic cond603_clk;
logic cond603_reset;
logic cond603_out;
logic cond603_done;
logic cond_wire603_in;
logic cond_wire603_out;
logic cond604_in;
logic cond604_write_en;
logic cond604_clk;
logic cond604_reset;
logic cond604_out;
logic cond604_done;
logic cond_wire604_in;
logic cond_wire604_out;
logic cond605_in;
logic cond605_write_en;
logic cond605_clk;
logic cond605_reset;
logic cond605_out;
logic cond605_done;
logic cond_wire605_in;
logic cond_wire605_out;
logic cond606_in;
logic cond606_write_en;
logic cond606_clk;
logic cond606_reset;
logic cond606_out;
logic cond606_done;
logic cond_wire606_in;
logic cond_wire606_out;
logic cond607_in;
logic cond607_write_en;
logic cond607_clk;
logic cond607_reset;
logic cond607_out;
logic cond607_done;
logic cond_wire607_in;
logic cond_wire607_out;
logic cond608_in;
logic cond608_write_en;
logic cond608_clk;
logic cond608_reset;
logic cond608_out;
logic cond608_done;
logic cond_wire608_in;
logic cond_wire608_out;
logic cond609_in;
logic cond609_write_en;
logic cond609_clk;
logic cond609_reset;
logic cond609_out;
logic cond609_done;
logic cond_wire609_in;
logic cond_wire609_out;
logic cond610_in;
logic cond610_write_en;
logic cond610_clk;
logic cond610_reset;
logic cond610_out;
logic cond610_done;
logic cond_wire610_in;
logic cond_wire610_out;
logic cond611_in;
logic cond611_write_en;
logic cond611_clk;
logic cond611_reset;
logic cond611_out;
logic cond611_done;
logic cond_wire611_in;
logic cond_wire611_out;
logic cond612_in;
logic cond612_write_en;
logic cond612_clk;
logic cond612_reset;
logic cond612_out;
logic cond612_done;
logic cond_wire612_in;
logic cond_wire612_out;
logic cond613_in;
logic cond613_write_en;
logic cond613_clk;
logic cond613_reset;
logic cond613_out;
logic cond613_done;
logic cond_wire613_in;
logic cond_wire613_out;
logic cond614_in;
logic cond614_write_en;
logic cond614_clk;
logic cond614_reset;
logic cond614_out;
logic cond614_done;
logic cond_wire614_in;
logic cond_wire614_out;
logic cond615_in;
logic cond615_write_en;
logic cond615_clk;
logic cond615_reset;
logic cond615_out;
logic cond615_done;
logic cond_wire615_in;
logic cond_wire615_out;
logic cond616_in;
logic cond616_write_en;
logic cond616_clk;
logic cond616_reset;
logic cond616_out;
logic cond616_done;
logic cond_wire616_in;
logic cond_wire616_out;
logic cond617_in;
logic cond617_write_en;
logic cond617_clk;
logic cond617_reset;
logic cond617_out;
logic cond617_done;
logic cond_wire617_in;
logic cond_wire617_out;
logic cond618_in;
logic cond618_write_en;
logic cond618_clk;
logic cond618_reset;
logic cond618_out;
logic cond618_done;
logic cond_wire618_in;
logic cond_wire618_out;
logic cond619_in;
logic cond619_write_en;
logic cond619_clk;
logic cond619_reset;
logic cond619_out;
logic cond619_done;
logic cond_wire619_in;
logic cond_wire619_out;
logic cond620_in;
logic cond620_write_en;
logic cond620_clk;
logic cond620_reset;
logic cond620_out;
logic cond620_done;
logic cond_wire620_in;
logic cond_wire620_out;
logic cond621_in;
logic cond621_write_en;
logic cond621_clk;
logic cond621_reset;
logic cond621_out;
logic cond621_done;
logic cond_wire621_in;
logic cond_wire621_out;
logic cond622_in;
logic cond622_write_en;
logic cond622_clk;
logic cond622_reset;
logic cond622_out;
logic cond622_done;
logic cond_wire622_in;
logic cond_wire622_out;
logic cond623_in;
logic cond623_write_en;
logic cond623_clk;
logic cond623_reset;
logic cond623_out;
logic cond623_done;
logic cond_wire623_in;
logic cond_wire623_out;
logic cond624_in;
logic cond624_write_en;
logic cond624_clk;
logic cond624_reset;
logic cond624_out;
logic cond624_done;
logic cond_wire624_in;
logic cond_wire624_out;
logic cond625_in;
logic cond625_write_en;
logic cond625_clk;
logic cond625_reset;
logic cond625_out;
logic cond625_done;
logic cond_wire625_in;
logic cond_wire625_out;
logic cond626_in;
logic cond626_write_en;
logic cond626_clk;
logic cond626_reset;
logic cond626_out;
logic cond626_done;
logic cond_wire626_in;
logic cond_wire626_out;
logic cond627_in;
logic cond627_write_en;
logic cond627_clk;
logic cond627_reset;
logic cond627_out;
logic cond627_done;
logic cond_wire627_in;
logic cond_wire627_out;
logic cond628_in;
logic cond628_write_en;
logic cond628_clk;
logic cond628_reset;
logic cond628_out;
logic cond628_done;
logic cond_wire628_in;
logic cond_wire628_out;
logic cond629_in;
logic cond629_write_en;
logic cond629_clk;
logic cond629_reset;
logic cond629_out;
logic cond629_done;
logic cond_wire629_in;
logic cond_wire629_out;
logic cond630_in;
logic cond630_write_en;
logic cond630_clk;
logic cond630_reset;
logic cond630_out;
logic cond630_done;
logic cond_wire630_in;
logic cond_wire630_out;
logic cond631_in;
logic cond631_write_en;
logic cond631_clk;
logic cond631_reset;
logic cond631_out;
logic cond631_done;
logic cond_wire631_in;
logic cond_wire631_out;
logic cond632_in;
logic cond632_write_en;
logic cond632_clk;
logic cond632_reset;
logic cond632_out;
logic cond632_done;
logic cond_wire632_in;
logic cond_wire632_out;
logic cond633_in;
logic cond633_write_en;
logic cond633_clk;
logic cond633_reset;
logic cond633_out;
logic cond633_done;
logic cond_wire633_in;
logic cond_wire633_out;
logic cond634_in;
logic cond634_write_en;
logic cond634_clk;
logic cond634_reset;
logic cond634_out;
logic cond634_done;
logic cond_wire634_in;
logic cond_wire634_out;
logic cond635_in;
logic cond635_write_en;
logic cond635_clk;
logic cond635_reset;
logic cond635_out;
logic cond635_done;
logic cond_wire635_in;
logic cond_wire635_out;
logic cond636_in;
logic cond636_write_en;
logic cond636_clk;
logic cond636_reset;
logic cond636_out;
logic cond636_done;
logic cond_wire636_in;
logic cond_wire636_out;
logic cond637_in;
logic cond637_write_en;
logic cond637_clk;
logic cond637_reset;
logic cond637_out;
logic cond637_done;
logic cond_wire637_in;
logic cond_wire637_out;
logic cond638_in;
logic cond638_write_en;
logic cond638_clk;
logic cond638_reset;
logic cond638_out;
logic cond638_done;
logic cond_wire638_in;
logic cond_wire638_out;
logic cond639_in;
logic cond639_write_en;
logic cond639_clk;
logic cond639_reset;
logic cond639_out;
logic cond639_done;
logic cond_wire639_in;
logic cond_wire639_out;
logic cond640_in;
logic cond640_write_en;
logic cond640_clk;
logic cond640_reset;
logic cond640_out;
logic cond640_done;
logic cond_wire640_in;
logic cond_wire640_out;
logic cond641_in;
logic cond641_write_en;
logic cond641_clk;
logic cond641_reset;
logic cond641_out;
logic cond641_done;
logic cond_wire641_in;
logic cond_wire641_out;
logic cond642_in;
logic cond642_write_en;
logic cond642_clk;
logic cond642_reset;
logic cond642_out;
logic cond642_done;
logic cond_wire642_in;
logic cond_wire642_out;
logic cond643_in;
logic cond643_write_en;
logic cond643_clk;
logic cond643_reset;
logic cond643_out;
logic cond643_done;
logic cond_wire643_in;
logic cond_wire643_out;
logic cond644_in;
logic cond644_write_en;
logic cond644_clk;
logic cond644_reset;
logic cond644_out;
logic cond644_done;
logic cond_wire644_in;
logic cond_wire644_out;
logic cond645_in;
logic cond645_write_en;
logic cond645_clk;
logic cond645_reset;
logic cond645_out;
logic cond645_done;
logic cond_wire645_in;
logic cond_wire645_out;
logic cond646_in;
logic cond646_write_en;
logic cond646_clk;
logic cond646_reset;
logic cond646_out;
logic cond646_done;
logic cond_wire646_in;
logic cond_wire646_out;
logic cond647_in;
logic cond647_write_en;
logic cond647_clk;
logic cond647_reset;
logic cond647_out;
logic cond647_done;
logic cond_wire647_in;
logic cond_wire647_out;
logic cond648_in;
logic cond648_write_en;
logic cond648_clk;
logic cond648_reset;
logic cond648_out;
logic cond648_done;
logic cond_wire648_in;
logic cond_wire648_out;
logic cond649_in;
logic cond649_write_en;
logic cond649_clk;
logic cond649_reset;
logic cond649_out;
logic cond649_done;
logic cond_wire649_in;
logic cond_wire649_out;
logic cond650_in;
logic cond650_write_en;
logic cond650_clk;
logic cond650_reset;
logic cond650_out;
logic cond650_done;
logic cond_wire650_in;
logic cond_wire650_out;
logic cond651_in;
logic cond651_write_en;
logic cond651_clk;
logic cond651_reset;
logic cond651_out;
logic cond651_done;
logic cond_wire651_in;
logic cond_wire651_out;
logic cond652_in;
logic cond652_write_en;
logic cond652_clk;
logic cond652_reset;
logic cond652_out;
logic cond652_done;
logic cond_wire652_in;
logic cond_wire652_out;
logic cond653_in;
logic cond653_write_en;
logic cond653_clk;
logic cond653_reset;
logic cond653_out;
logic cond653_done;
logic cond_wire653_in;
logic cond_wire653_out;
logic cond654_in;
logic cond654_write_en;
logic cond654_clk;
logic cond654_reset;
logic cond654_out;
logic cond654_done;
logic cond_wire654_in;
logic cond_wire654_out;
logic cond655_in;
logic cond655_write_en;
logic cond655_clk;
logic cond655_reset;
logic cond655_out;
logic cond655_done;
logic cond_wire655_in;
logic cond_wire655_out;
logic cond656_in;
logic cond656_write_en;
logic cond656_clk;
logic cond656_reset;
logic cond656_out;
logic cond656_done;
logic cond_wire656_in;
logic cond_wire656_out;
logic cond657_in;
logic cond657_write_en;
logic cond657_clk;
logic cond657_reset;
logic cond657_out;
logic cond657_done;
logic cond_wire657_in;
logic cond_wire657_out;
logic cond658_in;
logic cond658_write_en;
logic cond658_clk;
logic cond658_reset;
logic cond658_out;
logic cond658_done;
logic cond_wire658_in;
logic cond_wire658_out;
logic cond659_in;
logic cond659_write_en;
logic cond659_clk;
logic cond659_reset;
logic cond659_out;
logic cond659_done;
logic cond_wire659_in;
logic cond_wire659_out;
logic cond660_in;
logic cond660_write_en;
logic cond660_clk;
logic cond660_reset;
logic cond660_out;
logic cond660_done;
logic cond_wire660_in;
logic cond_wire660_out;
logic cond661_in;
logic cond661_write_en;
logic cond661_clk;
logic cond661_reset;
logic cond661_out;
logic cond661_done;
logic cond_wire661_in;
logic cond_wire661_out;
logic cond662_in;
logic cond662_write_en;
logic cond662_clk;
logic cond662_reset;
logic cond662_out;
logic cond662_done;
logic cond_wire662_in;
logic cond_wire662_out;
logic cond663_in;
logic cond663_write_en;
logic cond663_clk;
logic cond663_reset;
logic cond663_out;
logic cond663_done;
logic cond_wire663_in;
logic cond_wire663_out;
logic cond664_in;
logic cond664_write_en;
logic cond664_clk;
logic cond664_reset;
logic cond664_out;
logic cond664_done;
logic cond_wire664_in;
logic cond_wire664_out;
logic cond665_in;
logic cond665_write_en;
logic cond665_clk;
logic cond665_reset;
logic cond665_out;
logic cond665_done;
logic cond_wire665_in;
logic cond_wire665_out;
logic cond666_in;
logic cond666_write_en;
logic cond666_clk;
logic cond666_reset;
logic cond666_out;
logic cond666_done;
logic cond_wire666_in;
logic cond_wire666_out;
logic cond667_in;
logic cond667_write_en;
logic cond667_clk;
logic cond667_reset;
logic cond667_out;
logic cond667_done;
logic cond_wire667_in;
logic cond_wire667_out;
logic cond668_in;
logic cond668_write_en;
logic cond668_clk;
logic cond668_reset;
logic cond668_out;
logic cond668_done;
logic cond_wire668_in;
logic cond_wire668_out;
logic cond669_in;
logic cond669_write_en;
logic cond669_clk;
logic cond669_reset;
logic cond669_out;
logic cond669_done;
logic cond_wire669_in;
logic cond_wire669_out;
logic cond670_in;
logic cond670_write_en;
logic cond670_clk;
logic cond670_reset;
logic cond670_out;
logic cond670_done;
logic cond_wire670_in;
logic cond_wire670_out;
logic cond671_in;
logic cond671_write_en;
logic cond671_clk;
logic cond671_reset;
logic cond671_out;
logic cond671_done;
logic cond_wire671_in;
logic cond_wire671_out;
logic cond672_in;
logic cond672_write_en;
logic cond672_clk;
logic cond672_reset;
logic cond672_out;
logic cond672_done;
logic cond_wire672_in;
logic cond_wire672_out;
logic cond673_in;
logic cond673_write_en;
logic cond673_clk;
logic cond673_reset;
logic cond673_out;
logic cond673_done;
logic cond_wire673_in;
logic cond_wire673_out;
logic cond674_in;
logic cond674_write_en;
logic cond674_clk;
logic cond674_reset;
logic cond674_out;
logic cond674_done;
logic cond_wire674_in;
logic cond_wire674_out;
logic cond675_in;
logic cond675_write_en;
logic cond675_clk;
logic cond675_reset;
logic cond675_out;
logic cond675_done;
logic cond_wire675_in;
logic cond_wire675_out;
logic cond676_in;
logic cond676_write_en;
logic cond676_clk;
logic cond676_reset;
logic cond676_out;
logic cond676_done;
logic cond_wire676_in;
logic cond_wire676_out;
logic cond677_in;
logic cond677_write_en;
logic cond677_clk;
logic cond677_reset;
logic cond677_out;
logic cond677_done;
logic cond_wire677_in;
logic cond_wire677_out;
logic cond678_in;
logic cond678_write_en;
logic cond678_clk;
logic cond678_reset;
logic cond678_out;
logic cond678_done;
logic cond_wire678_in;
logic cond_wire678_out;
logic cond679_in;
logic cond679_write_en;
logic cond679_clk;
logic cond679_reset;
logic cond679_out;
logic cond679_done;
logic cond_wire679_in;
logic cond_wire679_out;
logic cond680_in;
logic cond680_write_en;
logic cond680_clk;
logic cond680_reset;
logic cond680_out;
logic cond680_done;
logic cond_wire680_in;
logic cond_wire680_out;
logic cond681_in;
logic cond681_write_en;
logic cond681_clk;
logic cond681_reset;
logic cond681_out;
logic cond681_done;
logic cond_wire681_in;
logic cond_wire681_out;
logic cond682_in;
logic cond682_write_en;
logic cond682_clk;
logic cond682_reset;
logic cond682_out;
logic cond682_done;
logic cond_wire682_in;
logic cond_wire682_out;
logic cond683_in;
logic cond683_write_en;
logic cond683_clk;
logic cond683_reset;
logic cond683_out;
logic cond683_done;
logic cond_wire683_in;
logic cond_wire683_out;
logic cond684_in;
logic cond684_write_en;
logic cond684_clk;
logic cond684_reset;
logic cond684_out;
logic cond684_done;
logic cond_wire684_in;
logic cond_wire684_out;
logic cond685_in;
logic cond685_write_en;
logic cond685_clk;
logic cond685_reset;
logic cond685_out;
logic cond685_done;
logic cond_wire685_in;
logic cond_wire685_out;
logic cond686_in;
logic cond686_write_en;
logic cond686_clk;
logic cond686_reset;
logic cond686_out;
logic cond686_done;
logic cond_wire686_in;
logic cond_wire686_out;
logic cond687_in;
logic cond687_write_en;
logic cond687_clk;
logic cond687_reset;
logic cond687_out;
logic cond687_done;
logic cond_wire687_in;
logic cond_wire687_out;
logic cond688_in;
logic cond688_write_en;
logic cond688_clk;
logic cond688_reset;
logic cond688_out;
logic cond688_done;
logic cond_wire688_in;
logic cond_wire688_out;
logic cond689_in;
logic cond689_write_en;
logic cond689_clk;
logic cond689_reset;
logic cond689_out;
logic cond689_done;
logic cond_wire689_in;
logic cond_wire689_out;
logic cond690_in;
logic cond690_write_en;
logic cond690_clk;
logic cond690_reset;
logic cond690_out;
logic cond690_done;
logic cond_wire690_in;
logic cond_wire690_out;
logic cond691_in;
logic cond691_write_en;
logic cond691_clk;
logic cond691_reset;
logic cond691_out;
logic cond691_done;
logic cond_wire691_in;
logic cond_wire691_out;
logic cond692_in;
logic cond692_write_en;
logic cond692_clk;
logic cond692_reset;
logic cond692_out;
logic cond692_done;
logic cond_wire692_in;
logic cond_wire692_out;
logic cond693_in;
logic cond693_write_en;
logic cond693_clk;
logic cond693_reset;
logic cond693_out;
logic cond693_done;
logic cond_wire693_in;
logic cond_wire693_out;
logic cond694_in;
logic cond694_write_en;
logic cond694_clk;
logic cond694_reset;
logic cond694_out;
logic cond694_done;
logic cond_wire694_in;
logic cond_wire694_out;
logic cond695_in;
logic cond695_write_en;
logic cond695_clk;
logic cond695_reset;
logic cond695_out;
logic cond695_done;
logic cond_wire695_in;
logic cond_wire695_out;
logic cond696_in;
logic cond696_write_en;
logic cond696_clk;
logic cond696_reset;
logic cond696_out;
logic cond696_done;
logic cond_wire696_in;
logic cond_wire696_out;
logic cond697_in;
logic cond697_write_en;
logic cond697_clk;
logic cond697_reset;
logic cond697_out;
logic cond697_done;
logic cond_wire697_in;
logic cond_wire697_out;
logic cond698_in;
logic cond698_write_en;
logic cond698_clk;
logic cond698_reset;
logic cond698_out;
logic cond698_done;
logic cond_wire698_in;
logic cond_wire698_out;
logic cond699_in;
logic cond699_write_en;
logic cond699_clk;
logic cond699_reset;
logic cond699_out;
logic cond699_done;
logic cond_wire699_in;
logic cond_wire699_out;
logic cond700_in;
logic cond700_write_en;
logic cond700_clk;
logic cond700_reset;
logic cond700_out;
logic cond700_done;
logic cond_wire700_in;
logic cond_wire700_out;
logic cond701_in;
logic cond701_write_en;
logic cond701_clk;
logic cond701_reset;
logic cond701_out;
logic cond701_done;
logic cond_wire701_in;
logic cond_wire701_out;
logic cond702_in;
logic cond702_write_en;
logic cond702_clk;
logic cond702_reset;
logic cond702_out;
logic cond702_done;
logic cond_wire702_in;
logic cond_wire702_out;
logic cond703_in;
logic cond703_write_en;
logic cond703_clk;
logic cond703_reset;
logic cond703_out;
logic cond703_done;
logic cond_wire703_in;
logic cond_wire703_out;
logic cond704_in;
logic cond704_write_en;
logic cond704_clk;
logic cond704_reset;
logic cond704_out;
logic cond704_done;
logic cond_wire704_in;
logic cond_wire704_out;
logic cond705_in;
logic cond705_write_en;
logic cond705_clk;
logic cond705_reset;
logic cond705_out;
logic cond705_done;
logic cond_wire705_in;
logic cond_wire705_out;
logic cond706_in;
logic cond706_write_en;
logic cond706_clk;
logic cond706_reset;
logic cond706_out;
logic cond706_done;
logic cond_wire706_in;
logic cond_wire706_out;
logic cond707_in;
logic cond707_write_en;
logic cond707_clk;
logic cond707_reset;
logic cond707_out;
logic cond707_done;
logic cond_wire707_in;
logic cond_wire707_out;
logic cond708_in;
logic cond708_write_en;
logic cond708_clk;
logic cond708_reset;
logic cond708_out;
logic cond708_done;
logic cond_wire708_in;
logic cond_wire708_out;
logic cond709_in;
logic cond709_write_en;
logic cond709_clk;
logic cond709_reset;
logic cond709_out;
logic cond709_done;
logic cond_wire709_in;
logic cond_wire709_out;
logic cond710_in;
logic cond710_write_en;
logic cond710_clk;
logic cond710_reset;
logic cond710_out;
logic cond710_done;
logic cond_wire710_in;
logic cond_wire710_out;
logic cond711_in;
logic cond711_write_en;
logic cond711_clk;
logic cond711_reset;
logic cond711_out;
logic cond711_done;
logic cond_wire711_in;
logic cond_wire711_out;
logic cond712_in;
logic cond712_write_en;
logic cond712_clk;
logic cond712_reset;
logic cond712_out;
logic cond712_done;
logic cond_wire712_in;
logic cond_wire712_out;
logic cond713_in;
logic cond713_write_en;
logic cond713_clk;
logic cond713_reset;
logic cond713_out;
logic cond713_done;
logic cond_wire713_in;
logic cond_wire713_out;
logic cond714_in;
logic cond714_write_en;
logic cond714_clk;
logic cond714_reset;
logic cond714_out;
logic cond714_done;
logic cond_wire714_in;
logic cond_wire714_out;
logic cond715_in;
logic cond715_write_en;
logic cond715_clk;
logic cond715_reset;
logic cond715_out;
logic cond715_done;
logic cond_wire715_in;
logic cond_wire715_out;
logic cond716_in;
logic cond716_write_en;
logic cond716_clk;
logic cond716_reset;
logic cond716_out;
logic cond716_done;
logic cond_wire716_in;
logic cond_wire716_out;
logic cond717_in;
logic cond717_write_en;
logic cond717_clk;
logic cond717_reset;
logic cond717_out;
logic cond717_done;
logic cond_wire717_in;
logic cond_wire717_out;
logic cond718_in;
logic cond718_write_en;
logic cond718_clk;
logic cond718_reset;
logic cond718_out;
logic cond718_done;
logic cond_wire718_in;
logic cond_wire718_out;
logic cond719_in;
logic cond719_write_en;
logic cond719_clk;
logic cond719_reset;
logic cond719_out;
logic cond719_done;
logic cond_wire719_in;
logic cond_wire719_out;
logic cond720_in;
logic cond720_write_en;
logic cond720_clk;
logic cond720_reset;
logic cond720_out;
logic cond720_done;
logic cond_wire720_in;
logic cond_wire720_out;
logic cond721_in;
logic cond721_write_en;
logic cond721_clk;
logic cond721_reset;
logic cond721_out;
logic cond721_done;
logic cond_wire721_in;
logic cond_wire721_out;
logic cond722_in;
logic cond722_write_en;
logic cond722_clk;
logic cond722_reset;
logic cond722_out;
logic cond722_done;
logic cond_wire722_in;
logic cond_wire722_out;
logic cond723_in;
logic cond723_write_en;
logic cond723_clk;
logic cond723_reset;
logic cond723_out;
logic cond723_done;
logic cond_wire723_in;
logic cond_wire723_out;
logic cond724_in;
logic cond724_write_en;
logic cond724_clk;
logic cond724_reset;
logic cond724_out;
logic cond724_done;
logic cond_wire724_in;
logic cond_wire724_out;
logic cond725_in;
logic cond725_write_en;
logic cond725_clk;
logic cond725_reset;
logic cond725_out;
logic cond725_done;
logic cond_wire725_in;
logic cond_wire725_out;
logic cond726_in;
logic cond726_write_en;
logic cond726_clk;
logic cond726_reset;
logic cond726_out;
logic cond726_done;
logic cond_wire726_in;
logic cond_wire726_out;
logic cond727_in;
logic cond727_write_en;
logic cond727_clk;
logic cond727_reset;
logic cond727_out;
logic cond727_done;
logic cond_wire727_in;
logic cond_wire727_out;
logic cond728_in;
logic cond728_write_en;
logic cond728_clk;
logic cond728_reset;
logic cond728_out;
logic cond728_done;
logic cond_wire728_in;
logic cond_wire728_out;
logic cond729_in;
logic cond729_write_en;
logic cond729_clk;
logic cond729_reset;
logic cond729_out;
logic cond729_done;
logic cond_wire729_in;
logic cond_wire729_out;
logic cond730_in;
logic cond730_write_en;
logic cond730_clk;
logic cond730_reset;
logic cond730_out;
logic cond730_done;
logic cond_wire730_in;
logic cond_wire730_out;
logic cond731_in;
logic cond731_write_en;
logic cond731_clk;
logic cond731_reset;
logic cond731_out;
logic cond731_done;
logic cond_wire731_in;
logic cond_wire731_out;
logic cond732_in;
logic cond732_write_en;
logic cond732_clk;
logic cond732_reset;
logic cond732_out;
logic cond732_done;
logic cond_wire732_in;
logic cond_wire732_out;
logic cond733_in;
logic cond733_write_en;
logic cond733_clk;
logic cond733_reset;
logic cond733_out;
logic cond733_done;
logic cond_wire733_in;
logic cond_wire733_out;
logic cond734_in;
logic cond734_write_en;
logic cond734_clk;
logic cond734_reset;
logic cond734_out;
logic cond734_done;
logic cond_wire734_in;
logic cond_wire734_out;
logic cond735_in;
logic cond735_write_en;
logic cond735_clk;
logic cond735_reset;
logic cond735_out;
logic cond735_done;
logic cond_wire735_in;
logic cond_wire735_out;
logic cond736_in;
logic cond736_write_en;
logic cond736_clk;
logic cond736_reset;
logic cond736_out;
logic cond736_done;
logic cond_wire736_in;
logic cond_wire736_out;
logic cond737_in;
logic cond737_write_en;
logic cond737_clk;
logic cond737_reset;
logic cond737_out;
logic cond737_done;
logic cond_wire737_in;
logic cond_wire737_out;
logic cond738_in;
logic cond738_write_en;
logic cond738_clk;
logic cond738_reset;
logic cond738_out;
logic cond738_done;
logic cond_wire738_in;
logic cond_wire738_out;
logic cond739_in;
logic cond739_write_en;
logic cond739_clk;
logic cond739_reset;
logic cond739_out;
logic cond739_done;
logic cond_wire739_in;
logic cond_wire739_out;
logic cond740_in;
logic cond740_write_en;
logic cond740_clk;
logic cond740_reset;
logic cond740_out;
logic cond740_done;
logic cond_wire740_in;
logic cond_wire740_out;
logic cond741_in;
logic cond741_write_en;
logic cond741_clk;
logic cond741_reset;
logic cond741_out;
logic cond741_done;
logic cond_wire741_in;
logic cond_wire741_out;
logic cond742_in;
logic cond742_write_en;
logic cond742_clk;
logic cond742_reset;
logic cond742_out;
logic cond742_done;
logic cond_wire742_in;
logic cond_wire742_out;
logic cond743_in;
logic cond743_write_en;
logic cond743_clk;
logic cond743_reset;
logic cond743_out;
logic cond743_done;
logic cond_wire743_in;
logic cond_wire743_out;
logic cond744_in;
logic cond744_write_en;
logic cond744_clk;
logic cond744_reset;
logic cond744_out;
logic cond744_done;
logic cond_wire744_in;
logic cond_wire744_out;
logic cond745_in;
logic cond745_write_en;
logic cond745_clk;
logic cond745_reset;
logic cond745_out;
logic cond745_done;
logic cond_wire745_in;
logic cond_wire745_out;
logic cond746_in;
logic cond746_write_en;
logic cond746_clk;
logic cond746_reset;
logic cond746_out;
logic cond746_done;
logic cond_wire746_in;
logic cond_wire746_out;
logic cond747_in;
logic cond747_write_en;
logic cond747_clk;
logic cond747_reset;
logic cond747_out;
logic cond747_done;
logic cond_wire747_in;
logic cond_wire747_out;
logic cond748_in;
logic cond748_write_en;
logic cond748_clk;
logic cond748_reset;
logic cond748_out;
logic cond748_done;
logic cond_wire748_in;
logic cond_wire748_out;
logic cond749_in;
logic cond749_write_en;
logic cond749_clk;
logic cond749_reset;
logic cond749_out;
logic cond749_done;
logic cond_wire749_in;
logic cond_wire749_out;
logic cond750_in;
logic cond750_write_en;
logic cond750_clk;
logic cond750_reset;
logic cond750_out;
logic cond750_done;
logic cond_wire750_in;
logic cond_wire750_out;
logic cond751_in;
logic cond751_write_en;
logic cond751_clk;
logic cond751_reset;
logic cond751_out;
logic cond751_done;
logic cond_wire751_in;
logic cond_wire751_out;
logic cond752_in;
logic cond752_write_en;
logic cond752_clk;
logic cond752_reset;
logic cond752_out;
logic cond752_done;
logic cond_wire752_in;
logic cond_wire752_out;
logic cond753_in;
logic cond753_write_en;
logic cond753_clk;
logic cond753_reset;
logic cond753_out;
logic cond753_done;
logic cond_wire753_in;
logic cond_wire753_out;
logic cond754_in;
logic cond754_write_en;
logic cond754_clk;
logic cond754_reset;
logic cond754_out;
logic cond754_done;
logic cond_wire754_in;
logic cond_wire754_out;
logic cond755_in;
logic cond755_write_en;
logic cond755_clk;
logic cond755_reset;
logic cond755_out;
logic cond755_done;
logic cond_wire755_in;
logic cond_wire755_out;
logic cond756_in;
logic cond756_write_en;
logic cond756_clk;
logic cond756_reset;
logic cond756_out;
logic cond756_done;
logic cond_wire756_in;
logic cond_wire756_out;
logic cond757_in;
logic cond757_write_en;
logic cond757_clk;
logic cond757_reset;
logic cond757_out;
logic cond757_done;
logic cond_wire757_in;
logic cond_wire757_out;
logic cond758_in;
logic cond758_write_en;
logic cond758_clk;
logic cond758_reset;
logic cond758_out;
logic cond758_done;
logic cond_wire758_in;
logic cond_wire758_out;
logic cond759_in;
logic cond759_write_en;
logic cond759_clk;
logic cond759_reset;
logic cond759_out;
logic cond759_done;
logic cond_wire759_in;
logic cond_wire759_out;
logic cond760_in;
logic cond760_write_en;
logic cond760_clk;
logic cond760_reset;
logic cond760_out;
logic cond760_done;
logic cond_wire760_in;
logic cond_wire760_out;
logic cond761_in;
logic cond761_write_en;
logic cond761_clk;
logic cond761_reset;
logic cond761_out;
logic cond761_done;
logic cond_wire761_in;
logic cond_wire761_out;
logic cond762_in;
logic cond762_write_en;
logic cond762_clk;
logic cond762_reset;
logic cond762_out;
logic cond762_done;
logic cond_wire762_in;
logic cond_wire762_out;
logic cond763_in;
logic cond763_write_en;
logic cond763_clk;
logic cond763_reset;
logic cond763_out;
logic cond763_done;
logic cond_wire763_in;
logic cond_wire763_out;
logic cond764_in;
logic cond764_write_en;
logic cond764_clk;
logic cond764_reset;
logic cond764_out;
logic cond764_done;
logic cond_wire764_in;
logic cond_wire764_out;
logic cond765_in;
logic cond765_write_en;
logic cond765_clk;
logic cond765_reset;
logic cond765_out;
logic cond765_done;
logic cond_wire765_in;
logic cond_wire765_out;
logic cond766_in;
logic cond766_write_en;
logic cond766_clk;
logic cond766_reset;
logic cond766_out;
logic cond766_done;
logic cond_wire766_in;
logic cond_wire766_out;
logic cond767_in;
logic cond767_write_en;
logic cond767_clk;
logic cond767_reset;
logic cond767_out;
logic cond767_done;
logic cond_wire767_in;
logic cond_wire767_out;
logic cond768_in;
logic cond768_write_en;
logic cond768_clk;
logic cond768_reset;
logic cond768_out;
logic cond768_done;
logic cond_wire768_in;
logic cond_wire768_out;
logic cond769_in;
logic cond769_write_en;
logic cond769_clk;
logic cond769_reset;
logic cond769_out;
logic cond769_done;
logic cond_wire769_in;
logic cond_wire769_out;
logic cond770_in;
logic cond770_write_en;
logic cond770_clk;
logic cond770_reset;
logic cond770_out;
logic cond770_done;
logic cond_wire770_in;
logic cond_wire770_out;
logic cond771_in;
logic cond771_write_en;
logic cond771_clk;
logic cond771_reset;
logic cond771_out;
logic cond771_done;
logic cond_wire771_in;
logic cond_wire771_out;
logic cond772_in;
logic cond772_write_en;
logic cond772_clk;
logic cond772_reset;
logic cond772_out;
logic cond772_done;
logic cond_wire772_in;
logic cond_wire772_out;
logic cond773_in;
logic cond773_write_en;
logic cond773_clk;
logic cond773_reset;
logic cond773_out;
logic cond773_done;
logic cond_wire773_in;
logic cond_wire773_out;
logic cond774_in;
logic cond774_write_en;
logic cond774_clk;
logic cond774_reset;
logic cond774_out;
logic cond774_done;
logic cond_wire774_in;
logic cond_wire774_out;
logic cond775_in;
logic cond775_write_en;
logic cond775_clk;
logic cond775_reset;
logic cond775_out;
logic cond775_done;
logic cond_wire775_in;
logic cond_wire775_out;
logic cond776_in;
logic cond776_write_en;
logic cond776_clk;
logic cond776_reset;
logic cond776_out;
logic cond776_done;
logic cond_wire776_in;
logic cond_wire776_out;
logic cond777_in;
logic cond777_write_en;
logic cond777_clk;
logic cond777_reset;
logic cond777_out;
logic cond777_done;
logic cond_wire777_in;
logic cond_wire777_out;
logic cond778_in;
logic cond778_write_en;
logic cond778_clk;
logic cond778_reset;
logic cond778_out;
logic cond778_done;
logic cond_wire778_in;
logic cond_wire778_out;
logic cond779_in;
logic cond779_write_en;
logic cond779_clk;
logic cond779_reset;
logic cond779_out;
logic cond779_done;
logic cond_wire779_in;
logic cond_wire779_out;
logic cond780_in;
logic cond780_write_en;
logic cond780_clk;
logic cond780_reset;
logic cond780_out;
logic cond780_done;
logic cond_wire780_in;
logic cond_wire780_out;
logic cond781_in;
logic cond781_write_en;
logic cond781_clk;
logic cond781_reset;
logic cond781_out;
logic cond781_done;
logic cond_wire781_in;
logic cond_wire781_out;
logic cond782_in;
logic cond782_write_en;
logic cond782_clk;
logic cond782_reset;
logic cond782_out;
logic cond782_done;
logic cond_wire782_in;
logic cond_wire782_out;
logic cond783_in;
logic cond783_write_en;
logic cond783_clk;
logic cond783_reset;
logic cond783_out;
logic cond783_done;
logic cond_wire783_in;
logic cond_wire783_out;
logic cond784_in;
logic cond784_write_en;
logic cond784_clk;
logic cond784_reset;
logic cond784_out;
logic cond784_done;
logic cond_wire784_in;
logic cond_wire784_out;
logic cond785_in;
logic cond785_write_en;
logic cond785_clk;
logic cond785_reset;
logic cond785_out;
logic cond785_done;
logic cond_wire785_in;
logic cond_wire785_out;
logic cond786_in;
logic cond786_write_en;
logic cond786_clk;
logic cond786_reset;
logic cond786_out;
logic cond786_done;
logic cond_wire786_in;
logic cond_wire786_out;
logic cond787_in;
logic cond787_write_en;
logic cond787_clk;
logic cond787_reset;
logic cond787_out;
logic cond787_done;
logic cond_wire787_in;
logic cond_wire787_out;
logic cond788_in;
logic cond788_write_en;
logic cond788_clk;
logic cond788_reset;
logic cond788_out;
logic cond788_done;
logic cond_wire788_in;
logic cond_wire788_out;
logic cond789_in;
logic cond789_write_en;
logic cond789_clk;
logic cond789_reset;
logic cond789_out;
logic cond789_done;
logic cond_wire789_in;
logic cond_wire789_out;
logic cond790_in;
logic cond790_write_en;
logic cond790_clk;
logic cond790_reset;
logic cond790_out;
logic cond790_done;
logic cond_wire790_in;
logic cond_wire790_out;
logic cond791_in;
logic cond791_write_en;
logic cond791_clk;
logic cond791_reset;
logic cond791_out;
logic cond791_done;
logic cond_wire791_in;
logic cond_wire791_out;
logic cond792_in;
logic cond792_write_en;
logic cond792_clk;
logic cond792_reset;
logic cond792_out;
logic cond792_done;
logic cond_wire792_in;
logic cond_wire792_out;
logic cond793_in;
logic cond793_write_en;
logic cond793_clk;
logic cond793_reset;
logic cond793_out;
logic cond793_done;
logic cond_wire793_in;
logic cond_wire793_out;
logic cond794_in;
logic cond794_write_en;
logic cond794_clk;
logic cond794_reset;
logic cond794_out;
logic cond794_done;
logic cond_wire794_in;
logic cond_wire794_out;
logic cond795_in;
logic cond795_write_en;
logic cond795_clk;
logic cond795_reset;
logic cond795_out;
logic cond795_done;
logic cond_wire795_in;
logic cond_wire795_out;
logic cond796_in;
logic cond796_write_en;
logic cond796_clk;
logic cond796_reset;
logic cond796_out;
logic cond796_done;
logic cond_wire796_in;
logic cond_wire796_out;
logic cond797_in;
logic cond797_write_en;
logic cond797_clk;
logic cond797_reset;
logic cond797_out;
logic cond797_done;
logic cond_wire797_in;
logic cond_wire797_out;
logic cond798_in;
logic cond798_write_en;
logic cond798_clk;
logic cond798_reset;
logic cond798_out;
logic cond798_done;
logic cond_wire798_in;
logic cond_wire798_out;
logic cond799_in;
logic cond799_write_en;
logic cond799_clk;
logic cond799_reset;
logic cond799_out;
logic cond799_done;
logic cond_wire799_in;
logic cond_wire799_out;
logic cond800_in;
logic cond800_write_en;
logic cond800_clk;
logic cond800_reset;
logic cond800_out;
logic cond800_done;
logic cond_wire800_in;
logic cond_wire800_out;
logic cond801_in;
logic cond801_write_en;
logic cond801_clk;
logic cond801_reset;
logic cond801_out;
logic cond801_done;
logic cond_wire801_in;
logic cond_wire801_out;
logic cond802_in;
logic cond802_write_en;
logic cond802_clk;
logic cond802_reset;
logic cond802_out;
logic cond802_done;
logic cond_wire802_in;
logic cond_wire802_out;
logic cond803_in;
logic cond803_write_en;
logic cond803_clk;
logic cond803_reset;
logic cond803_out;
logic cond803_done;
logic cond_wire803_in;
logic cond_wire803_out;
logic cond804_in;
logic cond804_write_en;
logic cond804_clk;
logic cond804_reset;
logic cond804_out;
logic cond804_done;
logic cond_wire804_in;
logic cond_wire804_out;
logic cond805_in;
logic cond805_write_en;
logic cond805_clk;
logic cond805_reset;
logic cond805_out;
logic cond805_done;
logic cond_wire805_in;
logic cond_wire805_out;
logic cond806_in;
logic cond806_write_en;
logic cond806_clk;
logic cond806_reset;
logic cond806_out;
logic cond806_done;
logic cond_wire806_in;
logic cond_wire806_out;
logic cond807_in;
logic cond807_write_en;
logic cond807_clk;
logic cond807_reset;
logic cond807_out;
logic cond807_done;
logic cond_wire807_in;
logic cond_wire807_out;
logic cond808_in;
logic cond808_write_en;
logic cond808_clk;
logic cond808_reset;
logic cond808_out;
logic cond808_done;
logic cond_wire808_in;
logic cond_wire808_out;
logic cond809_in;
logic cond809_write_en;
logic cond809_clk;
logic cond809_reset;
logic cond809_out;
logic cond809_done;
logic cond_wire809_in;
logic cond_wire809_out;
logic cond810_in;
logic cond810_write_en;
logic cond810_clk;
logic cond810_reset;
logic cond810_out;
logic cond810_done;
logic cond_wire810_in;
logic cond_wire810_out;
logic cond811_in;
logic cond811_write_en;
logic cond811_clk;
logic cond811_reset;
logic cond811_out;
logic cond811_done;
logic cond_wire811_in;
logic cond_wire811_out;
logic cond812_in;
logic cond812_write_en;
logic cond812_clk;
logic cond812_reset;
logic cond812_out;
logic cond812_done;
logic cond_wire812_in;
logic cond_wire812_out;
logic cond813_in;
logic cond813_write_en;
logic cond813_clk;
logic cond813_reset;
logic cond813_out;
logic cond813_done;
logic cond_wire813_in;
logic cond_wire813_out;
logic cond814_in;
logic cond814_write_en;
logic cond814_clk;
logic cond814_reset;
logic cond814_out;
logic cond814_done;
logic cond_wire814_in;
logic cond_wire814_out;
logic cond815_in;
logic cond815_write_en;
logic cond815_clk;
logic cond815_reset;
logic cond815_out;
logic cond815_done;
logic cond_wire815_in;
logic cond_wire815_out;
logic cond816_in;
logic cond816_write_en;
logic cond816_clk;
logic cond816_reset;
logic cond816_out;
logic cond816_done;
logic cond_wire816_in;
logic cond_wire816_out;
logic cond817_in;
logic cond817_write_en;
logic cond817_clk;
logic cond817_reset;
logic cond817_out;
logic cond817_done;
logic cond_wire817_in;
logic cond_wire817_out;
logic cond818_in;
logic cond818_write_en;
logic cond818_clk;
logic cond818_reset;
logic cond818_out;
logic cond818_done;
logic cond_wire818_in;
logic cond_wire818_out;
logic cond819_in;
logic cond819_write_en;
logic cond819_clk;
logic cond819_reset;
logic cond819_out;
logic cond819_done;
logic cond_wire819_in;
logic cond_wire819_out;
logic cond820_in;
logic cond820_write_en;
logic cond820_clk;
logic cond820_reset;
logic cond820_out;
logic cond820_done;
logic cond_wire820_in;
logic cond_wire820_out;
logic cond821_in;
logic cond821_write_en;
logic cond821_clk;
logic cond821_reset;
logic cond821_out;
logic cond821_done;
logic cond_wire821_in;
logic cond_wire821_out;
logic cond822_in;
logic cond822_write_en;
logic cond822_clk;
logic cond822_reset;
logic cond822_out;
logic cond822_done;
logic cond_wire822_in;
logic cond_wire822_out;
logic cond823_in;
logic cond823_write_en;
logic cond823_clk;
logic cond823_reset;
logic cond823_out;
logic cond823_done;
logic cond_wire823_in;
logic cond_wire823_out;
logic cond824_in;
logic cond824_write_en;
logic cond824_clk;
logic cond824_reset;
logic cond824_out;
logic cond824_done;
logic cond_wire824_in;
logic cond_wire824_out;
logic cond825_in;
logic cond825_write_en;
logic cond825_clk;
logic cond825_reset;
logic cond825_out;
logic cond825_done;
logic cond_wire825_in;
logic cond_wire825_out;
logic cond826_in;
logic cond826_write_en;
logic cond826_clk;
logic cond826_reset;
logic cond826_out;
logic cond826_done;
logic cond_wire826_in;
logic cond_wire826_out;
logic cond827_in;
logic cond827_write_en;
logic cond827_clk;
logic cond827_reset;
logic cond827_out;
logic cond827_done;
logic cond_wire827_in;
logic cond_wire827_out;
logic cond828_in;
logic cond828_write_en;
logic cond828_clk;
logic cond828_reset;
logic cond828_out;
logic cond828_done;
logic cond_wire828_in;
logic cond_wire828_out;
logic cond829_in;
logic cond829_write_en;
logic cond829_clk;
logic cond829_reset;
logic cond829_out;
logic cond829_done;
logic cond_wire829_in;
logic cond_wire829_out;
logic cond830_in;
logic cond830_write_en;
logic cond830_clk;
logic cond830_reset;
logic cond830_out;
logic cond830_done;
logic cond_wire830_in;
logic cond_wire830_out;
logic cond831_in;
logic cond831_write_en;
logic cond831_clk;
logic cond831_reset;
logic cond831_out;
logic cond831_done;
logic cond_wire831_in;
logic cond_wire831_out;
logic cond832_in;
logic cond832_write_en;
logic cond832_clk;
logic cond832_reset;
logic cond832_out;
logic cond832_done;
logic cond_wire832_in;
logic cond_wire832_out;
logic cond833_in;
logic cond833_write_en;
logic cond833_clk;
logic cond833_reset;
logic cond833_out;
logic cond833_done;
logic cond_wire833_in;
logic cond_wire833_out;
logic cond834_in;
logic cond834_write_en;
logic cond834_clk;
logic cond834_reset;
logic cond834_out;
logic cond834_done;
logic cond_wire834_in;
logic cond_wire834_out;
logic cond835_in;
logic cond835_write_en;
logic cond835_clk;
logic cond835_reset;
logic cond835_out;
logic cond835_done;
logic cond_wire835_in;
logic cond_wire835_out;
logic cond836_in;
logic cond836_write_en;
logic cond836_clk;
logic cond836_reset;
logic cond836_out;
logic cond836_done;
logic cond_wire836_in;
logic cond_wire836_out;
logic cond837_in;
logic cond837_write_en;
logic cond837_clk;
logic cond837_reset;
logic cond837_out;
logic cond837_done;
logic cond_wire837_in;
logic cond_wire837_out;
logic cond838_in;
logic cond838_write_en;
logic cond838_clk;
logic cond838_reset;
logic cond838_out;
logic cond838_done;
logic cond_wire838_in;
logic cond_wire838_out;
logic cond839_in;
logic cond839_write_en;
logic cond839_clk;
logic cond839_reset;
logic cond839_out;
logic cond839_done;
logic cond_wire839_in;
logic cond_wire839_out;
logic cond840_in;
logic cond840_write_en;
logic cond840_clk;
logic cond840_reset;
logic cond840_out;
logic cond840_done;
logic cond_wire840_in;
logic cond_wire840_out;
logic cond841_in;
logic cond841_write_en;
logic cond841_clk;
logic cond841_reset;
logic cond841_out;
logic cond841_done;
logic cond_wire841_in;
logic cond_wire841_out;
logic cond842_in;
logic cond842_write_en;
logic cond842_clk;
logic cond842_reset;
logic cond842_out;
logic cond842_done;
logic cond_wire842_in;
logic cond_wire842_out;
logic cond843_in;
logic cond843_write_en;
logic cond843_clk;
logic cond843_reset;
logic cond843_out;
logic cond843_done;
logic cond_wire843_in;
logic cond_wire843_out;
logic cond844_in;
logic cond844_write_en;
logic cond844_clk;
logic cond844_reset;
logic cond844_out;
logic cond844_done;
logic cond_wire844_in;
logic cond_wire844_out;
logic cond845_in;
logic cond845_write_en;
logic cond845_clk;
logic cond845_reset;
logic cond845_out;
logic cond845_done;
logic cond_wire845_in;
logic cond_wire845_out;
logic cond846_in;
logic cond846_write_en;
logic cond846_clk;
logic cond846_reset;
logic cond846_out;
logic cond846_done;
logic cond_wire846_in;
logic cond_wire846_out;
logic cond847_in;
logic cond847_write_en;
logic cond847_clk;
logic cond847_reset;
logic cond847_out;
logic cond847_done;
logic cond_wire847_in;
logic cond_wire847_out;
logic cond848_in;
logic cond848_write_en;
logic cond848_clk;
logic cond848_reset;
logic cond848_out;
logic cond848_done;
logic cond_wire848_in;
logic cond_wire848_out;
logic cond849_in;
logic cond849_write_en;
logic cond849_clk;
logic cond849_reset;
logic cond849_out;
logic cond849_done;
logic cond_wire849_in;
logic cond_wire849_out;
logic cond850_in;
logic cond850_write_en;
logic cond850_clk;
logic cond850_reset;
logic cond850_out;
logic cond850_done;
logic cond_wire850_in;
logic cond_wire850_out;
logic cond851_in;
logic cond851_write_en;
logic cond851_clk;
logic cond851_reset;
logic cond851_out;
logic cond851_done;
logic cond_wire851_in;
logic cond_wire851_out;
logic cond852_in;
logic cond852_write_en;
logic cond852_clk;
logic cond852_reset;
logic cond852_out;
logic cond852_done;
logic cond_wire852_in;
logic cond_wire852_out;
logic cond853_in;
logic cond853_write_en;
logic cond853_clk;
logic cond853_reset;
logic cond853_out;
logic cond853_done;
logic cond_wire853_in;
logic cond_wire853_out;
logic cond854_in;
logic cond854_write_en;
logic cond854_clk;
logic cond854_reset;
logic cond854_out;
logic cond854_done;
logic cond_wire854_in;
logic cond_wire854_out;
logic cond855_in;
logic cond855_write_en;
logic cond855_clk;
logic cond855_reset;
logic cond855_out;
logic cond855_done;
logic cond_wire855_in;
logic cond_wire855_out;
logic cond856_in;
logic cond856_write_en;
logic cond856_clk;
logic cond856_reset;
logic cond856_out;
logic cond856_done;
logic cond_wire856_in;
logic cond_wire856_out;
logic cond857_in;
logic cond857_write_en;
logic cond857_clk;
logic cond857_reset;
logic cond857_out;
logic cond857_done;
logic cond_wire857_in;
logic cond_wire857_out;
logic cond858_in;
logic cond858_write_en;
logic cond858_clk;
logic cond858_reset;
logic cond858_out;
logic cond858_done;
logic cond_wire858_in;
logic cond_wire858_out;
logic cond859_in;
logic cond859_write_en;
logic cond859_clk;
logic cond859_reset;
logic cond859_out;
logic cond859_done;
logic cond_wire859_in;
logic cond_wire859_out;
logic cond860_in;
logic cond860_write_en;
logic cond860_clk;
logic cond860_reset;
logic cond860_out;
logic cond860_done;
logic cond_wire860_in;
logic cond_wire860_out;
logic cond861_in;
logic cond861_write_en;
logic cond861_clk;
logic cond861_reset;
logic cond861_out;
logic cond861_done;
logic cond_wire861_in;
logic cond_wire861_out;
logic cond862_in;
logic cond862_write_en;
logic cond862_clk;
logic cond862_reset;
logic cond862_out;
logic cond862_done;
logic cond_wire862_in;
logic cond_wire862_out;
logic cond863_in;
logic cond863_write_en;
logic cond863_clk;
logic cond863_reset;
logic cond863_out;
logic cond863_done;
logic cond_wire863_in;
logic cond_wire863_out;
logic cond864_in;
logic cond864_write_en;
logic cond864_clk;
logic cond864_reset;
logic cond864_out;
logic cond864_done;
logic cond_wire864_in;
logic cond_wire864_out;
logic cond865_in;
logic cond865_write_en;
logic cond865_clk;
logic cond865_reset;
logic cond865_out;
logic cond865_done;
logic cond_wire865_in;
logic cond_wire865_out;
logic cond866_in;
logic cond866_write_en;
logic cond866_clk;
logic cond866_reset;
logic cond866_out;
logic cond866_done;
logic cond_wire866_in;
logic cond_wire866_out;
logic cond867_in;
logic cond867_write_en;
logic cond867_clk;
logic cond867_reset;
logic cond867_out;
logic cond867_done;
logic cond_wire867_in;
logic cond_wire867_out;
logic cond868_in;
logic cond868_write_en;
logic cond868_clk;
logic cond868_reset;
logic cond868_out;
logic cond868_done;
logic cond_wire868_in;
logic cond_wire868_out;
logic cond869_in;
logic cond869_write_en;
logic cond869_clk;
logic cond869_reset;
logic cond869_out;
logic cond869_done;
logic cond_wire869_in;
logic cond_wire869_out;
logic cond870_in;
logic cond870_write_en;
logic cond870_clk;
logic cond870_reset;
logic cond870_out;
logic cond870_done;
logic cond_wire870_in;
logic cond_wire870_out;
logic cond871_in;
logic cond871_write_en;
logic cond871_clk;
logic cond871_reset;
logic cond871_out;
logic cond871_done;
logic cond_wire871_in;
logic cond_wire871_out;
logic cond872_in;
logic cond872_write_en;
logic cond872_clk;
logic cond872_reset;
logic cond872_out;
logic cond872_done;
logic cond_wire872_in;
logic cond_wire872_out;
logic cond873_in;
logic cond873_write_en;
logic cond873_clk;
logic cond873_reset;
logic cond873_out;
logic cond873_done;
logic cond_wire873_in;
logic cond_wire873_out;
logic cond874_in;
logic cond874_write_en;
logic cond874_clk;
logic cond874_reset;
logic cond874_out;
logic cond874_done;
logic cond_wire874_in;
logic cond_wire874_out;
logic cond875_in;
logic cond875_write_en;
logic cond875_clk;
logic cond875_reset;
logic cond875_out;
logic cond875_done;
logic cond_wire875_in;
logic cond_wire875_out;
logic cond876_in;
logic cond876_write_en;
logic cond876_clk;
logic cond876_reset;
logic cond876_out;
logic cond876_done;
logic cond_wire876_in;
logic cond_wire876_out;
logic cond877_in;
logic cond877_write_en;
logic cond877_clk;
logic cond877_reset;
logic cond877_out;
logic cond877_done;
logic cond_wire877_in;
logic cond_wire877_out;
logic cond878_in;
logic cond878_write_en;
logic cond878_clk;
logic cond878_reset;
logic cond878_out;
logic cond878_done;
logic cond_wire878_in;
logic cond_wire878_out;
logic cond879_in;
logic cond879_write_en;
logic cond879_clk;
logic cond879_reset;
logic cond879_out;
logic cond879_done;
logic cond_wire879_in;
logic cond_wire879_out;
logic cond880_in;
logic cond880_write_en;
logic cond880_clk;
logic cond880_reset;
logic cond880_out;
logic cond880_done;
logic cond_wire880_in;
logic cond_wire880_out;
logic cond881_in;
logic cond881_write_en;
logic cond881_clk;
logic cond881_reset;
logic cond881_out;
logic cond881_done;
logic cond_wire881_in;
logic cond_wire881_out;
logic cond882_in;
logic cond882_write_en;
logic cond882_clk;
logic cond882_reset;
logic cond882_out;
logic cond882_done;
logic cond_wire882_in;
logic cond_wire882_out;
logic cond883_in;
logic cond883_write_en;
logic cond883_clk;
logic cond883_reset;
logic cond883_out;
logic cond883_done;
logic cond_wire883_in;
logic cond_wire883_out;
logic cond884_in;
logic cond884_write_en;
logic cond884_clk;
logic cond884_reset;
logic cond884_out;
logic cond884_done;
logic cond_wire884_in;
logic cond_wire884_out;
logic cond885_in;
logic cond885_write_en;
logic cond885_clk;
logic cond885_reset;
logic cond885_out;
logic cond885_done;
logic cond_wire885_in;
logic cond_wire885_out;
logic cond886_in;
logic cond886_write_en;
logic cond886_clk;
logic cond886_reset;
logic cond886_out;
logic cond886_done;
logic cond_wire886_in;
logic cond_wire886_out;
logic cond887_in;
logic cond887_write_en;
logic cond887_clk;
logic cond887_reset;
logic cond887_out;
logic cond887_done;
logic cond_wire887_in;
logic cond_wire887_out;
logic cond888_in;
logic cond888_write_en;
logic cond888_clk;
logic cond888_reset;
logic cond888_out;
logic cond888_done;
logic cond_wire888_in;
logic cond_wire888_out;
logic cond889_in;
logic cond889_write_en;
logic cond889_clk;
logic cond889_reset;
logic cond889_out;
logic cond889_done;
logic cond_wire889_in;
logic cond_wire889_out;
logic cond890_in;
logic cond890_write_en;
logic cond890_clk;
logic cond890_reset;
logic cond890_out;
logic cond890_done;
logic cond_wire890_in;
logic cond_wire890_out;
logic cond891_in;
logic cond891_write_en;
logic cond891_clk;
logic cond891_reset;
logic cond891_out;
logic cond891_done;
logic cond_wire891_in;
logic cond_wire891_out;
logic cond892_in;
logic cond892_write_en;
logic cond892_clk;
logic cond892_reset;
logic cond892_out;
logic cond892_done;
logic cond_wire892_in;
logic cond_wire892_out;
logic cond893_in;
logic cond893_write_en;
logic cond893_clk;
logic cond893_reset;
logic cond893_out;
logic cond893_done;
logic cond_wire893_in;
logic cond_wire893_out;
logic cond894_in;
logic cond894_write_en;
logic cond894_clk;
logic cond894_reset;
logic cond894_out;
logic cond894_done;
logic cond_wire894_in;
logic cond_wire894_out;
logic cond895_in;
logic cond895_write_en;
logic cond895_clk;
logic cond895_reset;
logic cond895_out;
logic cond895_done;
logic cond_wire895_in;
logic cond_wire895_out;
logic cond896_in;
logic cond896_write_en;
logic cond896_clk;
logic cond896_reset;
logic cond896_out;
logic cond896_done;
logic cond_wire896_in;
logic cond_wire896_out;
logic cond897_in;
logic cond897_write_en;
logic cond897_clk;
logic cond897_reset;
logic cond897_out;
logic cond897_done;
logic cond_wire897_in;
logic cond_wire897_out;
logic cond898_in;
logic cond898_write_en;
logic cond898_clk;
logic cond898_reset;
logic cond898_out;
logic cond898_done;
logic cond_wire898_in;
logic cond_wire898_out;
logic cond899_in;
logic cond899_write_en;
logic cond899_clk;
logic cond899_reset;
logic cond899_out;
logic cond899_done;
logic cond_wire899_in;
logic cond_wire899_out;
logic cond900_in;
logic cond900_write_en;
logic cond900_clk;
logic cond900_reset;
logic cond900_out;
logic cond900_done;
logic cond_wire900_in;
logic cond_wire900_out;
logic cond901_in;
logic cond901_write_en;
logic cond901_clk;
logic cond901_reset;
logic cond901_out;
logic cond901_done;
logic cond_wire901_in;
logic cond_wire901_out;
logic cond902_in;
logic cond902_write_en;
logic cond902_clk;
logic cond902_reset;
logic cond902_out;
logic cond902_done;
logic cond_wire902_in;
logic cond_wire902_out;
logic cond903_in;
logic cond903_write_en;
logic cond903_clk;
logic cond903_reset;
logic cond903_out;
logic cond903_done;
logic cond_wire903_in;
logic cond_wire903_out;
logic cond904_in;
logic cond904_write_en;
logic cond904_clk;
logic cond904_reset;
logic cond904_out;
logic cond904_done;
logic cond_wire904_in;
logic cond_wire904_out;
logic cond905_in;
logic cond905_write_en;
logic cond905_clk;
logic cond905_reset;
logic cond905_out;
logic cond905_done;
logic cond_wire905_in;
logic cond_wire905_out;
logic cond906_in;
logic cond906_write_en;
logic cond906_clk;
logic cond906_reset;
logic cond906_out;
logic cond906_done;
logic cond_wire906_in;
logic cond_wire906_out;
logic cond907_in;
logic cond907_write_en;
logic cond907_clk;
logic cond907_reset;
logic cond907_out;
logic cond907_done;
logic cond_wire907_in;
logic cond_wire907_out;
logic cond908_in;
logic cond908_write_en;
logic cond908_clk;
logic cond908_reset;
logic cond908_out;
logic cond908_done;
logic cond_wire908_in;
logic cond_wire908_out;
logic cond909_in;
logic cond909_write_en;
logic cond909_clk;
logic cond909_reset;
logic cond909_out;
logic cond909_done;
logic cond_wire909_in;
logic cond_wire909_out;
logic cond910_in;
logic cond910_write_en;
logic cond910_clk;
logic cond910_reset;
logic cond910_out;
logic cond910_done;
logic cond_wire910_in;
logic cond_wire910_out;
logic cond911_in;
logic cond911_write_en;
logic cond911_clk;
logic cond911_reset;
logic cond911_out;
logic cond911_done;
logic cond_wire911_in;
logic cond_wire911_out;
logic cond912_in;
logic cond912_write_en;
logic cond912_clk;
logic cond912_reset;
logic cond912_out;
logic cond912_done;
logic cond_wire912_in;
logic cond_wire912_out;
logic cond913_in;
logic cond913_write_en;
logic cond913_clk;
logic cond913_reset;
logic cond913_out;
logic cond913_done;
logic cond_wire913_in;
logic cond_wire913_out;
logic cond914_in;
logic cond914_write_en;
logic cond914_clk;
logic cond914_reset;
logic cond914_out;
logic cond914_done;
logic cond_wire914_in;
logic cond_wire914_out;
logic cond915_in;
logic cond915_write_en;
logic cond915_clk;
logic cond915_reset;
logic cond915_out;
logic cond915_done;
logic cond_wire915_in;
logic cond_wire915_out;
logic cond916_in;
logic cond916_write_en;
logic cond916_clk;
logic cond916_reset;
logic cond916_out;
logic cond916_done;
logic cond_wire916_in;
logic cond_wire916_out;
logic cond917_in;
logic cond917_write_en;
logic cond917_clk;
logic cond917_reset;
logic cond917_out;
logic cond917_done;
logic cond_wire917_in;
logic cond_wire917_out;
logic cond918_in;
logic cond918_write_en;
logic cond918_clk;
logic cond918_reset;
logic cond918_out;
logic cond918_done;
logic cond_wire918_in;
logic cond_wire918_out;
logic cond919_in;
logic cond919_write_en;
logic cond919_clk;
logic cond919_reset;
logic cond919_out;
logic cond919_done;
logic cond_wire919_in;
logic cond_wire919_out;
logic cond920_in;
logic cond920_write_en;
logic cond920_clk;
logic cond920_reset;
logic cond920_out;
logic cond920_done;
logic cond_wire920_in;
logic cond_wire920_out;
logic cond921_in;
logic cond921_write_en;
logic cond921_clk;
logic cond921_reset;
logic cond921_out;
logic cond921_done;
logic cond_wire921_in;
logic cond_wire921_out;
logic cond922_in;
logic cond922_write_en;
logic cond922_clk;
logic cond922_reset;
logic cond922_out;
logic cond922_done;
logic cond_wire922_in;
logic cond_wire922_out;
logic cond923_in;
logic cond923_write_en;
logic cond923_clk;
logic cond923_reset;
logic cond923_out;
logic cond923_done;
logic cond_wire923_in;
logic cond_wire923_out;
logic cond924_in;
logic cond924_write_en;
logic cond924_clk;
logic cond924_reset;
logic cond924_out;
logic cond924_done;
logic cond_wire924_in;
logic cond_wire924_out;
logic cond925_in;
logic cond925_write_en;
logic cond925_clk;
logic cond925_reset;
logic cond925_out;
logic cond925_done;
logic cond_wire925_in;
logic cond_wire925_out;
logic cond926_in;
logic cond926_write_en;
logic cond926_clk;
logic cond926_reset;
logic cond926_out;
logic cond926_done;
logic cond_wire926_in;
logic cond_wire926_out;
logic cond927_in;
logic cond927_write_en;
logic cond927_clk;
logic cond927_reset;
logic cond927_out;
logic cond927_done;
logic cond_wire927_in;
logic cond_wire927_out;
logic cond928_in;
logic cond928_write_en;
logic cond928_clk;
logic cond928_reset;
logic cond928_out;
logic cond928_done;
logic cond_wire928_in;
logic cond_wire928_out;
logic cond929_in;
logic cond929_write_en;
logic cond929_clk;
logic cond929_reset;
logic cond929_out;
logic cond929_done;
logic cond_wire929_in;
logic cond_wire929_out;
logic cond930_in;
logic cond930_write_en;
logic cond930_clk;
logic cond930_reset;
logic cond930_out;
logic cond930_done;
logic cond_wire930_in;
logic cond_wire930_out;
logic cond931_in;
logic cond931_write_en;
logic cond931_clk;
logic cond931_reset;
logic cond931_out;
logic cond931_done;
logic cond_wire931_in;
logic cond_wire931_out;
logic cond932_in;
logic cond932_write_en;
logic cond932_clk;
logic cond932_reset;
logic cond932_out;
logic cond932_done;
logic cond_wire932_in;
logic cond_wire932_out;
logic cond933_in;
logic cond933_write_en;
logic cond933_clk;
logic cond933_reset;
logic cond933_out;
logic cond933_done;
logic cond_wire933_in;
logic cond_wire933_out;
logic cond934_in;
logic cond934_write_en;
logic cond934_clk;
logic cond934_reset;
logic cond934_out;
logic cond934_done;
logic cond_wire934_in;
logic cond_wire934_out;
logic cond935_in;
logic cond935_write_en;
logic cond935_clk;
logic cond935_reset;
logic cond935_out;
logic cond935_done;
logic cond_wire935_in;
logic cond_wire935_out;
logic cond936_in;
logic cond936_write_en;
logic cond936_clk;
logic cond936_reset;
logic cond936_out;
logic cond936_done;
logic cond_wire936_in;
logic cond_wire936_out;
logic cond937_in;
logic cond937_write_en;
logic cond937_clk;
logic cond937_reset;
logic cond937_out;
logic cond937_done;
logic cond_wire937_in;
logic cond_wire937_out;
logic cond938_in;
logic cond938_write_en;
logic cond938_clk;
logic cond938_reset;
logic cond938_out;
logic cond938_done;
logic cond_wire938_in;
logic cond_wire938_out;
logic cond939_in;
logic cond939_write_en;
logic cond939_clk;
logic cond939_reset;
logic cond939_out;
logic cond939_done;
logic cond_wire939_in;
logic cond_wire939_out;
logic cond940_in;
logic cond940_write_en;
logic cond940_clk;
logic cond940_reset;
logic cond940_out;
logic cond940_done;
logic cond_wire940_in;
logic cond_wire940_out;
logic cond941_in;
logic cond941_write_en;
logic cond941_clk;
logic cond941_reset;
logic cond941_out;
logic cond941_done;
logic cond_wire941_in;
logic cond_wire941_out;
logic cond942_in;
logic cond942_write_en;
logic cond942_clk;
logic cond942_reset;
logic cond942_out;
logic cond942_done;
logic cond_wire942_in;
logic cond_wire942_out;
logic cond943_in;
logic cond943_write_en;
logic cond943_clk;
logic cond943_reset;
logic cond943_out;
logic cond943_done;
logic cond_wire943_in;
logic cond_wire943_out;
logic cond944_in;
logic cond944_write_en;
logic cond944_clk;
logic cond944_reset;
logic cond944_out;
logic cond944_done;
logic cond_wire944_in;
logic cond_wire944_out;
logic cond945_in;
logic cond945_write_en;
logic cond945_clk;
logic cond945_reset;
logic cond945_out;
logic cond945_done;
logic cond_wire945_in;
logic cond_wire945_out;
logic cond946_in;
logic cond946_write_en;
logic cond946_clk;
logic cond946_reset;
logic cond946_out;
logic cond946_done;
logic cond_wire946_in;
logic cond_wire946_out;
logic cond947_in;
logic cond947_write_en;
logic cond947_clk;
logic cond947_reset;
logic cond947_out;
logic cond947_done;
logic cond_wire947_in;
logic cond_wire947_out;
logic cond948_in;
logic cond948_write_en;
logic cond948_clk;
logic cond948_reset;
logic cond948_out;
logic cond948_done;
logic cond_wire948_in;
logic cond_wire948_out;
logic cond949_in;
logic cond949_write_en;
logic cond949_clk;
logic cond949_reset;
logic cond949_out;
logic cond949_done;
logic cond_wire949_in;
logic cond_wire949_out;
logic cond950_in;
logic cond950_write_en;
logic cond950_clk;
logic cond950_reset;
logic cond950_out;
logic cond950_done;
logic cond_wire950_in;
logic cond_wire950_out;
logic cond951_in;
logic cond951_write_en;
logic cond951_clk;
logic cond951_reset;
logic cond951_out;
logic cond951_done;
logic cond_wire951_in;
logic cond_wire951_out;
logic cond952_in;
logic cond952_write_en;
logic cond952_clk;
logic cond952_reset;
logic cond952_out;
logic cond952_done;
logic cond_wire952_in;
logic cond_wire952_out;
logic cond953_in;
logic cond953_write_en;
logic cond953_clk;
logic cond953_reset;
logic cond953_out;
logic cond953_done;
logic cond_wire953_in;
logic cond_wire953_out;
logic cond954_in;
logic cond954_write_en;
logic cond954_clk;
logic cond954_reset;
logic cond954_out;
logic cond954_done;
logic cond_wire954_in;
logic cond_wire954_out;
logic cond955_in;
logic cond955_write_en;
logic cond955_clk;
logic cond955_reset;
logic cond955_out;
logic cond955_done;
logic cond_wire955_in;
logic cond_wire955_out;
logic cond956_in;
logic cond956_write_en;
logic cond956_clk;
logic cond956_reset;
logic cond956_out;
logic cond956_done;
logic cond_wire956_in;
logic cond_wire956_out;
logic cond957_in;
logic cond957_write_en;
logic cond957_clk;
logic cond957_reset;
logic cond957_out;
logic cond957_done;
logic cond_wire957_in;
logic cond_wire957_out;
logic cond958_in;
logic cond958_write_en;
logic cond958_clk;
logic cond958_reset;
logic cond958_out;
logic cond958_done;
logic cond_wire958_in;
logic cond_wire958_out;
logic cond959_in;
logic cond959_write_en;
logic cond959_clk;
logic cond959_reset;
logic cond959_out;
logic cond959_done;
logic cond_wire959_in;
logic cond_wire959_out;
logic cond960_in;
logic cond960_write_en;
logic cond960_clk;
logic cond960_reset;
logic cond960_out;
logic cond960_done;
logic cond_wire960_in;
logic cond_wire960_out;
logic cond961_in;
logic cond961_write_en;
logic cond961_clk;
logic cond961_reset;
logic cond961_out;
logic cond961_done;
logic cond_wire961_in;
logic cond_wire961_out;
logic cond962_in;
logic cond962_write_en;
logic cond962_clk;
logic cond962_reset;
logic cond962_out;
logic cond962_done;
logic cond_wire962_in;
logic cond_wire962_out;
logic cond963_in;
logic cond963_write_en;
logic cond963_clk;
logic cond963_reset;
logic cond963_out;
logic cond963_done;
logic cond_wire963_in;
logic cond_wire963_out;
logic cond964_in;
logic cond964_write_en;
logic cond964_clk;
logic cond964_reset;
logic cond964_out;
logic cond964_done;
logic cond_wire964_in;
logic cond_wire964_out;
logic cond965_in;
logic cond965_write_en;
logic cond965_clk;
logic cond965_reset;
logic cond965_out;
logic cond965_done;
logic cond_wire965_in;
logic cond_wire965_out;
logic cond966_in;
logic cond966_write_en;
logic cond966_clk;
logic cond966_reset;
logic cond966_out;
logic cond966_done;
logic cond_wire966_in;
logic cond_wire966_out;
logic cond967_in;
logic cond967_write_en;
logic cond967_clk;
logic cond967_reset;
logic cond967_out;
logic cond967_done;
logic cond_wire967_in;
logic cond_wire967_out;
logic cond968_in;
logic cond968_write_en;
logic cond968_clk;
logic cond968_reset;
logic cond968_out;
logic cond968_done;
logic cond_wire968_in;
logic cond_wire968_out;
logic cond969_in;
logic cond969_write_en;
logic cond969_clk;
logic cond969_reset;
logic cond969_out;
logic cond969_done;
logic cond_wire969_in;
logic cond_wire969_out;
logic cond970_in;
logic cond970_write_en;
logic cond970_clk;
logic cond970_reset;
logic cond970_out;
logic cond970_done;
logic cond_wire970_in;
logic cond_wire970_out;
logic cond971_in;
logic cond971_write_en;
logic cond971_clk;
logic cond971_reset;
logic cond971_out;
logic cond971_done;
logic cond_wire971_in;
logic cond_wire971_out;
logic cond972_in;
logic cond972_write_en;
logic cond972_clk;
logic cond972_reset;
logic cond972_out;
logic cond972_done;
logic cond_wire972_in;
logic cond_wire972_out;
logic cond973_in;
logic cond973_write_en;
logic cond973_clk;
logic cond973_reset;
logic cond973_out;
logic cond973_done;
logic cond_wire973_in;
logic cond_wire973_out;
logic cond974_in;
logic cond974_write_en;
logic cond974_clk;
logic cond974_reset;
logic cond974_out;
logic cond974_done;
logic cond_wire974_in;
logic cond_wire974_out;
logic cond975_in;
logic cond975_write_en;
logic cond975_clk;
logic cond975_reset;
logic cond975_out;
logic cond975_done;
logic cond_wire975_in;
logic cond_wire975_out;
logic cond976_in;
logic cond976_write_en;
logic cond976_clk;
logic cond976_reset;
logic cond976_out;
logic cond976_done;
logic cond_wire976_in;
logic cond_wire976_out;
logic cond977_in;
logic cond977_write_en;
logic cond977_clk;
logic cond977_reset;
logic cond977_out;
logic cond977_done;
logic cond_wire977_in;
logic cond_wire977_out;
logic cond978_in;
logic cond978_write_en;
logic cond978_clk;
logic cond978_reset;
logic cond978_out;
logic cond978_done;
logic cond_wire978_in;
logic cond_wire978_out;
logic cond979_in;
logic cond979_write_en;
logic cond979_clk;
logic cond979_reset;
logic cond979_out;
logic cond979_done;
logic cond_wire979_in;
logic cond_wire979_out;
logic cond980_in;
logic cond980_write_en;
logic cond980_clk;
logic cond980_reset;
logic cond980_out;
logic cond980_done;
logic cond_wire980_in;
logic cond_wire980_out;
logic cond981_in;
logic cond981_write_en;
logic cond981_clk;
logic cond981_reset;
logic cond981_out;
logic cond981_done;
logic cond_wire981_in;
logic cond_wire981_out;
logic cond982_in;
logic cond982_write_en;
logic cond982_clk;
logic cond982_reset;
logic cond982_out;
logic cond982_done;
logic cond_wire982_in;
logic cond_wire982_out;
logic cond983_in;
logic cond983_write_en;
logic cond983_clk;
logic cond983_reset;
logic cond983_out;
logic cond983_done;
logic cond_wire983_in;
logic cond_wire983_out;
logic cond984_in;
logic cond984_write_en;
logic cond984_clk;
logic cond984_reset;
logic cond984_out;
logic cond984_done;
logic cond_wire984_in;
logic cond_wire984_out;
logic cond985_in;
logic cond985_write_en;
logic cond985_clk;
logic cond985_reset;
logic cond985_out;
logic cond985_done;
logic cond_wire985_in;
logic cond_wire985_out;
logic cond986_in;
logic cond986_write_en;
logic cond986_clk;
logic cond986_reset;
logic cond986_out;
logic cond986_done;
logic cond_wire986_in;
logic cond_wire986_out;
logic cond987_in;
logic cond987_write_en;
logic cond987_clk;
logic cond987_reset;
logic cond987_out;
logic cond987_done;
logic cond_wire987_in;
logic cond_wire987_out;
logic cond988_in;
logic cond988_write_en;
logic cond988_clk;
logic cond988_reset;
logic cond988_out;
logic cond988_done;
logic cond_wire988_in;
logic cond_wire988_out;
logic cond989_in;
logic cond989_write_en;
logic cond989_clk;
logic cond989_reset;
logic cond989_out;
logic cond989_done;
logic cond_wire989_in;
logic cond_wire989_out;
logic cond990_in;
logic cond990_write_en;
logic cond990_clk;
logic cond990_reset;
logic cond990_out;
logic cond990_done;
logic cond_wire990_in;
logic cond_wire990_out;
logic cond991_in;
logic cond991_write_en;
logic cond991_clk;
logic cond991_reset;
logic cond991_out;
logic cond991_done;
logic cond_wire991_in;
logic cond_wire991_out;
logic cond992_in;
logic cond992_write_en;
logic cond992_clk;
logic cond992_reset;
logic cond992_out;
logic cond992_done;
logic cond_wire992_in;
logic cond_wire992_out;
logic cond993_in;
logic cond993_write_en;
logic cond993_clk;
logic cond993_reset;
logic cond993_out;
logic cond993_done;
logic cond_wire993_in;
logic cond_wire993_out;
logic cond994_in;
logic cond994_write_en;
logic cond994_clk;
logic cond994_reset;
logic cond994_out;
logic cond994_done;
logic cond_wire994_in;
logic cond_wire994_out;
logic cond995_in;
logic cond995_write_en;
logic cond995_clk;
logic cond995_reset;
logic cond995_out;
logic cond995_done;
logic cond_wire995_in;
logic cond_wire995_out;
logic cond996_in;
logic cond996_write_en;
logic cond996_clk;
logic cond996_reset;
logic cond996_out;
logic cond996_done;
logic cond_wire996_in;
logic cond_wire996_out;
logic cond997_in;
logic cond997_write_en;
logic cond997_clk;
logic cond997_reset;
logic cond997_out;
logic cond997_done;
logic cond_wire997_in;
logic cond_wire997_out;
logic cond998_in;
logic cond998_write_en;
logic cond998_clk;
logic cond998_reset;
logic cond998_out;
logic cond998_done;
logic cond_wire998_in;
logic cond_wire998_out;
logic cond999_in;
logic cond999_write_en;
logic cond999_clk;
logic cond999_reset;
logic cond999_out;
logic cond999_done;
logic cond_wire999_in;
logic cond_wire999_out;
logic cond1000_in;
logic cond1000_write_en;
logic cond1000_clk;
logic cond1000_reset;
logic cond1000_out;
logic cond1000_done;
logic cond_wire1000_in;
logic cond_wire1000_out;
logic cond1001_in;
logic cond1001_write_en;
logic cond1001_clk;
logic cond1001_reset;
logic cond1001_out;
logic cond1001_done;
logic cond_wire1001_in;
logic cond_wire1001_out;
logic cond1002_in;
logic cond1002_write_en;
logic cond1002_clk;
logic cond1002_reset;
logic cond1002_out;
logic cond1002_done;
logic cond_wire1002_in;
logic cond_wire1002_out;
logic cond1003_in;
logic cond1003_write_en;
logic cond1003_clk;
logic cond1003_reset;
logic cond1003_out;
logic cond1003_done;
logic cond_wire1003_in;
logic cond_wire1003_out;
logic cond1004_in;
logic cond1004_write_en;
logic cond1004_clk;
logic cond1004_reset;
logic cond1004_out;
logic cond1004_done;
logic cond_wire1004_in;
logic cond_wire1004_out;
logic cond1005_in;
logic cond1005_write_en;
logic cond1005_clk;
logic cond1005_reset;
logic cond1005_out;
logic cond1005_done;
logic cond_wire1005_in;
logic cond_wire1005_out;
logic cond1006_in;
logic cond1006_write_en;
logic cond1006_clk;
logic cond1006_reset;
logic cond1006_out;
logic cond1006_done;
logic cond_wire1006_in;
logic cond_wire1006_out;
logic cond1007_in;
logic cond1007_write_en;
logic cond1007_clk;
logic cond1007_reset;
logic cond1007_out;
logic cond1007_done;
logic cond_wire1007_in;
logic cond_wire1007_out;
logic cond1008_in;
logic cond1008_write_en;
logic cond1008_clk;
logic cond1008_reset;
logic cond1008_out;
logic cond1008_done;
logic cond_wire1008_in;
logic cond_wire1008_out;
logic cond1009_in;
logic cond1009_write_en;
logic cond1009_clk;
logic cond1009_reset;
logic cond1009_out;
logic cond1009_done;
logic cond_wire1009_in;
logic cond_wire1009_out;
logic cond1010_in;
logic cond1010_write_en;
logic cond1010_clk;
logic cond1010_reset;
logic cond1010_out;
logic cond1010_done;
logic cond_wire1010_in;
logic cond_wire1010_out;
logic cond1011_in;
logic cond1011_write_en;
logic cond1011_clk;
logic cond1011_reset;
logic cond1011_out;
logic cond1011_done;
logic cond_wire1011_in;
logic cond_wire1011_out;
logic cond1012_in;
logic cond1012_write_en;
logic cond1012_clk;
logic cond1012_reset;
logic cond1012_out;
logic cond1012_done;
logic cond_wire1012_in;
logic cond_wire1012_out;
logic cond1013_in;
logic cond1013_write_en;
logic cond1013_clk;
logic cond1013_reset;
logic cond1013_out;
logic cond1013_done;
logic cond_wire1013_in;
logic cond_wire1013_out;
logic cond1014_in;
logic cond1014_write_en;
logic cond1014_clk;
logic cond1014_reset;
logic cond1014_out;
logic cond1014_done;
logic cond_wire1014_in;
logic cond_wire1014_out;
logic cond1015_in;
logic cond1015_write_en;
logic cond1015_clk;
logic cond1015_reset;
logic cond1015_out;
logic cond1015_done;
logic cond_wire1015_in;
logic cond_wire1015_out;
logic cond1016_in;
logic cond1016_write_en;
logic cond1016_clk;
logic cond1016_reset;
logic cond1016_out;
logic cond1016_done;
logic cond_wire1016_in;
logic cond_wire1016_out;
logic cond1017_in;
logic cond1017_write_en;
logic cond1017_clk;
logic cond1017_reset;
logic cond1017_out;
logic cond1017_done;
logic cond_wire1017_in;
logic cond_wire1017_out;
logic cond1018_in;
logic cond1018_write_en;
logic cond1018_clk;
logic cond1018_reset;
logic cond1018_out;
logic cond1018_done;
logic cond_wire1018_in;
logic cond_wire1018_out;
logic cond1019_in;
logic cond1019_write_en;
logic cond1019_clk;
logic cond1019_reset;
logic cond1019_out;
logic cond1019_done;
logic cond_wire1019_in;
logic cond_wire1019_out;
logic cond1020_in;
logic cond1020_write_en;
logic cond1020_clk;
logic cond1020_reset;
logic cond1020_out;
logic cond1020_done;
logic cond_wire1020_in;
logic cond_wire1020_out;
logic cond1021_in;
logic cond1021_write_en;
logic cond1021_clk;
logic cond1021_reset;
logic cond1021_out;
logic cond1021_done;
logic cond_wire1021_in;
logic cond_wire1021_out;
logic cond1022_in;
logic cond1022_write_en;
logic cond1022_clk;
logic cond1022_reset;
logic cond1022_out;
logic cond1022_done;
logic cond_wire1022_in;
logic cond_wire1022_out;
logic cond1023_in;
logic cond1023_write_en;
logic cond1023_clk;
logic cond1023_reset;
logic cond1023_out;
logic cond1023_done;
logic cond_wire1023_in;
logic cond_wire1023_out;
logic cond1024_in;
logic cond1024_write_en;
logic cond1024_clk;
logic cond1024_reset;
logic cond1024_out;
logic cond1024_done;
logic cond_wire1024_in;
logic cond_wire1024_out;
logic cond1025_in;
logic cond1025_write_en;
logic cond1025_clk;
logic cond1025_reset;
logic cond1025_out;
logic cond1025_done;
logic cond_wire1025_in;
logic cond_wire1025_out;
logic cond1026_in;
logic cond1026_write_en;
logic cond1026_clk;
logic cond1026_reset;
logic cond1026_out;
logic cond1026_done;
logic cond_wire1026_in;
logic cond_wire1026_out;
logic cond1027_in;
logic cond1027_write_en;
logic cond1027_clk;
logic cond1027_reset;
logic cond1027_out;
logic cond1027_done;
logic cond_wire1027_in;
logic cond_wire1027_out;
logic cond1028_in;
logic cond1028_write_en;
logic cond1028_clk;
logic cond1028_reset;
logic cond1028_out;
logic cond1028_done;
logic cond_wire1028_in;
logic cond_wire1028_out;
logic cond1029_in;
logic cond1029_write_en;
logic cond1029_clk;
logic cond1029_reset;
logic cond1029_out;
logic cond1029_done;
logic cond_wire1029_in;
logic cond_wire1029_out;
logic cond1030_in;
logic cond1030_write_en;
logic cond1030_clk;
logic cond1030_reset;
logic cond1030_out;
logic cond1030_done;
logic cond_wire1030_in;
logic cond_wire1030_out;
logic cond1031_in;
logic cond1031_write_en;
logic cond1031_clk;
logic cond1031_reset;
logic cond1031_out;
logic cond1031_done;
logic cond_wire1031_in;
logic cond_wire1031_out;
logic cond1032_in;
logic cond1032_write_en;
logic cond1032_clk;
logic cond1032_reset;
logic cond1032_out;
logic cond1032_done;
logic cond_wire1032_in;
logic cond_wire1032_out;
logic cond1033_in;
logic cond1033_write_en;
logic cond1033_clk;
logic cond1033_reset;
logic cond1033_out;
logic cond1033_done;
logic cond_wire1033_in;
logic cond_wire1033_out;
logic cond1034_in;
logic cond1034_write_en;
logic cond1034_clk;
logic cond1034_reset;
logic cond1034_out;
logic cond1034_done;
logic cond_wire1034_in;
logic cond_wire1034_out;
logic cond1035_in;
logic cond1035_write_en;
logic cond1035_clk;
logic cond1035_reset;
logic cond1035_out;
logic cond1035_done;
logic cond_wire1035_in;
logic cond_wire1035_out;
logic cond1036_in;
logic cond1036_write_en;
logic cond1036_clk;
logic cond1036_reset;
logic cond1036_out;
logic cond1036_done;
logic cond_wire1036_in;
logic cond_wire1036_out;
logic cond1037_in;
logic cond1037_write_en;
logic cond1037_clk;
logic cond1037_reset;
logic cond1037_out;
logic cond1037_done;
logic cond_wire1037_in;
logic cond_wire1037_out;
logic cond1038_in;
logic cond1038_write_en;
logic cond1038_clk;
logic cond1038_reset;
logic cond1038_out;
logic cond1038_done;
logic cond_wire1038_in;
logic cond_wire1038_out;
logic cond1039_in;
logic cond1039_write_en;
logic cond1039_clk;
logic cond1039_reset;
logic cond1039_out;
logic cond1039_done;
logic cond_wire1039_in;
logic cond_wire1039_out;
logic cond1040_in;
logic cond1040_write_en;
logic cond1040_clk;
logic cond1040_reset;
logic cond1040_out;
logic cond1040_done;
logic cond_wire1040_in;
logic cond_wire1040_out;
logic cond1041_in;
logic cond1041_write_en;
logic cond1041_clk;
logic cond1041_reset;
logic cond1041_out;
logic cond1041_done;
logic cond_wire1041_in;
logic cond_wire1041_out;
logic cond1042_in;
logic cond1042_write_en;
logic cond1042_clk;
logic cond1042_reset;
logic cond1042_out;
logic cond1042_done;
logic cond_wire1042_in;
logic cond_wire1042_out;
logic cond1043_in;
logic cond1043_write_en;
logic cond1043_clk;
logic cond1043_reset;
logic cond1043_out;
logic cond1043_done;
logic cond_wire1043_in;
logic cond_wire1043_out;
logic cond1044_in;
logic cond1044_write_en;
logic cond1044_clk;
logic cond1044_reset;
logic cond1044_out;
logic cond1044_done;
logic cond_wire1044_in;
logic cond_wire1044_out;
logic cond1045_in;
logic cond1045_write_en;
logic cond1045_clk;
logic cond1045_reset;
logic cond1045_out;
logic cond1045_done;
logic cond_wire1045_in;
logic cond_wire1045_out;
logic cond1046_in;
logic cond1046_write_en;
logic cond1046_clk;
logic cond1046_reset;
logic cond1046_out;
logic cond1046_done;
logic cond_wire1046_in;
logic cond_wire1046_out;
logic cond1047_in;
logic cond1047_write_en;
logic cond1047_clk;
logic cond1047_reset;
logic cond1047_out;
logic cond1047_done;
logic cond_wire1047_in;
logic cond_wire1047_out;
logic cond1048_in;
logic cond1048_write_en;
logic cond1048_clk;
logic cond1048_reset;
logic cond1048_out;
logic cond1048_done;
logic cond_wire1048_in;
logic cond_wire1048_out;
logic cond1049_in;
logic cond1049_write_en;
logic cond1049_clk;
logic cond1049_reset;
logic cond1049_out;
logic cond1049_done;
logic cond_wire1049_in;
logic cond_wire1049_out;
logic cond1050_in;
logic cond1050_write_en;
logic cond1050_clk;
logic cond1050_reset;
logic cond1050_out;
logic cond1050_done;
logic cond_wire1050_in;
logic cond_wire1050_out;
logic cond1051_in;
logic cond1051_write_en;
logic cond1051_clk;
logic cond1051_reset;
logic cond1051_out;
logic cond1051_done;
logic cond_wire1051_in;
logic cond_wire1051_out;
logic cond1052_in;
logic cond1052_write_en;
logic cond1052_clk;
logic cond1052_reset;
logic cond1052_out;
logic cond1052_done;
logic cond_wire1052_in;
logic cond_wire1052_out;
logic fsm_in;
logic fsm_write_en;
logic fsm_clk;
logic fsm_reset;
logic fsm_out;
logic fsm_done;
logic [5:0] fsm0_in;
logic fsm0_write_en;
logic fsm0_clk;
logic fsm0_reset;
logic [5:0] fsm0_out;
logic fsm0_done;
logic ud_out;
logic [5:0] adder_left;
logic [5:0] adder_right;
logic [5:0] adder_out;
logic ud0_out;
logic adder0_left;
logic adder0_right;
logic adder0_out;
logic signal_reg_in;
logic signal_reg_write_en;
logic signal_reg_clk;
logic signal_reg_reset;
logic signal_reg_out;
logic signal_reg_done;
logic early_reset_static_seq_go_in;
logic early_reset_static_seq_go_out;
logic early_reset_static_seq_done_in;
logic early_reset_static_seq_done_out;
logic early_reset_static_par0_go_in;
logic early_reset_static_par0_go_out;
logic early_reset_static_par0_done_in;
logic early_reset_static_par0_done_out;
logic wrapper_early_reset_static_seq_go_in;
logic wrapper_early_reset_static_seq_go_out;
logic wrapper_early_reset_static_seq_done_in;
logic wrapper_early_reset_static_seq_done_out;
mac_pe pe_0_0 (
    .clk(pe_0_0_clk),
    .done(pe_0_0_done),
    .go(pe_0_0_go),
    .left(pe_0_0_left),
    .mul_ready(pe_0_0_mul_ready),
    .out(pe_0_0_out),
    .reset(pe_0_0_reset),
    .top(pe_0_0_top)
);
std_reg # (
    .WIDTH(32)
) top_0_0 (
    .clk(top_0_0_clk),
    .done(top_0_0_done),
    .in(top_0_0_in),
    .out(top_0_0_out),
    .reset(top_0_0_reset),
    .write_en(top_0_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_0 (
    .clk(left_0_0_clk),
    .done(left_0_0_done),
    .in(left_0_0_in),
    .out(left_0_0_out),
    .reset(left_0_0_reset),
    .write_en(left_0_0_write_en)
);
mac_pe pe_0_1 (
    .clk(pe_0_1_clk),
    .done(pe_0_1_done),
    .go(pe_0_1_go),
    .left(pe_0_1_left),
    .mul_ready(pe_0_1_mul_ready),
    .out(pe_0_1_out),
    .reset(pe_0_1_reset),
    .top(pe_0_1_top)
);
std_reg # (
    .WIDTH(32)
) top_0_1 (
    .clk(top_0_1_clk),
    .done(top_0_1_done),
    .in(top_0_1_in),
    .out(top_0_1_out),
    .reset(top_0_1_reset),
    .write_en(top_0_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_1 (
    .clk(left_0_1_clk),
    .done(left_0_1_done),
    .in(left_0_1_in),
    .out(left_0_1_out),
    .reset(left_0_1_reset),
    .write_en(left_0_1_write_en)
);
mac_pe pe_0_2 (
    .clk(pe_0_2_clk),
    .done(pe_0_2_done),
    .go(pe_0_2_go),
    .left(pe_0_2_left),
    .mul_ready(pe_0_2_mul_ready),
    .out(pe_0_2_out),
    .reset(pe_0_2_reset),
    .top(pe_0_2_top)
);
std_reg # (
    .WIDTH(32)
) top_0_2 (
    .clk(top_0_2_clk),
    .done(top_0_2_done),
    .in(top_0_2_in),
    .out(top_0_2_out),
    .reset(top_0_2_reset),
    .write_en(top_0_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_2 (
    .clk(left_0_2_clk),
    .done(left_0_2_done),
    .in(left_0_2_in),
    .out(left_0_2_out),
    .reset(left_0_2_reset),
    .write_en(left_0_2_write_en)
);
mac_pe pe_0_3 (
    .clk(pe_0_3_clk),
    .done(pe_0_3_done),
    .go(pe_0_3_go),
    .left(pe_0_3_left),
    .mul_ready(pe_0_3_mul_ready),
    .out(pe_0_3_out),
    .reset(pe_0_3_reset),
    .top(pe_0_3_top)
);
std_reg # (
    .WIDTH(32)
) top_0_3 (
    .clk(top_0_3_clk),
    .done(top_0_3_done),
    .in(top_0_3_in),
    .out(top_0_3_out),
    .reset(top_0_3_reset),
    .write_en(top_0_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_3 (
    .clk(left_0_3_clk),
    .done(left_0_3_done),
    .in(left_0_3_in),
    .out(left_0_3_out),
    .reset(left_0_3_reset),
    .write_en(left_0_3_write_en)
);
mac_pe pe_0_4 (
    .clk(pe_0_4_clk),
    .done(pe_0_4_done),
    .go(pe_0_4_go),
    .left(pe_0_4_left),
    .mul_ready(pe_0_4_mul_ready),
    .out(pe_0_4_out),
    .reset(pe_0_4_reset),
    .top(pe_0_4_top)
);
std_reg # (
    .WIDTH(32)
) top_0_4 (
    .clk(top_0_4_clk),
    .done(top_0_4_done),
    .in(top_0_4_in),
    .out(top_0_4_out),
    .reset(top_0_4_reset),
    .write_en(top_0_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_4 (
    .clk(left_0_4_clk),
    .done(left_0_4_done),
    .in(left_0_4_in),
    .out(left_0_4_out),
    .reset(left_0_4_reset),
    .write_en(left_0_4_write_en)
);
mac_pe pe_0_5 (
    .clk(pe_0_5_clk),
    .done(pe_0_5_done),
    .go(pe_0_5_go),
    .left(pe_0_5_left),
    .mul_ready(pe_0_5_mul_ready),
    .out(pe_0_5_out),
    .reset(pe_0_5_reset),
    .top(pe_0_5_top)
);
std_reg # (
    .WIDTH(32)
) top_0_5 (
    .clk(top_0_5_clk),
    .done(top_0_5_done),
    .in(top_0_5_in),
    .out(top_0_5_out),
    .reset(top_0_5_reset),
    .write_en(top_0_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_5 (
    .clk(left_0_5_clk),
    .done(left_0_5_done),
    .in(left_0_5_in),
    .out(left_0_5_out),
    .reset(left_0_5_reset),
    .write_en(left_0_5_write_en)
);
mac_pe pe_0_6 (
    .clk(pe_0_6_clk),
    .done(pe_0_6_done),
    .go(pe_0_6_go),
    .left(pe_0_6_left),
    .mul_ready(pe_0_6_mul_ready),
    .out(pe_0_6_out),
    .reset(pe_0_6_reset),
    .top(pe_0_6_top)
);
std_reg # (
    .WIDTH(32)
) top_0_6 (
    .clk(top_0_6_clk),
    .done(top_0_6_done),
    .in(top_0_6_in),
    .out(top_0_6_out),
    .reset(top_0_6_reset),
    .write_en(top_0_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_6 (
    .clk(left_0_6_clk),
    .done(left_0_6_done),
    .in(left_0_6_in),
    .out(left_0_6_out),
    .reset(left_0_6_reset),
    .write_en(left_0_6_write_en)
);
mac_pe pe_0_7 (
    .clk(pe_0_7_clk),
    .done(pe_0_7_done),
    .go(pe_0_7_go),
    .left(pe_0_7_left),
    .mul_ready(pe_0_7_mul_ready),
    .out(pe_0_7_out),
    .reset(pe_0_7_reset),
    .top(pe_0_7_top)
);
std_reg # (
    .WIDTH(32)
) top_0_7 (
    .clk(top_0_7_clk),
    .done(top_0_7_done),
    .in(top_0_7_in),
    .out(top_0_7_out),
    .reset(top_0_7_reset),
    .write_en(top_0_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_7 (
    .clk(left_0_7_clk),
    .done(left_0_7_done),
    .in(left_0_7_in),
    .out(left_0_7_out),
    .reset(left_0_7_reset),
    .write_en(left_0_7_write_en)
);
mac_pe pe_0_8 (
    .clk(pe_0_8_clk),
    .done(pe_0_8_done),
    .go(pe_0_8_go),
    .left(pe_0_8_left),
    .mul_ready(pe_0_8_mul_ready),
    .out(pe_0_8_out),
    .reset(pe_0_8_reset),
    .top(pe_0_8_top)
);
std_reg # (
    .WIDTH(32)
) top_0_8 (
    .clk(top_0_8_clk),
    .done(top_0_8_done),
    .in(top_0_8_in),
    .out(top_0_8_out),
    .reset(top_0_8_reset),
    .write_en(top_0_8_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_8 (
    .clk(left_0_8_clk),
    .done(left_0_8_done),
    .in(left_0_8_in),
    .out(left_0_8_out),
    .reset(left_0_8_reset),
    .write_en(left_0_8_write_en)
);
mac_pe pe_0_9 (
    .clk(pe_0_9_clk),
    .done(pe_0_9_done),
    .go(pe_0_9_go),
    .left(pe_0_9_left),
    .mul_ready(pe_0_9_mul_ready),
    .out(pe_0_9_out),
    .reset(pe_0_9_reset),
    .top(pe_0_9_top)
);
std_reg # (
    .WIDTH(32)
) top_0_9 (
    .clk(top_0_9_clk),
    .done(top_0_9_done),
    .in(top_0_9_in),
    .out(top_0_9_out),
    .reset(top_0_9_reset),
    .write_en(top_0_9_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_9 (
    .clk(left_0_9_clk),
    .done(left_0_9_done),
    .in(left_0_9_in),
    .out(left_0_9_out),
    .reset(left_0_9_reset),
    .write_en(left_0_9_write_en)
);
mac_pe pe_0_10 (
    .clk(pe_0_10_clk),
    .done(pe_0_10_done),
    .go(pe_0_10_go),
    .left(pe_0_10_left),
    .mul_ready(pe_0_10_mul_ready),
    .out(pe_0_10_out),
    .reset(pe_0_10_reset),
    .top(pe_0_10_top)
);
std_reg # (
    .WIDTH(32)
) top_0_10 (
    .clk(top_0_10_clk),
    .done(top_0_10_done),
    .in(top_0_10_in),
    .out(top_0_10_out),
    .reset(top_0_10_reset),
    .write_en(top_0_10_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_10 (
    .clk(left_0_10_clk),
    .done(left_0_10_done),
    .in(left_0_10_in),
    .out(left_0_10_out),
    .reset(left_0_10_reset),
    .write_en(left_0_10_write_en)
);
mac_pe pe_0_11 (
    .clk(pe_0_11_clk),
    .done(pe_0_11_done),
    .go(pe_0_11_go),
    .left(pe_0_11_left),
    .mul_ready(pe_0_11_mul_ready),
    .out(pe_0_11_out),
    .reset(pe_0_11_reset),
    .top(pe_0_11_top)
);
std_reg # (
    .WIDTH(32)
) top_0_11 (
    .clk(top_0_11_clk),
    .done(top_0_11_done),
    .in(top_0_11_in),
    .out(top_0_11_out),
    .reset(top_0_11_reset),
    .write_en(top_0_11_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_11 (
    .clk(left_0_11_clk),
    .done(left_0_11_done),
    .in(left_0_11_in),
    .out(left_0_11_out),
    .reset(left_0_11_reset),
    .write_en(left_0_11_write_en)
);
mac_pe pe_0_12 (
    .clk(pe_0_12_clk),
    .done(pe_0_12_done),
    .go(pe_0_12_go),
    .left(pe_0_12_left),
    .mul_ready(pe_0_12_mul_ready),
    .out(pe_0_12_out),
    .reset(pe_0_12_reset),
    .top(pe_0_12_top)
);
std_reg # (
    .WIDTH(32)
) top_0_12 (
    .clk(top_0_12_clk),
    .done(top_0_12_done),
    .in(top_0_12_in),
    .out(top_0_12_out),
    .reset(top_0_12_reset),
    .write_en(top_0_12_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_12 (
    .clk(left_0_12_clk),
    .done(left_0_12_done),
    .in(left_0_12_in),
    .out(left_0_12_out),
    .reset(left_0_12_reset),
    .write_en(left_0_12_write_en)
);
mac_pe pe_0_13 (
    .clk(pe_0_13_clk),
    .done(pe_0_13_done),
    .go(pe_0_13_go),
    .left(pe_0_13_left),
    .mul_ready(pe_0_13_mul_ready),
    .out(pe_0_13_out),
    .reset(pe_0_13_reset),
    .top(pe_0_13_top)
);
std_reg # (
    .WIDTH(32)
) top_0_13 (
    .clk(top_0_13_clk),
    .done(top_0_13_done),
    .in(top_0_13_in),
    .out(top_0_13_out),
    .reset(top_0_13_reset),
    .write_en(top_0_13_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_13 (
    .clk(left_0_13_clk),
    .done(left_0_13_done),
    .in(left_0_13_in),
    .out(left_0_13_out),
    .reset(left_0_13_reset),
    .write_en(left_0_13_write_en)
);
mac_pe pe_0_14 (
    .clk(pe_0_14_clk),
    .done(pe_0_14_done),
    .go(pe_0_14_go),
    .left(pe_0_14_left),
    .mul_ready(pe_0_14_mul_ready),
    .out(pe_0_14_out),
    .reset(pe_0_14_reset),
    .top(pe_0_14_top)
);
std_reg # (
    .WIDTH(32)
) top_0_14 (
    .clk(top_0_14_clk),
    .done(top_0_14_done),
    .in(top_0_14_in),
    .out(top_0_14_out),
    .reset(top_0_14_reset),
    .write_en(top_0_14_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_14 (
    .clk(left_0_14_clk),
    .done(left_0_14_done),
    .in(left_0_14_in),
    .out(left_0_14_out),
    .reset(left_0_14_reset),
    .write_en(left_0_14_write_en)
);
mac_pe pe_0_15 (
    .clk(pe_0_15_clk),
    .done(pe_0_15_done),
    .go(pe_0_15_go),
    .left(pe_0_15_left),
    .mul_ready(pe_0_15_mul_ready),
    .out(pe_0_15_out),
    .reset(pe_0_15_reset),
    .top(pe_0_15_top)
);
std_reg # (
    .WIDTH(32)
) top_0_15 (
    .clk(top_0_15_clk),
    .done(top_0_15_done),
    .in(top_0_15_in),
    .out(top_0_15_out),
    .reset(top_0_15_reset),
    .write_en(top_0_15_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_15 (
    .clk(left_0_15_clk),
    .done(left_0_15_done),
    .in(left_0_15_in),
    .out(left_0_15_out),
    .reset(left_0_15_reset),
    .write_en(left_0_15_write_en)
);
mac_pe pe_1_0 (
    .clk(pe_1_0_clk),
    .done(pe_1_0_done),
    .go(pe_1_0_go),
    .left(pe_1_0_left),
    .mul_ready(pe_1_0_mul_ready),
    .out(pe_1_0_out),
    .reset(pe_1_0_reset),
    .top(pe_1_0_top)
);
std_reg # (
    .WIDTH(32)
) top_1_0 (
    .clk(top_1_0_clk),
    .done(top_1_0_done),
    .in(top_1_0_in),
    .out(top_1_0_out),
    .reset(top_1_0_reset),
    .write_en(top_1_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_0 (
    .clk(left_1_0_clk),
    .done(left_1_0_done),
    .in(left_1_0_in),
    .out(left_1_0_out),
    .reset(left_1_0_reset),
    .write_en(left_1_0_write_en)
);
mac_pe pe_1_1 (
    .clk(pe_1_1_clk),
    .done(pe_1_1_done),
    .go(pe_1_1_go),
    .left(pe_1_1_left),
    .mul_ready(pe_1_1_mul_ready),
    .out(pe_1_1_out),
    .reset(pe_1_1_reset),
    .top(pe_1_1_top)
);
std_reg # (
    .WIDTH(32)
) top_1_1 (
    .clk(top_1_1_clk),
    .done(top_1_1_done),
    .in(top_1_1_in),
    .out(top_1_1_out),
    .reset(top_1_1_reset),
    .write_en(top_1_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_1 (
    .clk(left_1_1_clk),
    .done(left_1_1_done),
    .in(left_1_1_in),
    .out(left_1_1_out),
    .reset(left_1_1_reset),
    .write_en(left_1_1_write_en)
);
mac_pe pe_1_2 (
    .clk(pe_1_2_clk),
    .done(pe_1_2_done),
    .go(pe_1_2_go),
    .left(pe_1_2_left),
    .mul_ready(pe_1_2_mul_ready),
    .out(pe_1_2_out),
    .reset(pe_1_2_reset),
    .top(pe_1_2_top)
);
std_reg # (
    .WIDTH(32)
) top_1_2 (
    .clk(top_1_2_clk),
    .done(top_1_2_done),
    .in(top_1_2_in),
    .out(top_1_2_out),
    .reset(top_1_2_reset),
    .write_en(top_1_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_2 (
    .clk(left_1_2_clk),
    .done(left_1_2_done),
    .in(left_1_2_in),
    .out(left_1_2_out),
    .reset(left_1_2_reset),
    .write_en(left_1_2_write_en)
);
mac_pe pe_1_3 (
    .clk(pe_1_3_clk),
    .done(pe_1_3_done),
    .go(pe_1_3_go),
    .left(pe_1_3_left),
    .mul_ready(pe_1_3_mul_ready),
    .out(pe_1_3_out),
    .reset(pe_1_3_reset),
    .top(pe_1_3_top)
);
std_reg # (
    .WIDTH(32)
) top_1_3 (
    .clk(top_1_3_clk),
    .done(top_1_3_done),
    .in(top_1_3_in),
    .out(top_1_3_out),
    .reset(top_1_3_reset),
    .write_en(top_1_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_3 (
    .clk(left_1_3_clk),
    .done(left_1_3_done),
    .in(left_1_3_in),
    .out(left_1_3_out),
    .reset(left_1_3_reset),
    .write_en(left_1_3_write_en)
);
mac_pe pe_1_4 (
    .clk(pe_1_4_clk),
    .done(pe_1_4_done),
    .go(pe_1_4_go),
    .left(pe_1_4_left),
    .mul_ready(pe_1_4_mul_ready),
    .out(pe_1_4_out),
    .reset(pe_1_4_reset),
    .top(pe_1_4_top)
);
std_reg # (
    .WIDTH(32)
) top_1_4 (
    .clk(top_1_4_clk),
    .done(top_1_4_done),
    .in(top_1_4_in),
    .out(top_1_4_out),
    .reset(top_1_4_reset),
    .write_en(top_1_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_4 (
    .clk(left_1_4_clk),
    .done(left_1_4_done),
    .in(left_1_4_in),
    .out(left_1_4_out),
    .reset(left_1_4_reset),
    .write_en(left_1_4_write_en)
);
mac_pe pe_1_5 (
    .clk(pe_1_5_clk),
    .done(pe_1_5_done),
    .go(pe_1_5_go),
    .left(pe_1_5_left),
    .mul_ready(pe_1_5_mul_ready),
    .out(pe_1_5_out),
    .reset(pe_1_5_reset),
    .top(pe_1_5_top)
);
std_reg # (
    .WIDTH(32)
) top_1_5 (
    .clk(top_1_5_clk),
    .done(top_1_5_done),
    .in(top_1_5_in),
    .out(top_1_5_out),
    .reset(top_1_5_reset),
    .write_en(top_1_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_5 (
    .clk(left_1_5_clk),
    .done(left_1_5_done),
    .in(left_1_5_in),
    .out(left_1_5_out),
    .reset(left_1_5_reset),
    .write_en(left_1_5_write_en)
);
mac_pe pe_1_6 (
    .clk(pe_1_6_clk),
    .done(pe_1_6_done),
    .go(pe_1_6_go),
    .left(pe_1_6_left),
    .mul_ready(pe_1_6_mul_ready),
    .out(pe_1_6_out),
    .reset(pe_1_6_reset),
    .top(pe_1_6_top)
);
std_reg # (
    .WIDTH(32)
) top_1_6 (
    .clk(top_1_6_clk),
    .done(top_1_6_done),
    .in(top_1_6_in),
    .out(top_1_6_out),
    .reset(top_1_6_reset),
    .write_en(top_1_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_6 (
    .clk(left_1_6_clk),
    .done(left_1_6_done),
    .in(left_1_6_in),
    .out(left_1_6_out),
    .reset(left_1_6_reset),
    .write_en(left_1_6_write_en)
);
mac_pe pe_1_7 (
    .clk(pe_1_7_clk),
    .done(pe_1_7_done),
    .go(pe_1_7_go),
    .left(pe_1_7_left),
    .mul_ready(pe_1_7_mul_ready),
    .out(pe_1_7_out),
    .reset(pe_1_7_reset),
    .top(pe_1_7_top)
);
std_reg # (
    .WIDTH(32)
) top_1_7 (
    .clk(top_1_7_clk),
    .done(top_1_7_done),
    .in(top_1_7_in),
    .out(top_1_7_out),
    .reset(top_1_7_reset),
    .write_en(top_1_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_7 (
    .clk(left_1_7_clk),
    .done(left_1_7_done),
    .in(left_1_7_in),
    .out(left_1_7_out),
    .reset(left_1_7_reset),
    .write_en(left_1_7_write_en)
);
mac_pe pe_1_8 (
    .clk(pe_1_8_clk),
    .done(pe_1_8_done),
    .go(pe_1_8_go),
    .left(pe_1_8_left),
    .mul_ready(pe_1_8_mul_ready),
    .out(pe_1_8_out),
    .reset(pe_1_8_reset),
    .top(pe_1_8_top)
);
std_reg # (
    .WIDTH(32)
) top_1_8 (
    .clk(top_1_8_clk),
    .done(top_1_8_done),
    .in(top_1_8_in),
    .out(top_1_8_out),
    .reset(top_1_8_reset),
    .write_en(top_1_8_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_8 (
    .clk(left_1_8_clk),
    .done(left_1_8_done),
    .in(left_1_8_in),
    .out(left_1_8_out),
    .reset(left_1_8_reset),
    .write_en(left_1_8_write_en)
);
mac_pe pe_1_9 (
    .clk(pe_1_9_clk),
    .done(pe_1_9_done),
    .go(pe_1_9_go),
    .left(pe_1_9_left),
    .mul_ready(pe_1_9_mul_ready),
    .out(pe_1_9_out),
    .reset(pe_1_9_reset),
    .top(pe_1_9_top)
);
std_reg # (
    .WIDTH(32)
) top_1_9 (
    .clk(top_1_9_clk),
    .done(top_1_9_done),
    .in(top_1_9_in),
    .out(top_1_9_out),
    .reset(top_1_9_reset),
    .write_en(top_1_9_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_9 (
    .clk(left_1_9_clk),
    .done(left_1_9_done),
    .in(left_1_9_in),
    .out(left_1_9_out),
    .reset(left_1_9_reset),
    .write_en(left_1_9_write_en)
);
mac_pe pe_1_10 (
    .clk(pe_1_10_clk),
    .done(pe_1_10_done),
    .go(pe_1_10_go),
    .left(pe_1_10_left),
    .mul_ready(pe_1_10_mul_ready),
    .out(pe_1_10_out),
    .reset(pe_1_10_reset),
    .top(pe_1_10_top)
);
std_reg # (
    .WIDTH(32)
) top_1_10 (
    .clk(top_1_10_clk),
    .done(top_1_10_done),
    .in(top_1_10_in),
    .out(top_1_10_out),
    .reset(top_1_10_reset),
    .write_en(top_1_10_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_10 (
    .clk(left_1_10_clk),
    .done(left_1_10_done),
    .in(left_1_10_in),
    .out(left_1_10_out),
    .reset(left_1_10_reset),
    .write_en(left_1_10_write_en)
);
mac_pe pe_1_11 (
    .clk(pe_1_11_clk),
    .done(pe_1_11_done),
    .go(pe_1_11_go),
    .left(pe_1_11_left),
    .mul_ready(pe_1_11_mul_ready),
    .out(pe_1_11_out),
    .reset(pe_1_11_reset),
    .top(pe_1_11_top)
);
std_reg # (
    .WIDTH(32)
) top_1_11 (
    .clk(top_1_11_clk),
    .done(top_1_11_done),
    .in(top_1_11_in),
    .out(top_1_11_out),
    .reset(top_1_11_reset),
    .write_en(top_1_11_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_11 (
    .clk(left_1_11_clk),
    .done(left_1_11_done),
    .in(left_1_11_in),
    .out(left_1_11_out),
    .reset(left_1_11_reset),
    .write_en(left_1_11_write_en)
);
mac_pe pe_1_12 (
    .clk(pe_1_12_clk),
    .done(pe_1_12_done),
    .go(pe_1_12_go),
    .left(pe_1_12_left),
    .mul_ready(pe_1_12_mul_ready),
    .out(pe_1_12_out),
    .reset(pe_1_12_reset),
    .top(pe_1_12_top)
);
std_reg # (
    .WIDTH(32)
) top_1_12 (
    .clk(top_1_12_clk),
    .done(top_1_12_done),
    .in(top_1_12_in),
    .out(top_1_12_out),
    .reset(top_1_12_reset),
    .write_en(top_1_12_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_12 (
    .clk(left_1_12_clk),
    .done(left_1_12_done),
    .in(left_1_12_in),
    .out(left_1_12_out),
    .reset(left_1_12_reset),
    .write_en(left_1_12_write_en)
);
mac_pe pe_1_13 (
    .clk(pe_1_13_clk),
    .done(pe_1_13_done),
    .go(pe_1_13_go),
    .left(pe_1_13_left),
    .mul_ready(pe_1_13_mul_ready),
    .out(pe_1_13_out),
    .reset(pe_1_13_reset),
    .top(pe_1_13_top)
);
std_reg # (
    .WIDTH(32)
) top_1_13 (
    .clk(top_1_13_clk),
    .done(top_1_13_done),
    .in(top_1_13_in),
    .out(top_1_13_out),
    .reset(top_1_13_reset),
    .write_en(top_1_13_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_13 (
    .clk(left_1_13_clk),
    .done(left_1_13_done),
    .in(left_1_13_in),
    .out(left_1_13_out),
    .reset(left_1_13_reset),
    .write_en(left_1_13_write_en)
);
mac_pe pe_1_14 (
    .clk(pe_1_14_clk),
    .done(pe_1_14_done),
    .go(pe_1_14_go),
    .left(pe_1_14_left),
    .mul_ready(pe_1_14_mul_ready),
    .out(pe_1_14_out),
    .reset(pe_1_14_reset),
    .top(pe_1_14_top)
);
std_reg # (
    .WIDTH(32)
) top_1_14 (
    .clk(top_1_14_clk),
    .done(top_1_14_done),
    .in(top_1_14_in),
    .out(top_1_14_out),
    .reset(top_1_14_reset),
    .write_en(top_1_14_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_14 (
    .clk(left_1_14_clk),
    .done(left_1_14_done),
    .in(left_1_14_in),
    .out(left_1_14_out),
    .reset(left_1_14_reset),
    .write_en(left_1_14_write_en)
);
mac_pe pe_1_15 (
    .clk(pe_1_15_clk),
    .done(pe_1_15_done),
    .go(pe_1_15_go),
    .left(pe_1_15_left),
    .mul_ready(pe_1_15_mul_ready),
    .out(pe_1_15_out),
    .reset(pe_1_15_reset),
    .top(pe_1_15_top)
);
std_reg # (
    .WIDTH(32)
) top_1_15 (
    .clk(top_1_15_clk),
    .done(top_1_15_done),
    .in(top_1_15_in),
    .out(top_1_15_out),
    .reset(top_1_15_reset),
    .write_en(top_1_15_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_15 (
    .clk(left_1_15_clk),
    .done(left_1_15_done),
    .in(left_1_15_in),
    .out(left_1_15_out),
    .reset(left_1_15_reset),
    .write_en(left_1_15_write_en)
);
mac_pe pe_2_0 (
    .clk(pe_2_0_clk),
    .done(pe_2_0_done),
    .go(pe_2_0_go),
    .left(pe_2_0_left),
    .mul_ready(pe_2_0_mul_ready),
    .out(pe_2_0_out),
    .reset(pe_2_0_reset),
    .top(pe_2_0_top)
);
std_reg # (
    .WIDTH(32)
) top_2_0 (
    .clk(top_2_0_clk),
    .done(top_2_0_done),
    .in(top_2_0_in),
    .out(top_2_0_out),
    .reset(top_2_0_reset),
    .write_en(top_2_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_0 (
    .clk(left_2_0_clk),
    .done(left_2_0_done),
    .in(left_2_0_in),
    .out(left_2_0_out),
    .reset(left_2_0_reset),
    .write_en(left_2_0_write_en)
);
mac_pe pe_2_1 (
    .clk(pe_2_1_clk),
    .done(pe_2_1_done),
    .go(pe_2_1_go),
    .left(pe_2_1_left),
    .mul_ready(pe_2_1_mul_ready),
    .out(pe_2_1_out),
    .reset(pe_2_1_reset),
    .top(pe_2_1_top)
);
std_reg # (
    .WIDTH(32)
) top_2_1 (
    .clk(top_2_1_clk),
    .done(top_2_1_done),
    .in(top_2_1_in),
    .out(top_2_1_out),
    .reset(top_2_1_reset),
    .write_en(top_2_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_1 (
    .clk(left_2_1_clk),
    .done(left_2_1_done),
    .in(left_2_1_in),
    .out(left_2_1_out),
    .reset(left_2_1_reset),
    .write_en(left_2_1_write_en)
);
mac_pe pe_2_2 (
    .clk(pe_2_2_clk),
    .done(pe_2_2_done),
    .go(pe_2_2_go),
    .left(pe_2_2_left),
    .mul_ready(pe_2_2_mul_ready),
    .out(pe_2_2_out),
    .reset(pe_2_2_reset),
    .top(pe_2_2_top)
);
std_reg # (
    .WIDTH(32)
) top_2_2 (
    .clk(top_2_2_clk),
    .done(top_2_2_done),
    .in(top_2_2_in),
    .out(top_2_2_out),
    .reset(top_2_2_reset),
    .write_en(top_2_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_2 (
    .clk(left_2_2_clk),
    .done(left_2_2_done),
    .in(left_2_2_in),
    .out(left_2_2_out),
    .reset(left_2_2_reset),
    .write_en(left_2_2_write_en)
);
mac_pe pe_2_3 (
    .clk(pe_2_3_clk),
    .done(pe_2_3_done),
    .go(pe_2_3_go),
    .left(pe_2_3_left),
    .mul_ready(pe_2_3_mul_ready),
    .out(pe_2_3_out),
    .reset(pe_2_3_reset),
    .top(pe_2_3_top)
);
std_reg # (
    .WIDTH(32)
) top_2_3 (
    .clk(top_2_3_clk),
    .done(top_2_3_done),
    .in(top_2_3_in),
    .out(top_2_3_out),
    .reset(top_2_3_reset),
    .write_en(top_2_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_3 (
    .clk(left_2_3_clk),
    .done(left_2_3_done),
    .in(left_2_3_in),
    .out(left_2_3_out),
    .reset(left_2_3_reset),
    .write_en(left_2_3_write_en)
);
mac_pe pe_2_4 (
    .clk(pe_2_4_clk),
    .done(pe_2_4_done),
    .go(pe_2_4_go),
    .left(pe_2_4_left),
    .mul_ready(pe_2_4_mul_ready),
    .out(pe_2_4_out),
    .reset(pe_2_4_reset),
    .top(pe_2_4_top)
);
std_reg # (
    .WIDTH(32)
) top_2_4 (
    .clk(top_2_4_clk),
    .done(top_2_4_done),
    .in(top_2_4_in),
    .out(top_2_4_out),
    .reset(top_2_4_reset),
    .write_en(top_2_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_4 (
    .clk(left_2_4_clk),
    .done(left_2_4_done),
    .in(left_2_4_in),
    .out(left_2_4_out),
    .reset(left_2_4_reset),
    .write_en(left_2_4_write_en)
);
mac_pe pe_2_5 (
    .clk(pe_2_5_clk),
    .done(pe_2_5_done),
    .go(pe_2_5_go),
    .left(pe_2_5_left),
    .mul_ready(pe_2_5_mul_ready),
    .out(pe_2_5_out),
    .reset(pe_2_5_reset),
    .top(pe_2_5_top)
);
std_reg # (
    .WIDTH(32)
) top_2_5 (
    .clk(top_2_5_clk),
    .done(top_2_5_done),
    .in(top_2_5_in),
    .out(top_2_5_out),
    .reset(top_2_5_reset),
    .write_en(top_2_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_5 (
    .clk(left_2_5_clk),
    .done(left_2_5_done),
    .in(left_2_5_in),
    .out(left_2_5_out),
    .reset(left_2_5_reset),
    .write_en(left_2_5_write_en)
);
mac_pe pe_2_6 (
    .clk(pe_2_6_clk),
    .done(pe_2_6_done),
    .go(pe_2_6_go),
    .left(pe_2_6_left),
    .mul_ready(pe_2_6_mul_ready),
    .out(pe_2_6_out),
    .reset(pe_2_6_reset),
    .top(pe_2_6_top)
);
std_reg # (
    .WIDTH(32)
) top_2_6 (
    .clk(top_2_6_clk),
    .done(top_2_6_done),
    .in(top_2_6_in),
    .out(top_2_6_out),
    .reset(top_2_6_reset),
    .write_en(top_2_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_6 (
    .clk(left_2_6_clk),
    .done(left_2_6_done),
    .in(left_2_6_in),
    .out(left_2_6_out),
    .reset(left_2_6_reset),
    .write_en(left_2_6_write_en)
);
mac_pe pe_2_7 (
    .clk(pe_2_7_clk),
    .done(pe_2_7_done),
    .go(pe_2_7_go),
    .left(pe_2_7_left),
    .mul_ready(pe_2_7_mul_ready),
    .out(pe_2_7_out),
    .reset(pe_2_7_reset),
    .top(pe_2_7_top)
);
std_reg # (
    .WIDTH(32)
) top_2_7 (
    .clk(top_2_7_clk),
    .done(top_2_7_done),
    .in(top_2_7_in),
    .out(top_2_7_out),
    .reset(top_2_7_reset),
    .write_en(top_2_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_7 (
    .clk(left_2_7_clk),
    .done(left_2_7_done),
    .in(left_2_7_in),
    .out(left_2_7_out),
    .reset(left_2_7_reset),
    .write_en(left_2_7_write_en)
);
mac_pe pe_2_8 (
    .clk(pe_2_8_clk),
    .done(pe_2_8_done),
    .go(pe_2_8_go),
    .left(pe_2_8_left),
    .mul_ready(pe_2_8_mul_ready),
    .out(pe_2_8_out),
    .reset(pe_2_8_reset),
    .top(pe_2_8_top)
);
std_reg # (
    .WIDTH(32)
) top_2_8 (
    .clk(top_2_8_clk),
    .done(top_2_8_done),
    .in(top_2_8_in),
    .out(top_2_8_out),
    .reset(top_2_8_reset),
    .write_en(top_2_8_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_8 (
    .clk(left_2_8_clk),
    .done(left_2_8_done),
    .in(left_2_8_in),
    .out(left_2_8_out),
    .reset(left_2_8_reset),
    .write_en(left_2_8_write_en)
);
mac_pe pe_2_9 (
    .clk(pe_2_9_clk),
    .done(pe_2_9_done),
    .go(pe_2_9_go),
    .left(pe_2_9_left),
    .mul_ready(pe_2_9_mul_ready),
    .out(pe_2_9_out),
    .reset(pe_2_9_reset),
    .top(pe_2_9_top)
);
std_reg # (
    .WIDTH(32)
) top_2_9 (
    .clk(top_2_9_clk),
    .done(top_2_9_done),
    .in(top_2_9_in),
    .out(top_2_9_out),
    .reset(top_2_9_reset),
    .write_en(top_2_9_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_9 (
    .clk(left_2_9_clk),
    .done(left_2_9_done),
    .in(left_2_9_in),
    .out(left_2_9_out),
    .reset(left_2_9_reset),
    .write_en(left_2_9_write_en)
);
mac_pe pe_2_10 (
    .clk(pe_2_10_clk),
    .done(pe_2_10_done),
    .go(pe_2_10_go),
    .left(pe_2_10_left),
    .mul_ready(pe_2_10_mul_ready),
    .out(pe_2_10_out),
    .reset(pe_2_10_reset),
    .top(pe_2_10_top)
);
std_reg # (
    .WIDTH(32)
) top_2_10 (
    .clk(top_2_10_clk),
    .done(top_2_10_done),
    .in(top_2_10_in),
    .out(top_2_10_out),
    .reset(top_2_10_reset),
    .write_en(top_2_10_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_10 (
    .clk(left_2_10_clk),
    .done(left_2_10_done),
    .in(left_2_10_in),
    .out(left_2_10_out),
    .reset(left_2_10_reset),
    .write_en(left_2_10_write_en)
);
mac_pe pe_2_11 (
    .clk(pe_2_11_clk),
    .done(pe_2_11_done),
    .go(pe_2_11_go),
    .left(pe_2_11_left),
    .mul_ready(pe_2_11_mul_ready),
    .out(pe_2_11_out),
    .reset(pe_2_11_reset),
    .top(pe_2_11_top)
);
std_reg # (
    .WIDTH(32)
) top_2_11 (
    .clk(top_2_11_clk),
    .done(top_2_11_done),
    .in(top_2_11_in),
    .out(top_2_11_out),
    .reset(top_2_11_reset),
    .write_en(top_2_11_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_11 (
    .clk(left_2_11_clk),
    .done(left_2_11_done),
    .in(left_2_11_in),
    .out(left_2_11_out),
    .reset(left_2_11_reset),
    .write_en(left_2_11_write_en)
);
mac_pe pe_2_12 (
    .clk(pe_2_12_clk),
    .done(pe_2_12_done),
    .go(pe_2_12_go),
    .left(pe_2_12_left),
    .mul_ready(pe_2_12_mul_ready),
    .out(pe_2_12_out),
    .reset(pe_2_12_reset),
    .top(pe_2_12_top)
);
std_reg # (
    .WIDTH(32)
) top_2_12 (
    .clk(top_2_12_clk),
    .done(top_2_12_done),
    .in(top_2_12_in),
    .out(top_2_12_out),
    .reset(top_2_12_reset),
    .write_en(top_2_12_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_12 (
    .clk(left_2_12_clk),
    .done(left_2_12_done),
    .in(left_2_12_in),
    .out(left_2_12_out),
    .reset(left_2_12_reset),
    .write_en(left_2_12_write_en)
);
mac_pe pe_2_13 (
    .clk(pe_2_13_clk),
    .done(pe_2_13_done),
    .go(pe_2_13_go),
    .left(pe_2_13_left),
    .mul_ready(pe_2_13_mul_ready),
    .out(pe_2_13_out),
    .reset(pe_2_13_reset),
    .top(pe_2_13_top)
);
std_reg # (
    .WIDTH(32)
) top_2_13 (
    .clk(top_2_13_clk),
    .done(top_2_13_done),
    .in(top_2_13_in),
    .out(top_2_13_out),
    .reset(top_2_13_reset),
    .write_en(top_2_13_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_13 (
    .clk(left_2_13_clk),
    .done(left_2_13_done),
    .in(left_2_13_in),
    .out(left_2_13_out),
    .reset(left_2_13_reset),
    .write_en(left_2_13_write_en)
);
mac_pe pe_2_14 (
    .clk(pe_2_14_clk),
    .done(pe_2_14_done),
    .go(pe_2_14_go),
    .left(pe_2_14_left),
    .mul_ready(pe_2_14_mul_ready),
    .out(pe_2_14_out),
    .reset(pe_2_14_reset),
    .top(pe_2_14_top)
);
std_reg # (
    .WIDTH(32)
) top_2_14 (
    .clk(top_2_14_clk),
    .done(top_2_14_done),
    .in(top_2_14_in),
    .out(top_2_14_out),
    .reset(top_2_14_reset),
    .write_en(top_2_14_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_14 (
    .clk(left_2_14_clk),
    .done(left_2_14_done),
    .in(left_2_14_in),
    .out(left_2_14_out),
    .reset(left_2_14_reset),
    .write_en(left_2_14_write_en)
);
mac_pe pe_2_15 (
    .clk(pe_2_15_clk),
    .done(pe_2_15_done),
    .go(pe_2_15_go),
    .left(pe_2_15_left),
    .mul_ready(pe_2_15_mul_ready),
    .out(pe_2_15_out),
    .reset(pe_2_15_reset),
    .top(pe_2_15_top)
);
std_reg # (
    .WIDTH(32)
) top_2_15 (
    .clk(top_2_15_clk),
    .done(top_2_15_done),
    .in(top_2_15_in),
    .out(top_2_15_out),
    .reset(top_2_15_reset),
    .write_en(top_2_15_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_15 (
    .clk(left_2_15_clk),
    .done(left_2_15_done),
    .in(left_2_15_in),
    .out(left_2_15_out),
    .reset(left_2_15_reset),
    .write_en(left_2_15_write_en)
);
mac_pe pe_3_0 (
    .clk(pe_3_0_clk),
    .done(pe_3_0_done),
    .go(pe_3_0_go),
    .left(pe_3_0_left),
    .mul_ready(pe_3_0_mul_ready),
    .out(pe_3_0_out),
    .reset(pe_3_0_reset),
    .top(pe_3_0_top)
);
std_reg # (
    .WIDTH(32)
) top_3_0 (
    .clk(top_3_0_clk),
    .done(top_3_0_done),
    .in(top_3_0_in),
    .out(top_3_0_out),
    .reset(top_3_0_reset),
    .write_en(top_3_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_0 (
    .clk(left_3_0_clk),
    .done(left_3_0_done),
    .in(left_3_0_in),
    .out(left_3_0_out),
    .reset(left_3_0_reset),
    .write_en(left_3_0_write_en)
);
mac_pe pe_3_1 (
    .clk(pe_3_1_clk),
    .done(pe_3_1_done),
    .go(pe_3_1_go),
    .left(pe_3_1_left),
    .mul_ready(pe_3_1_mul_ready),
    .out(pe_3_1_out),
    .reset(pe_3_1_reset),
    .top(pe_3_1_top)
);
std_reg # (
    .WIDTH(32)
) top_3_1 (
    .clk(top_3_1_clk),
    .done(top_3_1_done),
    .in(top_3_1_in),
    .out(top_3_1_out),
    .reset(top_3_1_reset),
    .write_en(top_3_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_1 (
    .clk(left_3_1_clk),
    .done(left_3_1_done),
    .in(left_3_1_in),
    .out(left_3_1_out),
    .reset(left_3_1_reset),
    .write_en(left_3_1_write_en)
);
mac_pe pe_3_2 (
    .clk(pe_3_2_clk),
    .done(pe_3_2_done),
    .go(pe_3_2_go),
    .left(pe_3_2_left),
    .mul_ready(pe_3_2_mul_ready),
    .out(pe_3_2_out),
    .reset(pe_3_2_reset),
    .top(pe_3_2_top)
);
std_reg # (
    .WIDTH(32)
) top_3_2 (
    .clk(top_3_2_clk),
    .done(top_3_2_done),
    .in(top_3_2_in),
    .out(top_3_2_out),
    .reset(top_3_2_reset),
    .write_en(top_3_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_2 (
    .clk(left_3_2_clk),
    .done(left_3_2_done),
    .in(left_3_2_in),
    .out(left_3_2_out),
    .reset(left_3_2_reset),
    .write_en(left_3_2_write_en)
);
mac_pe pe_3_3 (
    .clk(pe_3_3_clk),
    .done(pe_3_3_done),
    .go(pe_3_3_go),
    .left(pe_3_3_left),
    .mul_ready(pe_3_3_mul_ready),
    .out(pe_3_3_out),
    .reset(pe_3_3_reset),
    .top(pe_3_3_top)
);
std_reg # (
    .WIDTH(32)
) top_3_3 (
    .clk(top_3_3_clk),
    .done(top_3_3_done),
    .in(top_3_3_in),
    .out(top_3_3_out),
    .reset(top_3_3_reset),
    .write_en(top_3_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_3 (
    .clk(left_3_3_clk),
    .done(left_3_3_done),
    .in(left_3_3_in),
    .out(left_3_3_out),
    .reset(left_3_3_reset),
    .write_en(left_3_3_write_en)
);
mac_pe pe_3_4 (
    .clk(pe_3_4_clk),
    .done(pe_3_4_done),
    .go(pe_3_4_go),
    .left(pe_3_4_left),
    .mul_ready(pe_3_4_mul_ready),
    .out(pe_3_4_out),
    .reset(pe_3_4_reset),
    .top(pe_3_4_top)
);
std_reg # (
    .WIDTH(32)
) top_3_4 (
    .clk(top_3_4_clk),
    .done(top_3_4_done),
    .in(top_3_4_in),
    .out(top_3_4_out),
    .reset(top_3_4_reset),
    .write_en(top_3_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_4 (
    .clk(left_3_4_clk),
    .done(left_3_4_done),
    .in(left_3_4_in),
    .out(left_3_4_out),
    .reset(left_3_4_reset),
    .write_en(left_3_4_write_en)
);
mac_pe pe_3_5 (
    .clk(pe_3_5_clk),
    .done(pe_3_5_done),
    .go(pe_3_5_go),
    .left(pe_3_5_left),
    .mul_ready(pe_3_5_mul_ready),
    .out(pe_3_5_out),
    .reset(pe_3_5_reset),
    .top(pe_3_5_top)
);
std_reg # (
    .WIDTH(32)
) top_3_5 (
    .clk(top_3_5_clk),
    .done(top_3_5_done),
    .in(top_3_5_in),
    .out(top_3_5_out),
    .reset(top_3_5_reset),
    .write_en(top_3_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_5 (
    .clk(left_3_5_clk),
    .done(left_3_5_done),
    .in(left_3_5_in),
    .out(left_3_5_out),
    .reset(left_3_5_reset),
    .write_en(left_3_5_write_en)
);
mac_pe pe_3_6 (
    .clk(pe_3_6_clk),
    .done(pe_3_6_done),
    .go(pe_3_6_go),
    .left(pe_3_6_left),
    .mul_ready(pe_3_6_mul_ready),
    .out(pe_3_6_out),
    .reset(pe_3_6_reset),
    .top(pe_3_6_top)
);
std_reg # (
    .WIDTH(32)
) top_3_6 (
    .clk(top_3_6_clk),
    .done(top_3_6_done),
    .in(top_3_6_in),
    .out(top_3_6_out),
    .reset(top_3_6_reset),
    .write_en(top_3_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_6 (
    .clk(left_3_6_clk),
    .done(left_3_6_done),
    .in(left_3_6_in),
    .out(left_3_6_out),
    .reset(left_3_6_reset),
    .write_en(left_3_6_write_en)
);
mac_pe pe_3_7 (
    .clk(pe_3_7_clk),
    .done(pe_3_7_done),
    .go(pe_3_7_go),
    .left(pe_3_7_left),
    .mul_ready(pe_3_7_mul_ready),
    .out(pe_3_7_out),
    .reset(pe_3_7_reset),
    .top(pe_3_7_top)
);
std_reg # (
    .WIDTH(32)
) top_3_7 (
    .clk(top_3_7_clk),
    .done(top_3_7_done),
    .in(top_3_7_in),
    .out(top_3_7_out),
    .reset(top_3_7_reset),
    .write_en(top_3_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_7 (
    .clk(left_3_7_clk),
    .done(left_3_7_done),
    .in(left_3_7_in),
    .out(left_3_7_out),
    .reset(left_3_7_reset),
    .write_en(left_3_7_write_en)
);
mac_pe pe_3_8 (
    .clk(pe_3_8_clk),
    .done(pe_3_8_done),
    .go(pe_3_8_go),
    .left(pe_3_8_left),
    .mul_ready(pe_3_8_mul_ready),
    .out(pe_3_8_out),
    .reset(pe_3_8_reset),
    .top(pe_3_8_top)
);
std_reg # (
    .WIDTH(32)
) top_3_8 (
    .clk(top_3_8_clk),
    .done(top_3_8_done),
    .in(top_3_8_in),
    .out(top_3_8_out),
    .reset(top_3_8_reset),
    .write_en(top_3_8_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_8 (
    .clk(left_3_8_clk),
    .done(left_3_8_done),
    .in(left_3_8_in),
    .out(left_3_8_out),
    .reset(left_3_8_reset),
    .write_en(left_3_8_write_en)
);
mac_pe pe_3_9 (
    .clk(pe_3_9_clk),
    .done(pe_3_9_done),
    .go(pe_3_9_go),
    .left(pe_3_9_left),
    .mul_ready(pe_3_9_mul_ready),
    .out(pe_3_9_out),
    .reset(pe_3_9_reset),
    .top(pe_3_9_top)
);
std_reg # (
    .WIDTH(32)
) top_3_9 (
    .clk(top_3_9_clk),
    .done(top_3_9_done),
    .in(top_3_9_in),
    .out(top_3_9_out),
    .reset(top_3_9_reset),
    .write_en(top_3_9_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_9 (
    .clk(left_3_9_clk),
    .done(left_3_9_done),
    .in(left_3_9_in),
    .out(left_3_9_out),
    .reset(left_3_9_reset),
    .write_en(left_3_9_write_en)
);
mac_pe pe_3_10 (
    .clk(pe_3_10_clk),
    .done(pe_3_10_done),
    .go(pe_3_10_go),
    .left(pe_3_10_left),
    .mul_ready(pe_3_10_mul_ready),
    .out(pe_3_10_out),
    .reset(pe_3_10_reset),
    .top(pe_3_10_top)
);
std_reg # (
    .WIDTH(32)
) top_3_10 (
    .clk(top_3_10_clk),
    .done(top_3_10_done),
    .in(top_3_10_in),
    .out(top_3_10_out),
    .reset(top_3_10_reset),
    .write_en(top_3_10_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_10 (
    .clk(left_3_10_clk),
    .done(left_3_10_done),
    .in(left_3_10_in),
    .out(left_3_10_out),
    .reset(left_3_10_reset),
    .write_en(left_3_10_write_en)
);
mac_pe pe_3_11 (
    .clk(pe_3_11_clk),
    .done(pe_3_11_done),
    .go(pe_3_11_go),
    .left(pe_3_11_left),
    .mul_ready(pe_3_11_mul_ready),
    .out(pe_3_11_out),
    .reset(pe_3_11_reset),
    .top(pe_3_11_top)
);
std_reg # (
    .WIDTH(32)
) top_3_11 (
    .clk(top_3_11_clk),
    .done(top_3_11_done),
    .in(top_3_11_in),
    .out(top_3_11_out),
    .reset(top_3_11_reset),
    .write_en(top_3_11_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_11 (
    .clk(left_3_11_clk),
    .done(left_3_11_done),
    .in(left_3_11_in),
    .out(left_3_11_out),
    .reset(left_3_11_reset),
    .write_en(left_3_11_write_en)
);
mac_pe pe_3_12 (
    .clk(pe_3_12_clk),
    .done(pe_3_12_done),
    .go(pe_3_12_go),
    .left(pe_3_12_left),
    .mul_ready(pe_3_12_mul_ready),
    .out(pe_3_12_out),
    .reset(pe_3_12_reset),
    .top(pe_3_12_top)
);
std_reg # (
    .WIDTH(32)
) top_3_12 (
    .clk(top_3_12_clk),
    .done(top_3_12_done),
    .in(top_3_12_in),
    .out(top_3_12_out),
    .reset(top_3_12_reset),
    .write_en(top_3_12_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_12 (
    .clk(left_3_12_clk),
    .done(left_3_12_done),
    .in(left_3_12_in),
    .out(left_3_12_out),
    .reset(left_3_12_reset),
    .write_en(left_3_12_write_en)
);
mac_pe pe_3_13 (
    .clk(pe_3_13_clk),
    .done(pe_3_13_done),
    .go(pe_3_13_go),
    .left(pe_3_13_left),
    .mul_ready(pe_3_13_mul_ready),
    .out(pe_3_13_out),
    .reset(pe_3_13_reset),
    .top(pe_3_13_top)
);
std_reg # (
    .WIDTH(32)
) top_3_13 (
    .clk(top_3_13_clk),
    .done(top_3_13_done),
    .in(top_3_13_in),
    .out(top_3_13_out),
    .reset(top_3_13_reset),
    .write_en(top_3_13_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_13 (
    .clk(left_3_13_clk),
    .done(left_3_13_done),
    .in(left_3_13_in),
    .out(left_3_13_out),
    .reset(left_3_13_reset),
    .write_en(left_3_13_write_en)
);
mac_pe pe_3_14 (
    .clk(pe_3_14_clk),
    .done(pe_3_14_done),
    .go(pe_3_14_go),
    .left(pe_3_14_left),
    .mul_ready(pe_3_14_mul_ready),
    .out(pe_3_14_out),
    .reset(pe_3_14_reset),
    .top(pe_3_14_top)
);
std_reg # (
    .WIDTH(32)
) top_3_14 (
    .clk(top_3_14_clk),
    .done(top_3_14_done),
    .in(top_3_14_in),
    .out(top_3_14_out),
    .reset(top_3_14_reset),
    .write_en(top_3_14_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_14 (
    .clk(left_3_14_clk),
    .done(left_3_14_done),
    .in(left_3_14_in),
    .out(left_3_14_out),
    .reset(left_3_14_reset),
    .write_en(left_3_14_write_en)
);
mac_pe pe_3_15 (
    .clk(pe_3_15_clk),
    .done(pe_3_15_done),
    .go(pe_3_15_go),
    .left(pe_3_15_left),
    .mul_ready(pe_3_15_mul_ready),
    .out(pe_3_15_out),
    .reset(pe_3_15_reset),
    .top(pe_3_15_top)
);
std_reg # (
    .WIDTH(32)
) top_3_15 (
    .clk(top_3_15_clk),
    .done(top_3_15_done),
    .in(top_3_15_in),
    .out(top_3_15_out),
    .reset(top_3_15_reset),
    .write_en(top_3_15_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_15 (
    .clk(left_3_15_clk),
    .done(left_3_15_done),
    .in(left_3_15_in),
    .out(left_3_15_out),
    .reset(left_3_15_reset),
    .write_en(left_3_15_write_en)
);
mac_pe pe_4_0 (
    .clk(pe_4_0_clk),
    .done(pe_4_0_done),
    .go(pe_4_0_go),
    .left(pe_4_0_left),
    .mul_ready(pe_4_0_mul_ready),
    .out(pe_4_0_out),
    .reset(pe_4_0_reset),
    .top(pe_4_0_top)
);
std_reg # (
    .WIDTH(32)
) top_4_0 (
    .clk(top_4_0_clk),
    .done(top_4_0_done),
    .in(top_4_0_in),
    .out(top_4_0_out),
    .reset(top_4_0_reset),
    .write_en(top_4_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_0 (
    .clk(left_4_0_clk),
    .done(left_4_0_done),
    .in(left_4_0_in),
    .out(left_4_0_out),
    .reset(left_4_0_reset),
    .write_en(left_4_0_write_en)
);
mac_pe pe_4_1 (
    .clk(pe_4_1_clk),
    .done(pe_4_1_done),
    .go(pe_4_1_go),
    .left(pe_4_1_left),
    .mul_ready(pe_4_1_mul_ready),
    .out(pe_4_1_out),
    .reset(pe_4_1_reset),
    .top(pe_4_1_top)
);
std_reg # (
    .WIDTH(32)
) top_4_1 (
    .clk(top_4_1_clk),
    .done(top_4_1_done),
    .in(top_4_1_in),
    .out(top_4_1_out),
    .reset(top_4_1_reset),
    .write_en(top_4_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_1 (
    .clk(left_4_1_clk),
    .done(left_4_1_done),
    .in(left_4_1_in),
    .out(left_4_1_out),
    .reset(left_4_1_reset),
    .write_en(left_4_1_write_en)
);
mac_pe pe_4_2 (
    .clk(pe_4_2_clk),
    .done(pe_4_2_done),
    .go(pe_4_2_go),
    .left(pe_4_2_left),
    .mul_ready(pe_4_2_mul_ready),
    .out(pe_4_2_out),
    .reset(pe_4_2_reset),
    .top(pe_4_2_top)
);
std_reg # (
    .WIDTH(32)
) top_4_2 (
    .clk(top_4_2_clk),
    .done(top_4_2_done),
    .in(top_4_2_in),
    .out(top_4_2_out),
    .reset(top_4_2_reset),
    .write_en(top_4_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_2 (
    .clk(left_4_2_clk),
    .done(left_4_2_done),
    .in(left_4_2_in),
    .out(left_4_2_out),
    .reset(left_4_2_reset),
    .write_en(left_4_2_write_en)
);
mac_pe pe_4_3 (
    .clk(pe_4_3_clk),
    .done(pe_4_3_done),
    .go(pe_4_3_go),
    .left(pe_4_3_left),
    .mul_ready(pe_4_3_mul_ready),
    .out(pe_4_3_out),
    .reset(pe_4_3_reset),
    .top(pe_4_3_top)
);
std_reg # (
    .WIDTH(32)
) top_4_3 (
    .clk(top_4_3_clk),
    .done(top_4_3_done),
    .in(top_4_3_in),
    .out(top_4_3_out),
    .reset(top_4_3_reset),
    .write_en(top_4_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_3 (
    .clk(left_4_3_clk),
    .done(left_4_3_done),
    .in(left_4_3_in),
    .out(left_4_3_out),
    .reset(left_4_3_reset),
    .write_en(left_4_3_write_en)
);
mac_pe pe_4_4 (
    .clk(pe_4_4_clk),
    .done(pe_4_4_done),
    .go(pe_4_4_go),
    .left(pe_4_4_left),
    .mul_ready(pe_4_4_mul_ready),
    .out(pe_4_4_out),
    .reset(pe_4_4_reset),
    .top(pe_4_4_top)
);
std_reg # (
    .WIDTH(32)
) top_4_4 (
    .clk(top_4_4_clk),
    .done(top_4_4_done),
    .in(top_4_4_in),
    .out(top_4_4_out),
    .reset(top_4_4_reset),
    .write_en(top_4_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_4 (
    .clk(left_4_4_clk),
    .done(left_4_4_done),
    .in(left_4_4_in),
    .out(left_4_4_out),
    .reset(left_4_4_reset),
    .write_en(left_4_4_write_en)
);
mac_pe pe_4_5 (
    .clk(pe_4_5_clk),
    .done(pe_4_5_done),
    .go(pe_4_5_go),
    .left(pe_4_5_left),
    .mul_ready(pe_4_5_mul_ready),
    .out(pe_4_5_out),
    .reset(pe_4_5_reset),
    .top(pe_4_5_top)
);
std_reg # (
    .WIDTH(32)
) top_4_5 (
    .clk(top_4_5_clk),
    .done(top_4_5_done),
    .in(top_4_5_in),
    .out(top_4_5_out),
    .reset(top_4_5_reset),
    .write_en(top_4_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_5 (
    .clk(left_4_5_clk),
    .done(left_4_5_done),
    .in(left_4_5_in),
    .out(left_4_5_out),
    .reset(left_4_5_reset),
    .write_en(left_4_5_write_en)
);
mac_pe pe_4_6 (
    .clk(pe_4_6_clk),
    .done(pe_4_6_done),
    .go(pe_4_6_go),
    .left(pe_4_6_left),
    .mul_ready(pe_4_6_mul_ready),
    .out(pe_4_6_out),
    .reset(pe_4_6_reset),
    .top(pe_4_6_top)
);
std_reg # (
    .WIDTH(32)
) top_4_6 (
    .clk(top_4_6_clk),
    .done(top_4_6_done),
    .in(top_4_6_in),
    .out(top_4_6_out),
    .reset(top_4_6_reset),
    .write_en(top_4_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_6 (
    .clk(left_4_6_clk),
    .done(left_4_6_done),
    .in(left_4_6_in),
    .out(left_4_6_out),
    .reset(left_4_6_reset),
    .write_en(left_4_6_write_en)
);
mac_pe pe_4_7 (
    .clk(pe_4_7_clk),
    .done(pe_4_7_done),
    .go(pe_4_7_go),
    .left(pe_4_7_left),
    .mul_ready(pe_4_7_mul_ready),
    .out(pe_4_7_out),
    .reset(pe_4_7_reset),
    .top(pe_4_7_top)
);
std_reg # (
    .WIDTH(32)
) top_4_7 (
    .clk(top_4_7_clk),
    .done(top_4_7_done),
    .in(top_4_7_in),
    .out(top_4_7_out),
    .reset(top_4_7_reset),
    .write_en(top_4_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_7 (
    .clk(left_4_7_clk),
    .done(left_4_7_done),
    .in(left_4_7_in),
    .out(left_4_7_out),
    .reset(left_4_7_reset),
    .write_en(left_4_7_write_en)
);
mac_pe pe_4_8 (
    .clk(pe_4_8_clk),
    .done(pe_4_8_done),
    .go(pe_4_8_go),
    .left(pe_4_8_left),
    .mul_ready(pe_4_8_mul_ready),
    .out(pe_4_8_out),
    .reset(pe_4_8_reset),
    .top(pe_4_8_top)
);
std_reg # (
    .WIDTH(32)
) top_4_8 (
    .clk(top_4_8_clk),
    .done(top_4_8_done),
    .in(top_4_8_in),
    .out(top_4_8_out),
    .reset(top_4_8_reset),
    .write_en(top_4_8_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_8 (
    .clk(left_4_8_clk),
    .done(left_4_8_done),
    .in(left_4_8_in),
    .out(left_4_8_out),
    .reset(left_4_8_reset),
    .write_en(left_4_8_write_en)
);
mac_pe pe_4_9 (
    .clk(pe_4_9_clk),
    .done(pe_4_9_done),
    .go(pe_4_9_go),
    .left(pe_4_9_left),
    .mul_ready(pe_4_9_mul_ready),
    .out(pe_4_9_out),
    .reset(pe_4_9_reset),
    .top(pe_4_9_top)
);
std_reg # (
    .WIDTH(32)
) top_4_9 (
    .clk(top_4_9_clk),
    .done(top_4_9_done),
    .in(top_4_9_in),
    .out(top_4_9_out),
    .reset(top_4_9_reset),
    .write_en(top_4_9_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_9 (
    .clk(left_4_9_clk),
    .done(left_4_9_done),
    .in(left_4_9_in),
    .out(left_4_9_out),
    .reset(left_4_9_reset),
    .write_en(left_4_9_write_en)
);
mac_pe pe_4_10 (
    .clk(pe_4_10_clk),
    .done(pe_4_10_done),
    .go(pe_4_10_go),
    .left(pe_4_10_left),
    .mul_ready(pe_4_10_mul_ready),
    .out(pe_4_10_out),
    .reset(pe_4_10_reset),
    .top(pe_4_10_top)
);
std_reg # (
    .WIDTH(32)
) top_4_10 (
    .clk(top_4_10_clk),
    .done(top_4_10_done),
    .in(top_4_10_in),
    .out(top_4_10_out),
    .reset(top_4_10_reset),
    .write_en(top_4_10_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_10 (
    .clk(left_4_10_clk),
    .done(left_4_10_done),
    .in(left_4_10_in),
    .out(left_4_10_out),
    .reset(left_4_10_reset),
    .write_en(left_4_10_write_en)
);
mac_pe pe_4_11 (
    .clk(pe_4_11_clk),
    .done(pe_4_11_done),
    .go(pe_4_11_go),
    .left(pe_4_11_left),
    .mul_ready(pe_4_11_mul_ready),
    .out(pe_4_11_out),
    .reset(pe_4_11_reset),
    .top(pe_4_11_top)
);
std_reg # (
    .WIDTH(32)
) top_4_11 (
    .clk(top_4_11_clk),
    .done(top_4_11_done),
    .in(top_4_11_in),
    .out(top_4_11_out),
    .reset(top_4_11_reset),
    .write_en(top_4_11_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_11 (
    .clk(left_4_11_clk),
    .done(left_4_11_done),
    .in(left_4_11_in),
    .out(left_4_11_out),
    .reset(left_4_11_reset),
    .write_en(left_4_11_write_en)
);
mac_pe pe_4_12 (
    .clk(pe_4_12_clk),
    .done(pe_4_12_done),
    .go(pe_4_12_go),
    .left(pe_4_12_left),
    .mul_ready(pe_4_12_mul_ready),
    .out(pe_4_12_out),
    .reset(pe_4_12_reset),
    .top(pe_4_12_top)
);
std_reg # (
    .WIDTH(32)
) top_4_12 (
    .clk(top_4_12_clk),
    .done(top_4_12_done),
    .in(top_4_12_in),
    .out(top_4_12_out),
    .reset(top_4_12_reset),
    .write_en(top_4_12_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_12 (
    .clk(left_4_12_clk),
    .done(left_4_12_done),
    .in(left_4_12_in),
    .out(left_4_12_out),
    .reset(left_4_12_reset),
    .write_en(left_4_12_write_en)
);
mac_pe pe_4_13 (
    .clk(pe_4_13_clk),
    .done(pe_4_13_done),
    .go(pe_4_13_go),
    .left(pe_4_13_left),
    .mul_ready(pe_4_13_mul_ready),
    .out(pe_4_13_out),
    .reset(pe_4_13_reset),
    .top(pe_4_13_top)
);
std_reg # (
    .WIDTH(32)
) top_4_13 (
    .clk(top_4_13_clk),
    .done(top_4_13_done),
    .in(top_4_13_in),
    .out(top_4_13_out),
    .reset(top_4_13_reset),
    .write_en(top_4_13_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_13 (
    .clk(left_4_13_clk),
    .done(left_4_13_done),
    .in(left_4_13_in),
    .out(left_4_13_out),
    .reset(left_4_13_reset),
    .write_en(left_4_13_write_en)
);
mac_pe pe_4_14 (
    .clk(pe_4_14_clk),
    .done(pe_4_14_done),
    .go(pe_4_14_go),
    .left(pe_4_14_left),
    .mul_ready(pe_4_14_mul_ready),
    .out(pe_4_14_out),
    .reset(pe_4_14_reset),
    .top(pe_4_14_top)
);
std_reg # (
    .WIDTH(32)
) top_4_14 (
    .clk(top_4_14_clk),
    .done(top_4_14_done),
    .in(top_4_14_in),
    .out(top_4_14_out),
    .reset(top_4_14_reset),
    .write_en(top_4_14_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_14 (
    .clk(left_4_14_clk),
    .done(left_4_14_done),
    .in(left_4_14_in),
    .out(left_4_14_out),
    .reset(left_4_14_reset),
    .write_en(left_4_14_write_en)
);
mac_pe pe_4_15 (
    .clk(pe_4_15_clk),
    .done(pe_4_15_done),
    .go(pe_4_15_go),
    .left(pe_4_15_left),
    .mul_ready(pe_4_15_mul_ready),
    .out(pe_4_15_out),
    .reset(pe_4_15_reset),
    .top(pe_4_15_top)
);
std_reg # (
    .WIDTH(32)
) top_4_15 (
    .clk(top_4_15_clk),
    .done(top_4_15_done),
    .in(top_4_15_in),
    .out(top_4_15_out),
    .reset(top_4_15_reset),
    .write_en(top_4_15_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_15 (
    .clk(left_4_15_clk),
    .done(left_4_15_done),
    .in(left_4_15_in),
    .out(left_4_15_out),
    .reset(left_4_15_reset),
    .write_en(left_4_15_write_en)
);
mac_pe pe_5_0 (
    .clk(pe_5_0_clk),
    .done(pe_5_0_done),
    .go(pe_5_0_go),
    .left(pe_5_0_left),
    .mul_ready(pe_5_0_mul_ready),
    .out(pe_5_0_out),
    .reset(pe_5_0_reset),
    .top(pe_5_0_top)
);
std_reg # (
    .WIDTH(32)
) top_5_0 (
    .clk(top_5_0_clk),
    .done(top_5_0_done),
    .in(top_5_0_in),
    .out(top_5_0_out),
    .reset(top_5_0_reset),
    .write_en(top_5_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_0 (
    .clk(left_5_0_clk),
    .done(left_5_0_done),
    .in(left_5_0_in),
    .out(left_5_0_out),
    .reset(left_5_0_reset),
    .write_en(left_5_0_write_en)
);
mac_pe pe_5_1 (
    .clk(pe_5_1_clk),
    .done(pe_5_1_done),
    .go(pe_5_1_go),
    .left(pe_5_1_left),
    .mul_ready(pe_5_1_mul_ready),
    .out(pe_5_1_out),
    .reset(pe_5_1_reset),
    .top(pe_5_1_top)
);
std_reg # (
    .WIDTH(32)
) top_5_1 (
    .clk(top_5_1_clk),
    .done(top_5_1_done),
    .in(top_5_1_in),
    .out(top_5_1_out),
    .reset(top_5_1_reset),
    .write_en(top_5_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_1 (
    .clk(left_5_1_clk),
    .done(left_5_1_done),
    .in(left_5_1_in),
    .out(left_5_1_out),
    .reset(left_5_1_reset),
    .write_en(left_5_1_write_en)
);
mac_pe pe_5_2 (
    .clk(pe_5_2_clk),
    .done(pe_5_2_done),
    .go(pe_5_2_go),
    .left(pe_5_2_left),
    .mul_ready(pe_5_2_mul_ready),
    .out(pe_5_2_out),
    .reset(pe_5_2_reset),
    .top(pe_5_2_top)
);
std_reg # (
    .WIDTH(32)
) top_5_2 (
    .clk(top_5_2_clk),
    .done(top_5_2_done),
    .in(top_5_2_in),
    .out(top_5_2_out),
    .reset(top_5_2_reset),
    .write_en(top_5_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_2 (
    .clk(left_5_2_clk),
    .done(left_5_2_done),
    .in(left_5_2_in),
    .out(left_5_2_out),
    .reset(left_5_2_reset),
    .write_en(left_5_2_write_en)
);
mac_pe pe_5_3 (
    .clk(pe_5_3_clk),
    .done(pe_5_3_done),
    .go(pe_5_3_go),
    .left(pe_5_3_left),
    .mul_ready(pe_5_3_mul_ready),
    .out(pe_5_3_out),
    .reset(pe_5_3_reset),
    .top(pe_5_3_top)
);
std_reg # (
    .WIDTH(32)
) top_5_3 (
    .clk(top_5_3_clk),
    .done(top_5_3_done),
    .in(top_5_3_in),
    .out(top_5_3_out),
    .reset(top_5_3_reset),
    .write_en(top_5_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_3 (
    .clk(left_5_3_clk),
    .done(left_5_3_done),
    .in(left_5_3_in),
    .out(left_5_3_out),
    .reset(left_5_3_reset),
    .write_en(left_5_3_write_en)
);
mac_pe pe_5_4 (
    .clk(pe_5_4_clk),
    .done(pe_5_4_done),
    .go(pe_5_4_go),
    .left(pe_5_4_left),
    .mul_ready(pe_5_4_mul_ready),
    .out(pe_5_4_out),
    .reset(pe_5_4_reset),
    .top(pe_5_4_top)
);
std_reg # (
    .WIDTH(32)
) top_5_4 (
    .clk(top_5_4_clk),
    .done(top_5_4_done),
    .in(top_5_4_in),
    .out(top_5_4_out),
    .reset(top_5_4_reset),
    .write_en(top_5_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_4 (
    .clk(left_5_4_clk),
    .done(left_5_4_done),
    .in(left_5_4_in),
    .out(left_5_4_out),
    .reset(left_5_4_reset),
    .write_en(left_5_4_write_en)
);
mac_pe pe_5_5 (
    .clk(pe_5_5_clk),
    .done(pe_5_5_done),
    .go(pe_5_5_go),
    .left(pe_5_5_left),
    .mul_ready(pe_5_5_mul_ready),
    .out(pe_5_5_out),
    .reset(pe_5_5_reset),
    .top(pe_5_5_top)
);
std_reg # (
    .WIDTH(32)
) top_5_5 (
    .clk(top_5_5_clk),
    .done(top_5_5_done),
    .in(top_5_5_in),
    .out(top_5_5_out),
    .reset(top_5_5_reset),
    .write_en(top_5_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_5 (
    .clk(left_5_5_clk),
    .done(left_5_5_done),
    .in(left_5_5_in),
    .out(left_5_5_out),
    .reset(left_5_5_reset),
    .write_en(left_5_5_write_en)
);
mac_pe pe_5_6 (
    .clk(pe_5_6_clk),
    .done(pe_5_6_done),
    .go(pe_5_6_go),
    .left(pe_5_6_left),
    .mul_ready(pe_5_6_mul_ready),
    .out(pe_5_6_out),
    .reset(pe_5_6_reset),
    .top(pe_5_6_top)
);
std_reg # (
    .WIDTH(32)
) top_5_6 (
    .clk(top_5_6_clk),
    .done(top_5_6_done),
    .in(top_5_6_in),
    .out(top_5_6_out),
    .reset(top_5_6_reset),
    .write_en(top_5_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_6 (
    .clk(left_5_6_clk),
    .done(left_5_6_done),
    .in(left_5_6_in),
    .out(left_5_6_out),
    .reset(left_5_6_reset),
    .write_en(left_5_6_write_en)
);
mac_pe pe_5_7 (
    .clk(pe_5_7_clk),
    .done(pe_5_7_done),
    .go(pe_5_7_go),
    .left(pe_5_7_left),
    .mul_ready(pe_5_7_mul_ready),
    .out(pe_5_7_out),
    .reset(pe_5_7_reset),
    .top(pe_5_7_top)
);
std_reg # (
    .WIDTH(32)
) top_5_7 (
    .clk(top_5_7_clk),
    .done(top_5_7_done),
    .in(top_5_7_in),
    .out(top_5_7_out),
    .reset(top_5_7_reset),
    .write_en(top_5_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_7 (
    .clk(left_5_7_clk),
    .done(left_5_7_done),
    .in(left_5_7_in),
    .out(left_5_7_out),
    .reset(left_5_7_reset),
    .write_en(left_5_7_write_en)
);
mac_pe pe_5_8 (
    .clk(pe_5_8_clk),
    .done(pe_5_8_done),
    .go(pe_5_8_go),
    .left(pe_5_8_left),
    .mul_ready(pe_5_8_mul_ready),
    .out(pe_5_8_out),
    .reset(pe_5_8_reset),
    .top(pe_5_8_top)
);
std_reg # (
    .WIDTH(32)
) top_5_8 (
    .clk(top_5_8_clk),
    .done(top_5_8_done),
    .in(top_5_8_in),
    .out(top_5_8_out),
    .reset(top_5_8_reset),
    .write_en(top_5_8_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_8 (
    .clk(left_5_8_clk),
    .done(left_5_8_done),
    .in(left_5_8_in),
    .out(left_5_8_out),
    .reset(left_5_8_reset),
    .write_en(left_5_8_write_en)
);
mac_pe pe_5_9 (
    .clk(pe_5_9_clk),
    .done(pe_5_9_done),
    .go(pe_5_9_go),
    .left(pe_5_9_left),
    .mul_ready(pe_5_9_mul_ready),
    .out(pe_5_9_out),
    .reset(pe_5_9_reset),
    .top(pe_5_9_top)
);
std_reg # (
    .WIDTH(32)
) top_5_9 (
    .clk(top_5_9_clk),
    .done(top_5_9_done),
    .in(top_5_9_in),
    .out(top_5_9_out),
    .reset(top_5_9_reset),
    .write_en(top_5_9_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_9 (
    .clk(left_5_9_clk),
    .done(left_5_9_done),
    .in(left_5_9_in),
    .out(left_5_9_out),
    .reset(left_5_9_reset),
    .write_en(left_5_9_write_en)
);
mac_pe pe_5_10 (
    .clk(pe_5_10_clk),
    .done(pe_5_10_done),
    .go(pe_5_10_go),
    .left(pe_5_10_left),
    .mul_ready(pe_5_10_mul_ready),
    .out(pe_5_10_out),
    .reset(pe_5_10_reset),
    .top(pe_5_10_top)
);
std_reg # (
    .WIDTH(32)
) top_5_10 (
    .clk(top_5_10_clk),
    .done(top_5_10_done),
    .in(top_5_10_in),
    .out(top_5_10_out),
    .reset(top_5_10_reset),
    .write_en(top_5_10_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_10 (
    .clk(left_5_10_clk),
    .done(left_5_10_done),
    .in(left_5_10_in),
    .out(left_5_10_out),
    .reset(left_5_10_reset),
    .write_en(left_5_10_write_en)
);
mac_pe pe_5_11 (
    .clk(pe_5_11_clk),
    .done(pe_5_11_done),
    .go(pe_5_11_go),
    .left(pe_5_11_left),
    .mul_ready(pe_5_11_mul_ready),
    .out(pe_5_11_out),
    .reset(pe_5_11_reset),
    .top(pe_5_11_top)
);
std_reg # (
    .WIDTH(32)
) top_5_11 (
    .clk(top_5_11_clk),
    .done(top_5_11_done),
    .in(top_5_11_in),
    .out(top_5_11_out),
    .reset(top_5_11_reset),
    .write_en(top_5_11_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_11 (
    .clk(left_5_11_clk),
    .done(left_5_11_done),
    .in(left_5_11_in),
    .out(left_5_11_out),
    .reset(left_5_11_reset),
    .write_en(left_5_11_write_en)
);
mac_pe pe_5_12 (
    .clk(pe_5_12_clk),
    .done(pe_5_12_done),
    .go(pe_5_12_go),
    .left(pe_5_12_left),
    .mul_ready(pe_5_12_mul_ready),
    .out(pe_5_12_out),
    .reset(pe_5_12_reset),
    .top(pe_5_12_top)
);
std_reg # (
    .WIDTH(32)
) top_5_12 (
    .clk(top_5_12_clk),
    .done(top_5_12_done),
    .in(top_5_12_in),
    .out(top_5_12_out),
    .reset(top_5_12_reset),
    .write_en(top_5_12_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_12 (
    .clk(left_5_12_clk),
    .done(left_5_12_done),
    .in(left_5_12_in),
    .out(left_5_12_out),
    .reset(left_5_12_reset),
    .write_en(left_5_12_write_en)
);
mac_pe pe_5_13 (
    .clk(pe_5_13_clk),
    .done(pe_5_13_done),
    .go(pe_5_13_go),
    .left(pe_5_13_left),
    .mul_ready(pe_5_13_mul_ready),
    .out(pe_5_13_out),
    .reset(pe_5_13_reset),
    .top(pe_5_13_top)
);
std_reg # (
    .WIDTH(32)
) top_5_13 (
    .clk(top_5_13_clk),
    .done(top_5_13_done),
    .in(top_5_13_in),
    .out(top_5_13_out),
    .reset(top_5_13_reset),
    .write_en(top_5_13_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_13 (
    .clk(left_5_13_clk),
    .done(left_5_13_done),
    .in(left_5_13_in),
    .out(left_5_13_out),
    .reset(left_5_13_reset),
    .write_en(left_5_13_write_en)
);
mac_pe pe_5_14 (
    .clk(pe_5_14_clk),
    .done(pe_5_14_done),
    .go(pe_5_14_go),
    .left(pe_5_14_left),
    .mul_ready(pe_5_14_mul_ready),
    .out(pe_5_14_out),
    .reset(pe_5_14_reset),
    .top(pe_5_14_top)
);
std_reg # (
    .WIDTH(32)
) top_5_14 (
    .clk(top_5_14_clk),
    .done(top_5_14_done),
    .in(top_5_14_in),
    .out(top_5_14_out),
    .reset(top_5_14_reset),
    .write_en(top_5_14_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_14 (
    .clk(left_5_14_clk),
    .done(left_5_14_done),
    .in(left_5_14_in),
    .out(left_5_14_out),
    .reset(left_5_14_reset),
    .write_en(left_5_14_write_en)
);
mac_pe pe_5_15 (
    .clk(pe_5_15_clk),
    .done(pe_5_15_done),
    .go(pe_5_15_go),
    .left(pe_5_15_left),
    .mul_ready(pe_5_15_mul_ready),
    .out(pe_5_15_out),
    .reset(pe_5_15_reset),
    .top(pe_5_15_top)
);
std_reg # (
    .WIDTH(32)
) top_5_15 (
    .clk(top_5_15_clk),
    .done(top_5_15_done),
    .in(top_5_15_in),
    .out(top_5_15_out),
    .reset(top_5_15_reset),
    .write_en(top_5_15_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_15 (
    .clk(left_5_15_clk),
    .done(left_5_15_done),
    .in(left_5_15_in),
    .out(left_5_15_out),
    .reset(left_5_15_reset),
    .write_en(left_5_15_write_en)
);
mac_pe pe_6_0 (
    .clk(pe_6_0_clk),
    .done(pe_6_0_done),
    .go(pe_6_0_go),
    .left(pe_6_0_left),
    .mul_ready(pe_6_0_mul_ready),
    .out(pe_6_0_out),
    .reset(pe_6_0_reset),
    .top(pe_6_0_top)
);
std_reg # (
    .WIDTH(32)
) top_6_0 (
    .clk(top_6_0_clk),
    .done(top_6_0_done),
    .in(top_6_0_in),
    .out(top_6_0_out),
    .reset(top_6_0_reset),
    .write_en(top_6_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_0 (
    .clk(left_6_0_clk),
    .done(left_6_0_done),
    .in(left_6_0_in),
    .out(left_6_0_out),
    .reset(left_6_0_reset),
    .write_en(left_6_0_write_en)
);
mac_pe pe_6_1 (
    .clk(pe_6_1_clk),
    .done(pe_6_1_done),
    .go(pe_6_1_go),
    .left(pe_6_1_left),
    .mul_ready(pe_6_1_mul_ready),
    .out(pe_6_1_out),
    .reset(pe_6_1_reset),
    .top(pe_6_1_top)
);
std_reg # (
    .WIDTH(32)
) top_6_1 (
    .clk(top_6_1_clk),
    .done(top_6_1_done),
    .in(top_6_1_in),
    .out(top_6_1_out),
    .reset(top_6_1_reset),
    .write_en(top_6_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_1 (
    .clk(left_6_1_clk),
    .done(left_6_1_done),
    .in(left_6_1_in),
    .out(left_6_1_out),
    .reset(left_6_1_reset),
    .write_en(left_6_1_write_en)
);
mac_pe pe_6_2 (
    .clk(pe_6_2_clk),
    .done(pe_6_2_done),
    .go(pe_6_2_go),
    .left(pe_6_2_left),
    .mul_ready(pe_6_2_mul_ready),
    .out(pe_6_2_out),
    .reset(pe_6_2_reset),
    .top(pe_6_2_top)
);
std_reg # (
    .WIDTH(32)
) top_6_2 (
    .clk(top_6_2_clk),
    .done(top_6_2_done),
    .in(top_6_2_in),
    .out(top_6_2_out),
    .reset(top_6_2_reset),
    .write_en(top_6_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_2 (
    .clk(left_6_2_clk),
    .done(left_6_2_done),
    .in(left_6_2_in),
    .out(left_6_2_out),
    .reset(left_6_2_reset),
    .write_en(left_6_2_write_en)
);
mac_pe pe_6_3 (
    .clk(pe_6_3_clk),
    .done(pe_6_3_done),
    .go(pe_6_3_go),
    .left(pe_6_3_left),
    .mul_ready(pe_6_3_mul_ready),
    .out(pe_6_3_out),
    .reset(pe_6_3_reset),
    .top(pe_6_3_top)
);
std_reg # (
    .WIDTH(32)
) top_6_3 (
    .clk(top_6_3_clk),
    .done(top_6_3_done),
    .in(top_6_3_in),
    .out(top_6_3_out),
    .reset(top_6_3_reset),
    .write_en(top_6_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_3 (
    .clk(left_6_3_clk),
    .done(left_6_3_done),
    .in(left_6_3_in),
    .out(left_6_3_out),
    .reset(left_6_3_reset),
    .write_en(left_6_3_write_en)
);
mac_pe pe_6_4 (
    .clk(pe_6_4_clk),
    .done(pe_6_4_done),
    .go(pe_6_4_go),
    .left(pe_6_4_left),
    .mul_ready(pe_6_4_mul_ready),
    .out(pe_6_4_out),
    .reset(pe_6_4_reset),
    .top(pe_6_4_top)
);
std_reg # (
    .WIDTH(32)
) top_6_4 (
    .clk(top_6_4_clk),
    .done(top_6_4_done),
    .in(top_6_4_in),
    .out(top_6_4_out),
    .reset(top_6_4_reset),
    .write_en(top_6_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_4 (
    .clk(left_6_4_clk),
    .done(left_6_4_done),
    .in(left_6_4_in),
    .out(left_6_4_out),
    .reset(left_6_4_reset),
    .write_en(left_6_4_write_en)
);
mac_pe pe_6_5 (
    .clk(pe_6_5_clk),
    .done(pe_6_5_done),
    .go(pe_6_5_go),
    .left(pe_6_5_left),
    .mul_ready(pe_6_5_mul_ready),
    .out(pe_6_5_out),
    .reset(pe_6_5_reset),
    .top(pe_6_5_top)
);
std_reg # (
    .WIDTH(32)
) top_6_5 (
    .clk(top_6_5_clk),
    .done(top_6_5_done),
    .in(top_6_5_in),
    .out(top_6_5_out),
    .reset(top_6_5_reset),
    .write_en(top_6_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_5 (
    .clk(left_6_5_clk),
    .done(left_6_5_done),
    .in(left_6_5_in),
    .out(left_6_5_out),
    .reset(left_6_5_reset),
    .write_en(left_6_5_write_en)
);
mac_pe pe_6_6 (
    .clk(pe_6_6_clk),
    .done(pe_6_6_done),
    .go(pe_6_6_go),
    .left(pe_6_6_left),
    .mul_ready(pe_6_6_mul_ready),
    .out(pe_6_6_out),
    .reset(pe_6_6_reset),
    .top(pe_6_6_top)
);
std_reg # (
    .WIDTH(32)
) top_6_6 (
    .clk(top_6_6_clk),
    .done(top_6_6_done),
    .in(top_6_6_in),
    .out(top_6_6_out),
    .reset(top_6_6_reset),
    .write_en(top_6_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_6 (
    .clk(left_6_6_clk),
    .done(left_6_6_done),
    .in(left_6_6_in),
    .out(left_6_6_out),
    .reset(left_6_6_reset),
    .write_en(left_6_6_write_en)
);
mac_pe pe_6_7 (
    .clk(pe_6_7_clk),
    .done(pe_6_7_done),
    .go(pe_6_7_go),
    .left(pe_6_7_left),
    .mul_ready(pe_6_7_mul_ready),
    .out(pe_6_7_out),
    .reset(pe_6_7_reset),
    .top(pe_6_7_top)
);
std_reg # (
    .WIDTH(32)
) top_6_7 (
    .clk(top_6_7_clk),
    .done(top_6_7_done),
    .in(top_6_7_in),
    .out(top_6_7_out),
    .reset(top_6_7_reset),
    .write_en(top_6_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_7 (
    .clk(left_6_7_clk),
    .done(left_6_7_done),
    .in(left_6_7_in),
    .out(left_6_7_out),
    .reset(left_6_7_reset),
    .write_en(left_6_7_write_en)
);
mac_pe pe_6_8 (
    .clk(pe_6_8_clk),
    .done(pe_6_8_done),
    .go(pe_6_8_go),
    .left(pe_6_8_left),
    .mul_ready(pe_6_8_mul_ready),
    .out(pe_6_8_out),
    .reset(pe_6_8_reset),
    .top(pe_6_8_top)
);
std_reg # (
    .WIDTH(32)
) top_6_8 (
    .clk(top_6_8_clk),
    .done(top_6_8_done),
    .in(top_6_8_in),
    .out(top_6_8_out),
    .reset(top_6_8_reset),
    .write_en(top_6_8_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_8 (
    .clk(left_6_8_clk),
    .done(left_6_8_done),
    .in(left_6_8_in),
    .out(left_6_8_out),
    .reset(left_6_8_reset),
    .write_en(left_6_8_write_en)
);
mac_pe pe_6_9 (
    .clk(pe_6_9_clk),
    .done(pe_6_9_done),
    .go(pe_6_9_go),
    .left(pe_6_9_left),
    .mul_ready(pe_6_9_mul_ready),
    .out(pe_6_9_out),
    .reset(pe_6_9_reset),
    .top(pe_6_9_top)
);
std_reg # (
    .WIDTH(32)
) top_6_9 (
    .clk(top_6_9_clk),
    .done(top_6_9_done),
    .in(top_6_9_in),
    .out(top_6_9_out),
    .reset(top_6_9_reset),
    .write_en(top_6_9_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_9 (
    .clk(left_6_9_clk),
    .done(left_6_9_done),
    .in(left_6_9_in),
    .out(left_6_9_out),
    .reset(left_6_9_reset),
    .write_en(left_6_9_write_en)
);
mac_pe pe_6_10 (
    .clk(pe_6_10_clk),
    .done(pe_6_10_done),
    .go(pe_6_10_go),
    .left(pe_6_10_left),
    .mul_ready(pe_6_10_mul_ready),
    .out(pe_6_10_out),
    .reset(pe_6_10_reset),
    .top(pe_6_10_top)
);
std_reg # (
    .WIDTH(32)
) top_6_10 (
    .clk(top_6_10_clk),
    .done(top_6_10_done),
    .in(top_6_10_in),
    .out(top_6_10_out),
    .reset(top_6_10_reset),
    .write_en(top_6_10_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_10 (
    .clk(left_6_10_clk),
    .done(left_6_10_done),
    .in(left_6_10_in),
    .out(left_6_10_out),
    .reset(left_6_10_reset),
    .write_en(left_6_10_write_en)
);
mac_pe pe_6_11 (
    .clk(pe_6_11_clk),
    .done(pe_6_11_done),
    .go(pe_6_11_go),
    .left(pe_6_11_left),
    .mul_ready(pe_6_11_mul_ready),
    .out(pe_6_11_out),
    .reset(pe_6_11_reset),
    .top(pe_6_11_top)
);
std_reg # (
    .WIDTH(32)
) top_6_11 (
    .clk(top_6_11_clk),
    .done(top_6_11_done),
    .in(top_6_11_in),
    .out(top_6_11_out),
    .reset(top_6_11_reset),
    .write_en(top_6_11_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_11 (
    .clk(left_6_11_clk),
    .done(left_6_11_done),
    .in(left_6_11_in),
    .out(left_6_11_out),
    .reset(left_6_11_reset),
    .write_en(left_6_11_write_en)
);
mac_pe pe_6_12 (
    .clk(pe_6_12_clk),
    .done(pe_6_12_done),
    .go(pe_6_12_go),
    .left(pe_6_12_left),
    .mul_ready(pe_6_12_mul_ready),
    .out(pe_6_12_out),
    .reset(pe_6_12_reset),
    .top(pe_6_12_top)
);
std_reg # (
    .WIDTH(32)
) top_6_12 (
    .clk(top_6_12_clk),
    .done(top_6_12_done),
    .in(top_6_12_in),
    .out(top_6_12_out),
    .reset(top_6_12_reset),
    .write_en(top_6_12_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_12 (
    .clk(left_6_12_clk),
    .done(left_6_12_done),
    .in(left_6_12_in),
    .out(left_6_12_out),
    .reset(left_6_12_reset),
    .write_en(left_6_12_write_en)
);
mac_pe pe_6_13 (
    .clk(pe_6_13_clk),
    .done(pe_6_13_done),
    .go(pe_6_13_go),
    .left(pe_6_13_left),
    .mul_ready(pe_6_13_mul_ready),
    .out(pe_6_13_out),
    .reset(pe_6_13_reset),
    .top(pe_6_13_top)
);
std_reg # (
    .WIDTH(32)
) top_6_13 (
    .clk(top_6_13_clk),
    .done(top_6_13_done),
    .in(top_6_13_in),
    .out(top_6_13_out),
    .reset(top_6_13_reset),
    .write_en(top_6_13_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_13 (
    .clk(left_6_13_clk),
    .done(left_6_13_done),
    .in(left_6_13_in),
    .out(left_6_13_out),
    .reset(left_6_13_reset),
    .write_en(left_6_13_write_en)
);
mac_pe pe_6_14 (
    .clk(pe_6_14_clk),
    .done(pe_6_14_done),
    .go(pe_6_14_go),
    .left(pe_6_14_left),
    .mul_ready(pe_6_14_mul_ready),
    .out(pe_6_14_out),
    .reset(pe_6_14_reset),
    .top(pe_6_14_top)
);
std_reg # (
    .WIDTH(32)
) top_6_14 (
    .clk(top_6_14_clk),
    .done(top_6_14_done),
    .in(top_6_14_in),
    .out(top_6_14_out),
    .reset(top_6_14_reset),
    .write_en(top_6_14_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_14 (
    .clk(left_6_14_clk),
    .done(left_6_14_done),
    .in(left_6_14_in),
    .out(left_6_14_out),
    .reset(left_6_14_reset),
    .write_en(left_6_14_write_en)
);
mac_pe pe_6_15 (
    .clk(pe_6_15_clk),
    .done(pe_6_15_done),
    .go(pe_6_15_go),
    .left(pe_6_15_left),
    .mul_ready(pe_6_15_mul_ready),
    .out(pe_6_15_out),
    .reset(pe_6_15_reset),
    .top(pe_6_15_top)
);
std_reg # (
    .WIDTH(32)
) top_6_15 (
    .clk(top_6_15_clk),
    .done(top_6_15_done),
    .in(top_6_15_in),
    .out(top_6_15_out),
    .reset(top_6_15_reset),
    .write_en(top_6_15_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_15 (
    .clk(left_6_15_clk),
    .done(left_6_15_done),
    .in(left_6_15_in),
    .out(left_6_15_out),
    .reset(left_6_15_reset),
    .write_en(left_6_15_write_en)
);
mac_pe pe_7_0 (
    .clk(pe_7_0_clk),
    .done(pe_7_0_done),
    .go(pe_7_0_go),
    .left(pe_7_0_left),
    .mul_ready(pe_7_0_mul_ready),
    .out(pe_7_0_out),
    .reset(pe_7_0_reset),
    .top(pe_7_0_top)
);
std_reg # (
    .WIDTH(32)
) top_7_0 (
    .clk(top_7_0_clk),
    .done(top_7_0_done),
    .in(top_7_0_in),
    .out(top_7_0_out),
    .reset(top_7_0_reset),
    .write_en(top_7_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_0 (
    .clk(left_7_0_clk),
    .done(left_7_0_done),
    .in(left_7_0_in),
    .out(left_7_0_out),
    .reset(left_7_0_reset),
    .write_en(left_7_0_write_en)
);
mac_pe pe_7_1 (
    .clk(pe_7_1_clk),
    .done(pe_7_1_done),
    .go(pe_7_1_go),
    .left(pe_7_1_left),
    .mul_ready(pe_7_1_mul_ready),
    .out(pe_7_1_out),
    .reset(pe_7_1_reset),
    .top(pe_7_1_top)
);
std_reg # (
    .WIDTH(32)
) top_7_1 (
    .clk(top_7_1_clk),
    .done(top_7_1_done),
    .in(top_7_1_in),
    .out(top_7_1_out),
    .reset(top_7_1_reset),
    .write_en(top_7_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_1 (
    .clk(left_7_1_clk),
    .done(left_7_1_done),
    .in(left_7_1_in),
    .out(left_7_1_out),
    .reset(left_7_1_reset),
    .write_en(left_7_1_write_en)
);
mac_pe pe_7_2 (
    .clk(pe_7_2_clk),
    .done(pe_7_2_done),
    .go(pe_7_2_go),
    .left(pe_7_2_left),
    .mul_ready(pe_7_2_mul_ready),
    .out(pe_7_2_out),
    .reset(pe_7_2_reset),
    .top(pe_7_2_top)
);
std_reg # (
    .WIDTH(32)
) top_7_2 (
    .clk(top_7_2_clk),
    .done(top_7_2_done),
    .in(top_7_2_in),
    .out(top_7_2_out),
    .reset(top_7_2_reset),
    .write_en(top_7_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_2 (
    .clk(left_7_2_clk),
    .done(left_7_2_done),
    .in(left_7_2_in),
    .out(left_7_2_out),
    .reset(left_7_2_reset),
    .write_en(left_7_2_write_en)
);
mac_pe pe_7_3 (
    .clk(pe_7_3_clk),
    .done(pe_7_3_done),
    .go(pe_7_3_go),
    .left(pe_7_3_left),
    .mul_ready(pe_7_3_mul_ready),
    .out(pe_7_3_out),
    .reset(pe_7_3_reset),
    .top(pe_7_3_top)
);
std_reg # (
    .WIDTH(32)
) top_7_3 (
    .clk(top_7_3_clk),
    .done(top_7_3_done),
    .in(top_7_3_in),
    .out(top_7_3_out),
    .reset(top_7_3_reset),
    .write_en(top_7_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_3 (
    .clk(left_7_3_clk),
    .done(left_7_3_done),
    .in(left_7_3_in),
    .out(left_7_3_out),
    .reset(left_7_3_reset),
    .write_en(left_7_3_write_en)
);
mac_pe pe_7_4 (
    .clk(pe_7_4_clk),
    .done(pe_7_4_done),
    .go(pe_7_4_go),
    .left(pe_7_4_left),
    .mul_ready(pe_7_4_mul_ready),
    .out(pe_7_4_out),
    .reset(pe_7_4_reset),
    .top(pe_7_4_top)
);
std_reg # (
    .WIDTH(32)
) top_7_4 (
    .clk(top_7_4_clk),
    .done(top_7_4_done),
    .in(top_7_4_in),
    .out(top_7_4_out),
    .reset(top_7_4_reset),
    .write_en(top_7_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_4 (
    .clk(left_7_4_clk),
    .done(left_7_4_done),
    .in(left_7_4_in),
    .out(left_7_4_out),
    .reset(left_7_4_reset),
    .write_en(left_7_4_write_en)
);
mac_pe pe_7_5 (
    .clk(pe_7_5_clk),
    .done(pe_7_5_done),
    .go(pe_7_5_go),
    .left(pe_7_5_left),
    .mul_ready(pe_7_5_mul_ready),
    .out(pe_7_5_out),
    .reset(pe_7_5_reset),
    .top(pe_7_5_top)
);
std_reg # (
    .WIDTH(32)
) top_7_5 (
    .clk(top_7_5_clk),
    .done(top_7_5_done),
    .in(top_7_5_in),
    .out(top_7_5_out),
    .reset(top_7_5_reset),
    .write_en(top_7_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_5 (
    .clk(left_7_5_clk),
    .done(left_7_5_done),
    .in(left_7_5_in),
    .out(left_7_5_out),
    .reset(left_7_5_reset),
    .write_en(left_7_5_write_en)
);
mac_pe pe_7_6 (
    .clk(pe_7_6_clk),
    .done(pe_7_6_done),
    .go(pe_7_6_go),
    .left(pe_7_6_left),
    .mul_ready(pe_7_6_mul_ready),
    .out(pe_7_6_out),
    .reset(pe_7_6_reset),
    .top(pe_7_6_top)
);
std_reg # (
    .WIDTH(32)
) top_7_6 (
    .clk(top_7_6_clk),
    .done(top_7_6_done),
    .in(top_7_6_in),
    .out(top_7_6_out),
    .reset(top_7_6_reset),
    .write_en(top_7_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_6 (
    .clk(left_7_6_clk),
    .done(left_7_6_done),
    .in(left_7_6_in),
    .out(left_7_6_out),
    .reset(left_7_6_reset),
    .write_en(left_7_6_write_en)
);
mac_pe pe_7_7 (
    .clk(pe_7_7_clk),
    .done(pe_7_7_done),
    .go(pe_7_7_go),
    .left(pe_7_7_left),
    .mul_ready(pe_7_7_mul_ready),
    .out(pe_7_7_out),
    .reset(pe_7_7_reset),
    .top(pe_7_7_top)
);
std_reg # (
    .WIDTH(32)
) top_7_7 (
    .clk(top_7_7_clk),
    .done(top_7_7_done),
    .in(top_7_7_in),
    .out(top_7_7_out),
    .reset(top_7_7_reset),
    .write_en(top_7_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_7 (
    .clk(left_7_7_clk),
    .done(left_7_7_done),
    .in(left_7_7_in),
    .out(left_7_7_out),
    .reset(left_7_7_reset),
    .write_en(left_7_7_write_en)
);
mac_pe pe_7_8 (
    .clk(pe_7_8_clk),
    .done(pe_7_8_done),
    .go(pe_7_8_go),
    .left(pe_7_8_left),
    .mul_ready(pe_7_8_mul_ready),
    .out(pe_7_8_out),
    .reset(pe_7_8_reset),
    .top(pe_7_8_top)
);
std_reg # (
    .WIDTH(32)
) top_7_8 (
    .clk(top_7_8_clk),
    .done(top_7_8_done),
    .in(top_7_8_in),
    .out(top_7_8_out),
    .reset(top_7_8_reset),
    .write_en(top_7_8_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_8 (
    .clk(left_7_8_clk),
    .done(left_7_8_done),
    .in(left_7_8_in),
    .out(left_7_8_out),
    .reset(left_7_8_reset),
    .write_en(left_7_8_write_en)
);
mac_pe pe_7_9 (
    .clk(pe_7_9_clk),
    .done(pe_7_9_done),
    .go(pe_7_9_go),
    .left(pe_7_9_left),
    .mul_ready(pe_7_9_mul_ready),
    .out(pe_7_9_out),
    .reset(pe_7_9_reset),
    .top(pe_7_9_top)
);
std_reg # (
    .WIDTH(32)
) top_7_9 (
    .clk(top_7_9_clk),
    .done(top_7_9_done),
    .in(top_7_9_in),
    .out(top_7_9_out),
    .reset(top_7_9_reset),
    .write_en(top_7_9_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_9 (
    .clk(left_7_9_clk),
    .done(left_7_9_done),
    .in(left_7_9_in),
    .out(left_7_9_out),
    .reset(left_7_9_reset),
    .write_en(left_7_9_write_en)
);
mac_pe pe_7_10 (
    .clk(pe_7_10_clk),
    .done(pe_7_10_done),
    .go(pe_7_10_go),
    .left(pe_7_10_left),
    .mul_ready(pe_7_10_mul_ready),
    .out(pe_7_10_out),
    .reset(pe_7_10_reset),
    .top(pe_7_10_top)
);
std_reg # (
    .WIDTH(32)
) top_7_10 (
    .clk(top_7_10_clk),
    .done(top_7_10_done),
    .in(top_7_10_in),
    .out(top_7_10_out),
    .reset(top_7_10_reset),
    .write_en(top_7_10_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_10 (
    .clk(left_7_10_clk),
    .done(left_7_10_done),
    .in(left_7_10_in),
    .out(left_7_10_out),
    .reset(left_7_10_reset),
    .write_en(left_7_10_write_en)
);
mac_pe pe_7_11 (
    .clk(pe_7_11_clk),
    .done(pe_7_11_done),
    .go(pe_7_11_go),
    .left(pe_7_11_left),
    .mul_ready(pe_7_11_mul_ready),
    .out(pe_7_11_out),
    .reset(pe_7_11_reset),
    .top(pe_7_11_top)
);
std_reg # (
    .WIDTH(32)
) top_7_11 (
    .clk(top_7_11_clk),
    .done(top_7_11_done),
    .in(top_7_11_in),
    .out(top_7_11_out),
    .reset(top_7_11_reset),
    .write_en(top_7_11_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_11 (
    .clk(left_7_11_clk),
    .done(left_7_11_done),
    .in(left_7_11_in),
    .out(left_7_11_out),
    .reset(left_7_11_reset),
    .write_en(left_7_11_write_en)
);
mac_pe pe_7_12 (
    .clk(pe_7_12_clk),
    .done(pe_7_12_done),
    .go(pe_7_12_go),
    .left(pe_7_12_left),
    .mul_ready(pe_7_12_mul_ready),
    .out(pe_7_12_out),
    .reset(pe_7_12_reset),
    .top(pe_7_12_top)
);
std_reg # (
    .WIDTH(32)
) top_7_12 (
    .clk(top_7_12_clk),
    .done(top_7_12_done),
    .in(top_7_12_in),
    .out(top_7_12_out),
    .reset(top_7_12_reset),
    .write_en(top_7_12_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_12 (
    .clk(left_7_12_clk),
    .done(left_7_12_done),
    .in(left_7_12_in),
    .out(left_7_12_out),
    .reset(left_7_12_reset),
    .write_en(left_7_12_write_en)
);
mac_pe pe_7_13 (
    .clk(pe_7_13_clk),
    .done(pe_7_13_done),
    .go(pe_7_13_go),
    .left(pe_7_13_left),
    .mul_ready(pe_7_13_mul_ready),
    .out(pe_7_13_out),
    .reset(pe_7_13_reset),
    .top(pe_7_13_top)
);
std_reg # (
    .WIDTH(32)
) top_7_13 (
    .clk(top_7_13_clk),
    .done(top_7_13_done),
    .in(top_7_13_in),
    .out(top_7_13_out),
    .reset(top_7_13_reset),
    .write_en(top_7_13_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_13 (
    .clk(left_7_13_clk),
    .done(left_7_13_done),
    .in(left_7_13_in),
    .out(left_7_13_out),
    .reset(left_7_13_reset),
    .write_en(left_7_13_write_en)
);
mac_pe pe_7_14 (
    .clk(pe_7_14_clk),
    .done(pe_7_14_done),
    .go(pe_7_14_go),
    .left(pe_7_14_left),
    .mul_ready(pe_7_14_mul_ready),
    .out(pe_7_14_out),
    .reset(pe_7_14_reset),
    .top(pe_7_14_top)
);
std_reg # (
    .WIDTH(32)
) top_7_14 (
    .clk(top_7_14_clk),
    .done(top_7_14_done),
    .in(top_7_14_in),
    .out(top_7_14_out),
    .reset(top_7_14_reset),
    .write_en(top_7_14_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_14 (
    .clk(left_7_14_clk),
    .done(left_7_14_done),
    .in(left_7_14_in),
    .out(left_7_14_out),
    .reset(left_7_14_reset),
    .write_en(left_7_14_write_en)
);
mac_pe pe_7_15 (
    .clk(pe_7_15_clk),
    .done(pe_7_15_done),
    .go(pe_7_15_go),
    .left(pe_7_15_left),
    .mul_ready(pe_7_15_mul_ready),
    .out(pe_7_15_out),
    .reset(pe_7_15_reset),
    .top(pe_7_15_top)
);
std_reg # (
    .WIDTH(32)
) top_7_15 (
    .clk(top_7_15_clk),
    .done(top_7_15_done),
    .in(top_7_15_in),
    .out(top_7_15_out),
    .reset(top_7_15_reset),
    .write_en(top_7_15_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_15 (
    .clk(left_7_15_clk),
    .done(left_7_15_done),
    .in(left_7_15_in),
    .out(left_7_15_out),
    .reset(left_7_15_reset),
    .write_en(left_7_15_write_en)
);
mac_pe pe_8_0 (
    .clk(pe_8_0_clk),
    .done(pe_8_0_done),
    .go(pe_8_0_go),
    .left(pe_8_0_left),
    .mul_ready(pe_8_0_mul_ready),
    .out(pe_8_0_out),
    .reset(pe_8_0_reset),
    .top(pe_8_0_top)
);
std_reg # (
    .WIDTH(32)
) top_8_0 (
    .clk(top_8_0_clk),
    .done(top_8_0_done),
    .in(top_8_0_in),
    .out(top_8_0_out),
    .reset(top_8_0_reset),
    .write_en(top_8_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_8_0 (
    .clk(left_8_0_clk),
    .done(left_8_0_done),
    .in(left_8_0_in),
    .out(left_8_0_out),
    .reset(left_8_0_reset),
    .write_en(left_8_0_write_en)
);
mac_pe pe_8_1 (
    .clk(pe_8_1_clk),
    .done(pe_8_1_done),
    .go(pe_8_1_go),
    .left(pe_8_1_left),
    .mul_ready(pe_8_1_mul_ready),
    .out(pe_8_1_out),
    .reset(pe_8_1_reset),
    .top(pe_8_1_top)
);
std_reg # (
    .WIDTH(32)
) top_8_1 (
    .clk(top_8_1_clk),
    .done(top_8_1_done),
    .in(top_8_1_in),
    .out(top_8_1_out),
    .reset(top_8_1_reset),
    .write_en(top_8_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_8_1 (
    .clk(left_8_1_clk),
    .done(left_8_1_done),
    .in(left_8_1_in),
    .out(left_8_1_out),
    .reset(left_8_1_reset),
    .write_en(left_8_1_write_en)
);
mac_pe pe_8_2 (
    .clk(pe_8_2_clk),
    .done(pe_8_2_done),
    .go(pe_8_2_go),
    .left(pe_8_2_left),
    .mul_ready(pe_8_2_mul_ready),
    .out(pe_8_2_out),
    .reset(pe_8_2_reset),
    .top(pe_8_2_top)
);
std_reg # (
    .WIDTH(32)
) top_8_2 (
    .clk(top_8_2_clk),
    .done(top_8_2_done),
    .in(top_8_2_in),
    .out(top_8_2_out),
    .reset(top_8_2_reset),
    .write_en(top_8_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_8_2 (
    .clk(left_8_2_clk),
    .done(left_8_2_done),
    .in(left_8_2_in),
    .out(left_8_2_out),
    .reset(left_8_2_reset),
    .write_en(left_8_2_write_en)
);
mac_pe pe_8_3 (
    .clk(pe_8_3_clk),
    .done(pe_8_3_done),
    .go(pe_8_3_go),
    .left(pe_8_3_left),
    .mul_ready(pe_8_3_mul_ready),
    .out(pe_8_3_out),
    .reset(pe_8_3_reset),
    .top(pe_8_3_top)
);
std_reg # (
    .WIDTH(32)
) top_8_3 (
    .clk(top_8_3_clk),
    .done(top_8_3_done),
    .in(top_8_3_in),
    .out(top_8_3_out),
    .reset(top_8_3_reset),
    .write_en(top_8_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_8_3 (
    .clk(left_8_3_clk),
    .done(left_8_3_done),
    .in(left_8_3_in),
    .out(left_8_3_out),
    .reset(left_8_3_reset),
    .write_en(left_8_3_write_en)
);
mac_pe pe_8_4 (
    .clk(pe_8_4_clk),
    .done(pe_8_4_done),
    .go(pe_8_4_go),
    .left(pe_8_4_left),
    .mul_ready(pe_8_4_mul_ready),
    .out(pe_8_4_out),
    .reset(pe_8_4_reset),
    .top(pe_8_4_top)
);
std_reg # (
    .WIDTH(32)
) top_8_4 (
    .clk(top_8_4_clk),
    .done(top_8_4_done),
    .in(top_8_4_in),
    .out(top_8_4_out),
    .reset(top_8_4_reset),
    .write_en(top_8_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_8_4 (
    .clk(left_8_4_clk),
    .done(left_8_4_done),
    .in(left_8_4_in),
    .out(left_8_4_out),
    .reset(left_8_4_reset),
    .write_en(left_8_4_write_en)
);
mac_pe pe_8_5 (
    .clk(pe_8_5_clk),
    .done(pe_8_5_done),
    .go(pe_8_5_go),
    .left(pe_8_5_left),
    .mul_ready(pe_8_5_mul_ready),
    .out(pe_8_5_out),
    .reset(pe_8_5_reset),
    .top(pe_8_5_top)
);
std_reg # (
    .WIDTH(32)
) top_8_5 (
    .clk(top_8_5_clk),
    .done(top_8_5_done),
    .in(top_8_5_in),
    .out(top_8_5_out),
    .reset(top_8_5_reset),
    .write_en(top_8_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_8_5 (
    .clk(left_8_5_clk),
    .done(left_8_5_done),
    .in(left_8_5_in),
    .out(left_8_5_out),
    .reset(left_8_5_reset),
    .write_en(left_8_5_write_en)
);
mac_pe pe_8_6 (
    .clk(pe_8_6_clk),
    .done(pe_8_6_done),
    .go(pe_8_6_go),
    .left(pe_8_6_left),
    .mul_ready(pe_8_6_mul_ready),
    .out(pe_8_6_out),
    .reset(pe_8_6_reset),
    .top(pe_8_6_top)
);
std_reg # (
    .WIDTH(32)
) top_8_6 (
    .clk(top_8_6_clk),
    .done(top_8_6_done),
    .in(top_8_6_in),
    .out(top_8_6_out),
    .reset(top_8_6_reset),
    .write_en(top_8_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_8_6 (
    .clk(left_8_6_clk),
    .done(left_8_6_done),
    .in(left_8_6_in),
    .out(left_8_6_out),
    .reset(left_8_6_reset),
    .write_en(left_8_6_write_en)
);
mac_pe pe_8_7 (
    .clk(pe_8_7_clk),
    .done(pe_8_7_done),
    .go(pe_8_7_go),
    .left(pe_8_7_left),
    .mul_ready(pe_8_7_mul_ready),
    .out(pe_8_7_out),
    .reset(pe_8_7_reset),
    .top(pe_8_7_top)
);
std_reg # (
    .WIDTH(32)
) top_8_7 (
    .clk(top_8_7_clk),
    .done(top_8_7_done),
    .in(top_8_7_in),
    .out(top_8_7_out),
    .reset(top_8_7_reset),
    .write_en(top_8_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_8_7 (
    .clk(left_8_7_clk),
    .done(left_8_7_done),
    .in(left_8_7_in),
    .out(left_8_7_out),
    .reset(left_8_7_reset),
    .write_en(left_8_7_write_en)
);
mac_pe pe_8_8 (
    .clk(pe_8_8_clk),
    .done(pe_8_8_done),
    .go(pe_8_8_go),
    .left(pe_8_8_left),
    .mul_ready(pe_8_8_mul_ready),
    .out(pe_8_8_out),
    .reset(pe_8_8_reset),
    .top(pe_8_8_top)
);
std_reg # (
    .WIDTH(32)
) top_8_8 (
    .clk(top_8_8_clk),
    .done(top_8_8_done),
    .in(top_8_8_in),
    .out(top_8_8_out),
    .reset(top_8_8_reset),
    .write_en(top_8_8_write_en)
);
std_reg # (
    .WIDTH(32)
) left_8_8 (
    .clk(left_8_8_clk),
    .done(left_8_8_done),
    .in(left_8_8_in),
    .out(left_8_8_out),
    .reset(left_8_8_reset),
    .write_en(left_8_8_write_en)
);
mac_pe pe_8_9 (
    .clk(pe_8_9_clk),
    .done(pe_8_9_done),
    .go(pe_8_9_go),
    .left(pe_8_9_left),
    .mul_ready(pe_8_9_mul_ready),
    .out(pe_8_9_out),
    .reset(pe_8_9_reset),
    .top(pe_8_9_top)
);
std_reg # (
    .WIDTH(32)
) top_8_9 (
    .clk(top_8_9_clk),
    .done(top_8_9_done),
    .in(top_8_9_in),
    .out(top_8_9_out),
    .reset(top_8_9_reset),
    .write_en(top_8_9_write_en)
);
std_reg # (
    .WIDTH(32)
) left_8_9 (
    .clk(left_8_9_clk),
    .done(left_8_9_done),
    .in(left_8_9_in),
    .out(left_8_9_out),
    .reset(left_8_9_reset),
    .write_en(left_8_9_write_en)
);
mac_pe pe_8_10 (
    .clk(pe_8_10_clk),
    .done(pe_8_10_done),
    .go(pe_8_10_go),
    .left(pe_8_10_left),
    .mul_ready(pe_8_10_mul_ready),
    .out(pe_8_10_out),
    .reset(pe_8_10_reset),
    .top(pe_8_10_top)
);
std_reg # (
    .WIDTH(32)
) top_8_10 (
    .clk(top_8_10_clk),
    .done(top_8_10_done),
    .in(top_8_10_in),
    .out(top_8_10_out),
    .reset(top_8_10_reset),
    .write_en(top_8_10_write_en)
);
std_reg # (
    .WIDTH(32)
) left_8_10 (
    .clk(left_8_10_clk),
    .done(left_8_10_done),
    .in(left_8_10_in),
    .out(left_8_10_out),
    .reset(left_8_10_reset),
    .write_en(left_8_10_write_en)
);
mac_pe pe_8_11 (
    .clk(pe_8_11_clk),
    .done(pe_8_11_done),
    .go(pe_8_11_go),
    .left(pe_8_11_left),
    .mul_ready(pe_8_11_mul_ready),
    .out(pe_8_11_out),
    .reset(pe_8_11_reset),
    .top(pe_8_11_top)
);
std_reg # (
    .WIDTH(32)
) top_8_11 (
    .clk(top_8_11_clk),
    .done(top_8_11_done),
    .in(top_8_11_in),
    .out(top_8_11_out),
    .reset(top_8_11_reset),
    .write_en(top_8_11_write_en)
);
std_reg # (
    .WIDTH(32)
) left_8_11 (
    .clk(left_8_11_clk),
    .done(left_8_11_done),
    .in(left_8_11_in),
    .out(left_8_11_out),
    .reset(left_8_11_reset),
    .write_en(left_8_11_write_en)
);
mac_pe pe_8_12 (
    .clk(pe_8_12_clk),
    .done(pe_8_12_done),
    .go(pe_8_12_go),
    .left(pe_8_12_left),
    .mul_ready(pe_8_12_mul_ready),
    .out(pe_8_12_out),
    .reset(pe_8_12_reset),
    .top(pe_8_12_top)
);
std_reg # (
    .WIDTH(32)
) top_8_12 (
    .clk(top_8_12_clk),
    .done(top_8_12_done),
    .in(top_8_12_in),
    .out(top_8_12_out),
    .reset(top_8_12_reset),
    .write_en(top_8_12_write_en)
);
std_reg # (
    .WIDTH(32)
) left_8_12 (
    .clk(left_8_12_clk),
    .done(left_8_12_done),
    .in(left_8_12_in),
    .out(left_8_12_out),
    .reset(left_8_12_reset),
    .write_en(left_8_12_write_en)
);
mac_pe pe_8_13 (
    .clk(pe_8_13_clk),
    .done(pe_8_13_done),
    .go(pe_8_13_go),
    .left(pe_8_13_left),
    .mul_ready(pe_8_13_mul_ready),
    .out(pe_8_13_out),
    .reset(pe_8_13_reset),
    .top(pe_8_13_top)
);
std_reg # (
    .WIDTH(32)
) top_8_13 (
    .clk(top_8_13_clk),
    .done(top_8_13_done),
    .in(top_8_13_in),
    .out(top_8_13_out),
    .reset(top_8_13_reset),
    .write_en(top_8_13_write_en)
);
std_reg # (
    .WIDTH(32)
) left_8_13 (
    .clk(left_8_13_clk),
    .done(left_8_13_done),
    .in(left_8_13_in),
    .out(left_8_13_out),
    .reset(left_8_13_reset),
    .write_en(left_8_13_write_en)
);
mac_pe pe_8_14 (
    .clk(pe_8_14_clk),
    .done(pe_8_14_done),
    .go(pe_8_14_go),
    .left(pe_8_14_left),
    .mul_ready(pe_8_14_mul_ready),
    .out(pe_8_14_out),
    .reset(pe_8_14_reset),
    .top(pe_8_14_top)
);
std_reg # (
    .WIDTH(32)
) top_8_14 (
    .clk(top_8_14_clk),
    .done(top_8_14_done),
    .in(top_8_14_in),
    .out(top_8_14_out),
    .reset(top_8_14_reset),
    .write_en(top_8_14_write_en)
);
std_reg # (
    .WIDTH(32)
) left_8_14 (
    .clk(left_8_14_clk),
    .done(left_8_14_done),
    .in(left_8_14_in),
    .out(left_8_14_out),
    .reset(left_8_14_reset),
    .write_en(left_8_14_write_en)
);
mac_pe pe_8_15 (
    .clk(pe_8_15_clk),
    .done(pe_8_15_done),
    .go(pe_8_15_go),
    .left(pe_8_15_left),
    .mul_ready(pe_8_15_mul_ready),
    .out(pe_8_15_out),
    .reset(pe_8_15_reset),
    .top(pe_8_15_top)
);
std_reg # (
    .WIDTH(32)
) top_8_15 (
    .clk(top_8_15_clk),
    .done(top_8_15_done),
    .in(top_8_15_in),
    .out(top_8_15_out),
    .reset(top_8_15_reset),
    .write_en(top_8_15_write_en)
);
std_reg # (
    .WIDTH(32)
) left_8_15 (
    .clk(left_8_15_clk),
    .done(left_8_15_done),
    .in(left_8_15_in),
    .out(left_8_15_out),
    .reset(left_8_15_reset),
    .write_en(left_8_15_write_en)
);
mac_pe pe_9_0 (
    .clk(pe_9_0_clk),
    .done(pe_9_0_done),
    .go(pe_9_0_go),
    .left(pe_9_0_left),
    .mul_ready(pe_9_0_mul_ready),
    .out(pe_9_0_out),
    .reset(pe_9_0_reset),
    .top(pe_9_0_top)
);
std_reg # (
    .WIDTH(32)
) top_9_0 (
    .clk(top_9_0_clk),
    .done(top_9_0_done),
    .in(top_9_0_in),
    .out(top_9_0_out),
    .reset(top_9_0_reset),
    .write_en(top_9_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_9_0 (
    .clk(left_9_0_clk),
    .done(left_9_0_done),
    .in(left_9_0_in),
    .out(left_9_0_out),
    .reset(left_9_0_reset),
    .write_en(left_9_0_write_en)
);
mac_pe pe_9_1 (
    .clk(pe_9_1_clk),
    .done(pe_9_1_done),
    .go(pe_9_1_go),
    .left(pe_9_1_left),
    .mul_ready(pe_9_1_mul_ready),
    .out(pe_9_1_out),
    .reset(pe_9_1_reset),
    .top(pe_9_1_top)
);
std_reg # (
    .WIDTH(32)
) top_9_1 (
    .clk(top_9_1_clk),
    .done(top_9_1_done),
    .in(top_9_1_in),
    .out(top_9_1_out),
    .reset(top_9_1_reset),
    .write_en(top_9_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_9_1 (
    .clk(left_9_1_clk),
    .done(left_9_1_done),
    .in(left_9_1_in),
    .out(left_9_1_out),
    .reset(left_9_1_reset),
    .write_en(left_9_1_write_en)
);
mac_pe pe_9_2 (
    .clk(pe_9_2_clk),
    .done(pe_9_2_done),
    .go(pe_9_2_go),
    .left(pe_9_2_left),
    .mul_ready(pe_9_2_mul_ready),
    .out(pe_9_2_out),
    .reset(pe_9_2_reset),
    .top(pe_9_2_top)
);
std_reg # (
    .WIDTH(32)
) top_9_2 (
    .clk(top_9_2_clk),
    .done(top_9_2_done),
    .in(top_9_2_in),
    .out(top_9_2_out),
    .reset(top_9_2_reset),
    .write_en(top_9_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_9_2 (
    .clk(left_9_2_clk),
    .done(left_9_2_done),
    .in(left_9_2_in),
    .out(left_9_2_out),
    .reset(left_9_2_reset),
    .write_en(left_9_2_write_en)
);
mac_pe pe_9_3 (
    .clk(pe_9_3_clk),
    .done(pe_9_3_done),
    .go(pe_9_3_go),
    .left(pe_9_3_left),
    .mul_ready(pe_9_3_mul_ready),
    .out(pe_9_3_out),
    .reset(pe_9_3_reset),
    .top(pe_9_3_top)
);
std_reg # (
    .WIDTH(32)
) top_9_3 (
    .clk(top_9_3_clk),
    .done(top_9_3_done),
    .in(top_9_3_in),
    .out(top_9_3_out),
    .reset(top_9_3_reset),
    .write_en(top_9_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_9_3 (
    .clk(left_9_3_clk),
    .done(left_9_3_done),
    .in(left_9_3_in),
    .out(left_9_3_out),
    .reset(left_9_3_reset),
    .write_en(left_9_3_write_en)
);
mac_pe pe_9_4 (
    .clk(pe_9_4_clk),
    .done(pe_9_4_done),
    .go(pe_9_4_go),
    .left(pe_9_4_left),
    .mul_ready(pe_9_4_mul_ready),
    .out(pe_9_4_out),
    .reset(pe_9_4_reset),
    .top(pe_9_4_top)
);
std_reg # (
    .WIDTH(32)
) top_9_4 (
    .clk(top_9_4_clk),
    .done(top_9_4_done),
    .in(top_9_4_in),
    .out(top_9_4_out),
    .reset(top_9_4_reset),
    .write_en(top_9_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_9_4 (
    .clk(left_9_4_clk),
    .done(left_9_4_done),
    .in(left_9_4_in),
    .out(left_9_4_out),
    .reset(left_9_4_reset),
    .write_en(left_9_4_write_en)
);
mac_pe pe_9_5 (
    .clk(pe_9_5_clk),
    .done(pe_9_5_done),
    .go(pe_9_5_go),
    .left(pe_9_5_left),
    .mul_ready(pe_9_5_mul_ready),
    .out(pe_9_5_out),
    .reset(pe_9_5_reset),
    .top(pe_9_5_top)
);
std_reg # (
    .WIDTH(32)
) top_9_5 (
    .clk(top_9_5_clk),
    .done(top_9_5_done),
    .in(top_9_5_in),
    .out(top_9_5_out),
    .reset(top_9_5_reset),
    .write_en(top_9_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_9_5 (
    .clk(left_9_5_clk),
    .done(left_9_5_done),
    .in(left_9_5_in),
    .out(left_9_5_out),
    .reset(left_9_5_reset),
    .write_en(left_9_5_write_en)
);
mac_pe pe_9_6 (
    .clk(pe_9_6_clk),
    .done(pe_9_6_done),
    .go(pe_9_6_go),
    .left(pe_9_6_left),
    .mul_ready(pe_9_6_mul_ready),
    .out(pe_9_6_out),
    .reset(pe_9_6_reset),
    .top(pe_9_6_top)
);
std_reg # (
    .WIDTH(32)
) top_9_6 (
    .clk(top_9_6_clk),
    .done(top_9_6_done),
    .in(top_9_6_in),
    .out(top_9_6_out),
    .reset(top_9_6_reset),
    .write_en(top_9_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_9_6 (
    .clk(left_9_6_clk),
    .done(left_9_6_done),
    .in(left_9_6_in),
    .out(left_9_6_out),
    .reset(left_9_6_reset),
    .write_en(left_9_6_write_en)
);
mac_pe pe_9_7 (
    .clk(pe_9_7_clk),
    .done(pe_9_7_done),
    .go(pe_9_7_go),
    .left(pe_9_7_left),
    .mul_ready(pe_9_7_mul_ready),
    .out(pe_9_7_out),
    .reset(pe_9_7_reset),
    .top(pe_9_7_top)
);
std_reg # (
    .WIDTH(32)
) top_9_7 (
    .clk(top_9_7_clk),
    .done(top_9_7_done),
    .in(top_9_7_in),
    .out(top_9_7_out),
    .reset(top_9_7_reset),
    .write_en(top_9_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_9_7 (
    .clk(left_9_7_clk),
    .done(left_9_7_done),
    .in(left_9_7_in),
    .out(left_9_7_out),
    .reset(left_9_7_reset),
    .write_en(left_9_7_write_en)
);
mac_pe pe_9_8 (
    .clk(pe_9_8_clk),
    .done(pe_9_8_done),
    .go(pe_9_8_go),
    .left(pe_9_8_left),
    .mul_ready(pe_9_8_mul_ready),
    .out(pe_9_8_out),
    .reset(pe_9_8_reset),
    .top(pe_9_8_top)
);
std_reg # (
    .WIDTH(32)
) top_9_8 (
    .clk(top_9_8_clk),
    .done(top_9_8_done),
    .in(top_9_8_in),
    .out(top_9_8_out),
    .reset(top_9_8_reset),
    .write_en(top_9_8_write_en)
);
std_reg # (
    .WIDTH(32)
) left_9_8 (
    .clk(left_9_8_clk),
    .done(left_9_8_done),
    .in(left_9_8_in),
    .out(left_9_8_out),
    .reset(left_9_8_reset),
    .write_en(left_9_8_write_en)
);
mac_pe pe_9_9 (
    .clk(pe_9_9_clk),
    .done(pe_9_9_done),
    .go(pe_9_9_go),
    .left(pe_9_9_left),
    .mul_ready(pe_9_9_mul_ready),
    .out(pe_9_9_out),
    .reset(pe_9_9_reset),
    .top(pe_9_9_top)
);
std_reg # (
    .WIDTH(32)
) top_9_9 (
    .clk(top_9_9_clk),
    .done(top_9_9_done),
    .in(top_9_9_in),
    .out(top_9_9_out),
    .reset(top_9_9_reset),
    .write_en(top_9_9_write_en)
);
std_reg # (
    .WIDTH(32)
) left_9_9 (
    .clk(left_9_9_clk),
    .done(left_9_9_done),
    .in(left_9_9_in),
    .out(left_9_9_out),
    .reset(left_9_9_reset),
    .write_en(left_9_9_write_en)
);
mac_pe pe_9_10 (
    .clk(pe_9_10_clk),
    .done(pe_9_10_done),
    .go(pe_9_10_go),
    .left(pe_9_10_left),
    .mul_ready(pe_9_10_mul_ready),
    .out(pe_9_10_out),
    .reset(pe_9_10_reset),
    .top(pe_9_10_top)
);
std_reg # (
    .WIDTH(32)
) top_9_10 (
    .clk(top_9_10_clk),
    .done(top_9_10_done),
    .in(top_9_10_in),
    .out(top_9_10_out),
    .reset(top_9_10_reset),
    .write_en(top_9_10_write_en)
);
std_reg # (
    .WIDTH(32)
) left_9_10 (
    .clk(left_9_10_clk),
    .done(left_9_10_done),
    .in(left_9_10_in),
    .out(left_9_10_out),
    .reset(left_9_10_reset),
    .write_en(left_9_10_write_en)
);
mac_pe pe_9_11 (
    .clk(pe_9_11_clk),
    .done(pe_9_11_done),
    .go(pe_9_11_go),
    .left(pe_9_11_left),
    .mul_ready(pe_9_11_mul_ready),
    .out(pe_9_11_out),
    .reset(pe_9_11_reset),
    .top(pe_9_11_top)
);
std_reg # (
    .WIDTH(32)
) top_9_11 (
    .clk(top_9_11_clk),
    .done(top_9_11_done),
    .in(top_9_11_in),
    .out(top_9_11_out),
    .reset(top_9_11_reset),
    .write_en(top_9_11_write_en)
);
std_reg # (
    .WIDTH(32)
) left_9_11 (
    .clk(left_9_11_clk),
    .done(left_9_11_done),
    .in(left_9_11_in),
    .out(left_9_11_out),
    .reset(left_9_11_reset),
    .write_en(left_9_11_write_en)
);
mac_pe pe_9_12 (
    .clk(pe_9_12_clk),
    .done(pe_9_12_done),
    .go(pe_9_12_go),
    .left(pe_9_12_left),
    .mul_ready(pe_9_12_mul_ready),
    .out(pe_9_12_out),
    .reset(pe_9_12_reset),
    .top(pe_9_12_top)
);
std_reg # (
    .WIDTH(32)
) top_9_12 (
    .clk(top_9_12_clk),
    .done(top_9_12_done),
    .in(top_9_12_in),
    .out(top_9_12_out),
    .reset(top_9_12_reset),
    .write_en(top_9_12_write_en)
);
std_reg # (
    .WIDTH(32)
) left_9_12 (
    .clk(left_9_12_clk),
    .done(left_9_12_done),
    .in(left_9_12_in),
    .out(left_9_12_out),
    .reset(left_9_12_reset),
    .write_en(left_9_12_write_en)
);
mac_pe pe_9_13 (
    .clk(pe_9_13_clk),
    .done(pe_9_13_done),
    .go(pe_9_13_go),
    .left(pe_9_13_left),
    .mul_ready(pe_9_13_mul_ready),
    .out(pe_9_13_out),
    .reset(pe_9_13_reset),
    .top(pe_9_13_top)
);
std_reg # (
    .WIDTH(32)
) top_9_13 (
    .clk(top_9_13_clk),
    .done(top_9_13_done),
    .in(top_9_13_in),
    .out(top_9_13_out),
    .reset(top_9_13_reset),
    .write_en(top_9_13_write_en)
);
std_reg # (
    .WIDTH(32)
) left_9_13 (
    .clk(left_9_13_clk),
    .done(left_9_13_done),
    .in(left_9_13_in),
    .out(left_9_13_out),
    .reset(left_9_13_reset),
    .write_en(left_9_13_write_en)
);
mac_pe pe_9_14 (
    .clk(pe_9_14_clk),
    .done(pe_9_14_done),
    .go(pe_9_14_go),
    .left(pe_9_14_left),
    .mul_ready(pe_9_14_mul_ready),
    .out(pe_9_14_out),
    .reset(pe_9_14_reset),
    .top(pe_9_14_top)
);
std_reg # (
    .WIDTH(32)
) top_9_14 (
    .clk(top_9_14_clk),
    .done(top_9_14_done),
    .in(top_9_14_in),
    .out(top_9_14_out),
    .reset(top_9_14_reset),
    .write_en(top_9_14_write_en)
);
std_reg # (
    .WIDTH(32)
) left_9_14 (
    .clk(left_9_14_clk),
    .done(left_9_14_done),
    .in(left_9_14_in),
    .out(left_9_14_out),
    .reset(left_9_14_reset),
    .write_en(left_9_14_write_en)
);
mac_pe pe_9_15 (
    .clk(pe_9_15_clk),
    .done(pe_9_15_done),
    .go(pe_9_15_go),
    .left(pe_9_15_left),
    .mul_ready(pe_9_15_mul_ready),
    .out(pe_9_15_out),
    .reset(pe_9_15_reset),
    .top(pe_9_15_top)
);
std_reg # (
    .WIDTH(32)
) top_9_15 (
    .clk(top_9_15_clk),
    .done(top_9_15_done),
    .in(top_9_15_in),
    .out(top_9_15_out),
    .reset(top_9_15_reset),
    .write_en(top_9_15_write_en)
);
std_reg # (
    .WIDTH(32)
) left_9_15 (
    .clk(left_9_15_clk),
    .done(left_9_15_done),
    .in(left_9_15_in),
    .out(left_9_15_out),
    .reset(left_9_15_reset),
    .write_en(left_9_15_write_en)
);
mac_pe pe_10_0 (
    .clk(pe_10_0_clk),
    .done(pe_10_0_done),
    .go(pe_10_0_go),
    .left(pe_10_0_left),
    .mul_ready(pe_10_0_mul_ready),
    .out(pe_10_0_out),
    .reset(pe_10_0_reset),
    .top(pe_10_0_top)
);
std_reg # (
    .WIDTH(32)
) top_10_0 (
    .clk(top_10_0_clk),
    .done(top_10_0_done),
    .in(top_10_0_in),
    .out(top_10_0_out),
    .reset(top_10_0_reset),
    .write_en(top_10_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_10_0 (
    .clk(left_10_0_clk),
    .done(left_10_0_done),
    .in(left_10_0_in),
    .out(left_10_0_out),
    .reset(left_10_0_reset),
    .write_en(left_10_0_write_en)
);
mac_pe pe_10_1 (
    .clk(pe_10_1_clk),
    .done(pe_10_1_done),
    .go(pe_10_1_go),
    .left(pe_10_1_left),
    .mul_ready(pe_10_1_mul_ready),
    .out(pe_10_1_out),
    .reset(pe_10_1_reset),
    .top(pe_10_1_top)
);
std_reg # (
    .WIDTH(32)
) top_10_1 (
    .clk(top_10_1_clk),
    .done(top_10_1_done),
    .in(top_10_1_in),
    .out(top_10_1_out),
    .reset(top_10_1_reset),
    .write_en(top_10_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_10_1 (
    .clk(left_10_1_clk),
    .done(left_10_1_done),
    .in(left_10_1_in),
    .out(left_10_1_out),
    .reset(left_10_1_reset),
    .write_en(left_10_1_write_en)
);
mac_pe pe_10_2 (
    .clk(pe_10_2_clk),
    .done(pe_10_2_done),
    .go(pe_10_2_go),
    .left(pe_10_2_left),
    .mul_ready(pe_10_2_mul_ready),
    .out(pe_10_2_out),
    .reset(pe_10_2_reset),
    .top(pe_10_2_top)
);
std_reg # (
    .WIDTH(32)
) top_10_2 (
    .clk(top_10_2_clk),
    .done(top_10_2_done),
    .in(top_10_2_in),
    .out(top_10_2_out),
    .reset(top_10_2_reset),
    .write_en(top_10_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_10_2 (
    .clk(left_10_2_clk),
    .done(left_10_2_done),
    .in(left_10_2_in),
    .out(left_10_2_out),
    .reset(left_10_2_reset),
    .write_en(left_10_2_write_en)
);
mac_pe pe_10_3 (
    .clk(pe_10_3_clk),
    .done(pe_10_3_done),
    .go(pe_10_3_go),
    .left(pe_10_3_left),
    .mul_ready(pe_10_3_mul_ready),
    .out(pe_10_3_out),
    .reset(pe_10_3_reset),
    .top(pe_10_3_top)
);
std_reg # (
    .WIDTH(32)
) top_10_3 (
    .clk(top_10_3_clk),
    .done(top_10_3_done),
    .in(top_10_3_in),
    .out(top_10_3_out),
    .reset(top_10_3_reset),
    .write_en(top_10_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_10_3 (
    .clk(left_10_3_clk),
    .done(left_10_3_done),
    .in(left_10_3_in),
    .out(left_10_3_out),
    .reset(left_10_3_reset),
    .write_en(left_10_3_write_en)
);
mac_pe pe_10_4 (
    .clk(pe_10_4_clk),
    .done(pe_10_4_done),
    .go(pe_10_4_go),
    .left(pe_10_4_left),
    .mul_ready(pe_10_4_mul_ready),
    .out(pe_10_4_out),
    .reset(pe_10_4_reset),
    .top(pe_10_4_top)
);
std_reg # (
    .WIDTH(32)
) top_10_4 (
    .clk(top_10_4_clk),
    .done(top_10_4_done),
    .in(top_10_4_in),
    .out(top_10_4_out),
    .reset(top_10_4_reset),
    .write_en(top_10_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_10_4 (
    .clk(left_10_4_clk),
    .done(left_10_4_done),
    .in(left_10_4_in),
    .out(left_10_4_out),
    .reset(left_10_4_reset),
    .write_en(left_10_4_write_en)
);
mac_pe pe_10_5 (
    .clk(pe_10_5_clk),
    .done(pe_10_5_done),
    .go(pe_10_5_go),
    .left(pe_10_5_left),
    .mul_ready(pe_10_5_mul_ready),
    .out(pe_10_5_out),
    .reset(pe_10_5_reset),
    .top(pe_10_5_top)
);
std_reg # (
    .WIDTH(32)
) top_10_5 (
    .clk(top_10_5_clk),
    .done(top_10_5_done),
    .in(top_10_5_in),
    .out(top_10_5_out),
    .reset(top_10_5_reset),
    .write_en(top_10_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_10_5 (
    .clk(left_10_5_clk),
    .done(left_10_5_done),
    .in(left_10_5_in),
    .out(left_10_5_out),
    .reset(left_10_5_reset),
    .write_en(left_10_5_write_en)
);
mac_pe pe_10_6 (
    .clk(pe_10_6_clk),
    .done(pe_10_6_done),
    .go(pe_10_6_go),
    .left(pe_10_6_left),
    .mul_ready(pe_10_6_mul_ready),
    .out(pe_10_6_out),
    .reset(pe_10_6_reset),
    .top(pe_10_6_top)
);
std_reg # (
    .WIDTH(32)
) top_10_6 (
    .clk(top_10_6_clk),
    .done(top_10_6_done),
    .in(top_10_6_in),
    .out(top_10_6_out),
    .reset(top_10_6_reset),
    .write_en(top_10_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_10_6 (
    .clk(left_10_6_clk),
    .done(left_10_6_done),
    .in(left_10_6_in),
    .out(left_10_6_out),
    .reset(left_10_6_reset),
    .write_en(left_10_6_write_en)
);
mac_pe pe_10_7 (
    .clk(pe_10_7_clk),
    .done(pe_10_7_done),
    .go(pe_10_7_go),
    .left(pe_10_7_left),
    .mul_ready(pe_10_7_mul_ready),
    .out(pe_10_7_out),
    .reset(pe_10_7_reset),
    .top(pe_10_7_top)
);
std_reg # (
    .WIDTH(32)
) top_10_7 (
    .clk(top_10_7_clk),
    .done(top_10_7_done),
    .in(top_10_7_in),
    .out(top_10_7_out),
    .reset(top_10_7_reset),
    .write_en(top_10_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_10_7 (
    .clk(left_10_7_clk),
    .done(left_10_7_done),
    .in(left_10_7_in),
    .out(left_10_7_out),
    .reset(left_10_7_reset),
    .write_en(left_10_7_write_en)
);
mac_pe pe_10_8 (
    .clk(pe_10_8_clk),
    .done(pe_10_8_done),
    .go(pe_10_8_go),
    .left(pe_10_8_left),
    .mul_ready(pe_10_8_mul_ready),
    .out(pe_10_8_out),
    .reset(pe_10_8_reset),
    .top(pe_10_8_top)
);
std_reg # (
    .WIDTH(32)
) top_10_8 (
    .clk(top_10_8_clk),
    .done(top_10_8_done),
    .in(top_10_8_in),
    .out(top_10_8_out),
    .reset(top_10_8_reset),
    .write_en(top_10_8_write_en)
);
std_reg # (
    .WIDTH(32)
) left_10_8 (
    .clk(left_10_8_clk),
    .done(left_10_8_done),
    .in(left_10_8_in),
    .out(left_10_8_out),
    .reset(left_10_8_reset),
    .write_en(left_10_8_write_en)
);
mac_pe pe_10_9 (
    .clk(pe_10_9_clk),
    .done(pe_10_9_done),
    .go(pe_10_9_go),
    .left(pe_10_9_left),
    .mul_ready(pe_10_9_mul_ready),
    .out(pe_10_9_out),
    .reset(pe_10_9_reset),
    .top(pe_10_9_top)
);
std_reg # (
    .WIDTH(32)
) top_10_9 (
    .clk(top_10_9_clk),
    .done(top_10_9_done),
    .in(top_10_9_in),
    .out(top_10_9_out),
    .reset(top_10_9_reset),
    .write_en(top_10_9_write_en)
);
std_reg # (
    .WIDTH(32)
) left_10_9 (
    .clk(left_10_9_clk),
    .done(left_10_9_done),
    .in(left_10_9_in),
    .out(left_10_9_out),
    .reset(left_10_9_reset),
    .write_en(left_10_9_write_en)
);
mac_pe pe_10_10 (
    .clk(pe_10_10_clk),
    .done(pe_10_10_done),
    .go(pe_10_10_go),
    .left(pe_10_10_left),
    .mul_ready(pe_10_10_mul_ready),
    .out(pe_10_10_out),
    .reset(pe_10_10_reset),
    .top(pe_10_10_top)
);
std_reg # (
    .WIDTH(32)
) top_10_10 (
    .clk(top_10_10_clk),
    .done(top_10_10_done),
    .in(top_10_10_in),
    .out(top_10_10_out),
    .reset(top_10_10_reset),
    .write_en(top_10_10_write_en)
);
std_reg # (
    .WIDTH(32)
) left_10_10 (
    .clk(left_10_10_clk),
    .done(left_10_10_done),
    .in(left_10_10_in),
    .out(left_10_10_out),
    .reset(left_10_10_reset),
    .write_en(left_10_10_write_en)
);
mac_pe pe_10_11 (
    .clk(pe_10_11_clk),
    .done(pe_10_11_done),
    .go(pe_10_11_go),
    .left(pe_10_11_left),
    .mul_ready(pe_10_11_mul_ready),
    .out(pe_10_11_out),
    .reset(pe_10_11_reset),
    .top(pe_10_11_top)
);
std_reg # (
    .WIDTH(32)
) top_10_11 (
    .clk(top_10_11_clk),
    .done(top_10_11_done),
    .in(top_10_11_in),
    .out(top_10_11_out),
    .reset(top_10_11_reset),
    .write_en(top_10_11_write_en)
);
std_reg # (
    .WIDTH(32)
) left_10_11 (
    .clk(left_10_11_clk),
    .done(left_10_11_done),
    .in(left_10_11_in),
    .out(left_10_11_out),
    .reset(left_10_11_reset),
    .write_en(left_10_11_write_en)
);
mac_pe pe_10_12 (
    .clk(pe_10_12_clk),
    .done(pe_10_12_done),
    .go(pe_10_12_go),
    .left(pe_10_12_left),
    .mul_ready(pe_10_12_mul_ready),
    .out(pe_10_12_out),
    .reset(pe_10_12_reset),
    .top(pe_10_12_top)
);
std_reg # (
    .WIDTH(32)
) top_10_12 (
    .clk(top_10_12_clk),
    .done(top_10_12_done),
    .in(top_10_12_in),
    .out(top_10_12_out),
    .reset(top_10_12_reset),
    .write_en(top_10_12_write_en)
);
std_reg # (
    .WIDTH(32)
) left_10_12 (
    .clk(left_10_12_clk),
    .done(left_10_12_done),
    .in(left_10_12_in),
    .out(left_10_12_out),
    .reset(left_10_12_reset),
    .write_en(left_10_12_write_en)
);
mac_pe pe_10_13 (
    .clk(pe_10_13_clk),
    .done(pe_10_13_done),
    .go(pe_10_13_go),
    .left(pe_10_13_left),
    .mul_ready(pe_10_13_mul_ready),
    .out(pe_10_13_out),
    .reset(pe_10_13_reset),
    .top(pe_10_13_top)
);
std_reg # (
    .WIDTH(32)
) top_10_13 (
    .clk(top_10_13_clk),
    .done(top_10_13_done),
    .in(top_10_13_in),
    .out(top_10_13_out),
    .reset(top_10_13_reset),
    .write_en(top_10_13_write_en)
);
std_reg # (
    .WIDTH(32)
) left_10_13 (
    .clk(left_10_13_clk),
    .done(left_10_13_done),
    .in(left_10_13_in),
    .out(left_10_13_out),
    .reset(left_10_13_reset),
    .write_en(left_10_13_write_en)
);
mac_pe pe_10_14 (
    .clk(pe_10_14_clk),
    .done(pe_10_14_done),
    .go(pe_10_14_go),
    .left(pe_10_14_left),
    .mul_ready(pe_10_14_mul_ready),
    .out(pe_10_14_out),
    .reset(pe_10_14_reset),
    .top(pe_10_14_top)
);
std_reg # (
    .WIDTH(32)
) top_10_14 (
    .clk(top_10_14_clk),
    .done(top_10_14_done),
    .in(top_10_14_in),
    .out(top_10_14_out),
    .reset(top_10_14_reset),
    .write_en(top_10_14_write_en)
);
std_reg # (
    .WIDTH(32)
) left_10_14 (
    .clk(left_10_14_clk),
    .done(left_10_14_done),
    .in(left_10_14_in),
    .out(left_10_14_out),
    .reset(left_10_14_reset),
    .write_en(left_10_14_write_en)
);
mac_pe pe_10_15 (
    .clk(pe_10_15_clk),
    .done(pe_10_15_done),
    .go(pe_10_15_go),
    .left(pe_10_15_left),
    .mul_ready(pe_10_15_mul_ready),
    .out(pe_10_15_out),
    .reset(pe_10_15_reset),
    .top(pe_10_15_top)
);
std_reg # (
    .WIDTH(32)
) top_10_15 (
    .clk(top_10_15_clk),
    .done(top_10_15_done),
    .in(top_10_15_in),
    .out(top_10_15_out),
    .reset(top_10_15_reset),
    .write_en(top_10_15_write_en)
);
std_reg # (
    .WIDTH(32)
) left_10_15 (
    .clk(left_10_15_clk),
    .done(left_10_15_done),
    .in(left_10_15_in),
    .out(left_10_15_out),
    .reset(left_10_15_reset),
    .write_en(left_10_15_write_en)
);
mac_pe pe_11_0 (
    .clk(pe_11_0_clk),
    .done(pe_11_0_done),
    .go(pe_11_0_go),
    .left(pe_11_0_left),
    .mul_ready(pe_11_0_mul_ready),
    .out(pe_11_0_out),
    .reset(pe_11_0_reset),
    .top(pe_11_0_top)
);
std_reg # (
    .WIDTH(32)
) top_11_0 (
    .clk(top_11_0_clk),
    .done(top_11_0_done),
    .in(top_11_0_in),
    .out(top_11_0_out),
    .reset(top_11_0_reset),
    .write_en(top_11_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_11_0 (
    .clk(left_11_0_clk),
    .done(left_11_0_done),
    .in(left_11_0_in),
    .out(left_11_0_out),
    .reset(left_11_0_reset),
    .write_en(left_11_0_write_en)
);
mac_pe pe_11_1 (
    .clk(pe_11_1_clk),
    .done(pe_11_1_done),
    .go(pe_11_1_go),
    .left(pe_11_1_left),
    .mul_ready(pe_11_1_mul_ready),
    .out(pe_11_1_out),
    .reset(pe_11_1_reset),
    .top(pe_11_1_top)
);
std_reg # (
    .WIDTH(32)
) top_11_1 (
    .clk(top_11_1_clk),
    .done(top_11_1_done),
    .in(top_11_1_in),
    .out(top_11_1_out),
    .reset(top_11_1_reset),
    .write_en(top_11_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_11_1 (
    .clk(left_11_1_clk),
    .done(left_11_1_done),
    .in(left_11_1_in),
    .out(left_11_1_out),
    .reset(left_11_1_reset),
    .write_en(left_11_1_write_en)
);
mac_pe pe_11_2 (
    .clk(pe_11_2_clk),
    .done(pe_11_2_done),
    .go(pe_11_2_go),
    .left(pe_11_2_left),
    .mul_ready(pe_11_2_mul_ready),
    .out(pe_11_2_out),
    .reset(pe_11_2_reset),
    .top(pe_11_2_top)
);
std_reg # (
    .WIDTH(32)
) top_11_2 (
    .clk(top_11_2_clk),
    .done(top_11_2_done),
    .in(top_11_2_in),
    .out(top_11_2_out),
    .reset(top_11_2_reset),
    .write_en(top_11_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_11_2 (
    .clk(left_11_2_clk),
    .done(left_11_2_done),
    .in(left_11_2_in),
    .out(left_11_2_out),
    .reset(left_11_2_reset),
    .write_en(left_11_2_write_en)
);
mac_pe pe_11_3 (
    .clk(pe_11_3_clk),
    .done(pe_11_3_done),
    .go(pe_11_3_go),
    .left(pe_11_3_left),
    .mul_ready(pe_11_3_mul_ready),
    .out(pe_11_3_out),
    .reset(pe_11_3_reset),
    .top(pe_11_3_top)
);
std_reg # (
    .WIDTH(32)
) top_11_3 (
    .clk(top_11_3_clk),
    .done(top_11_3_done),
    .in(top_11_3_in),
    .out(top_11_3_out),
    .reset(top_11_3_reset),
    .write_en(top_11_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_11_3 (
    .clk(left_11_3_clk),
    .done(left_11_3_done),
    .in(left_11_3_in),
    .out(left_11_3_out),
    .reset(left_11_3_reset),
    .write_en(left_11_3_write_en)
);
mac_pe pe_11_4 (
    .clk(pe_11_4_clk),
    .done(pe_11_4_done),
    .go(pe_11_4_go),
    .left(pe_11_4_left),
    .mul_ready(pe_11_4_mul_ready),
    .out(pe_11_4_out),
    .reset(pe_11_4_reset),
    .top(pe_11_4_top)
);
std_reg # (
    .WIDTH(32)
) top_11_4 (
    .clk(top_11_4_clk),
    .done(top_11_4_done),
    .in(top_11_4_in),
    .out(top_11_4_out),
    .reset(top_11_4_reset),
    .write_en(top_11_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_11_4 (
    .clk(left_11_4_clk),
    .done(left_11_4_done),
    .in(left_11_4_in),
    .out(left_11_4_out),
    .reset(left_11_4_reset),
    .write_en(left_11_4_write_en)
);
mac_pe pe_11_5 (
    .clk(pe_11_5_clk),
    .done(pe_11_5_done),
    .go(pe_11_5_go),
    .left(pe_11_5_left),
    .mul_ready(pe_11_5_mul_ready),
    .out(pe_11_5_out),
    .reset(pe_11_5_reset),
    .top(pe_11_5_top)
);
std_reg # (
    .WIDTH(32)
) top_11_5 (
    .clk(top_11_5_clk),
    .done(top_11_5_done),
    .in(top_11_5_in),
    .out(top_11_5_out),
    .reset(top_11_5_reset),
    .write_en(top_11_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_11_5 (
    .clk(left_11_5_clk),
    .done(left_11_5_done),
    .in(left_11_5_in),
    .out(left_11_5_out),
    .reset(left_11_5_reset),
    .write_en(left_11_5_write_en)
);
mac_pe pe_11_6 (
    .clk(pe_11_6_clk),
    .done(pe_11_6_done),
    .go(pe_11_6_go),
    .left(pe_11_6_left),
    .mul_ready(pe_11_6_mul_ready),
    .out(pe_11_6_out),
    .reset(pe_11_6_reset),
    .top(pe_11_6_top)
);
std_reg # (
    .WIDTH(32)
) top_11_6 (
    .clk(top_11_6_clk),
    .done(top_11_6_done),
    .in(top_11_6_in),
    .out(top_11_6_out),
    .reset(top_11_6_reset),
    .write_en(top_11_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_11_6 (
    .clk(left_11_6_clk),
    .done(left_11_6_done),
    .in(left_11_6_in),
    .out(left_11_6_out),
    .reset(left_11_6_reset),
    .write_en(left_11_6_write_en)
);
mac_pe pe_11_7 (
    .clk(pe_11_7_clk),
    .done(pe_11_7_done),
    .go(pe_11_7_go),
    .left(pe_11_7_left),
    .mul_ready(pe_11_7_mul_ready),
    .out(pe_11_7_out),
    .reset(pe_11_7_reset),
    .top(pe_11_7_top)
);
std_reg # (
    .WIDTH(32)
) top_11_7 (
    .clk(top_11_7_clk),
    .done(top_11_7_done),
    .in(top_11_7_in),
    .out(top_11_7_out),
    .reset(top_11_7_reset),
    .write_en(top_11_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_11_7 (
    .clk(left_11_7_clk),
    .done(left_11_7_done),
    .in(left_11_7_in),
    .out(left_11_7_out),
    .reset(left_11_7_reset),
    .write_en(left_11_7_write_en)
);
mac_pe pe_11_8 (
    .clk(pe_11_8_clk),
    .done(pe_11_8_done),
    .go(pe_11_8_go),
    .left(pe_11_8_left),
    .mul_ready(pe_11_8_mul_ready),
    .out(pe_11_8_out),
    .reset(pe_11_8_reset),
    .top(pe_11_8_top)
);
std_reg # (
    .WIDTH(32)
) top_11_8 (
    .clk(top_11_8_clk),
    .done(top_11_8_done),
    .in(top_11_8_in),
    .out(top_11_8_out),
    .reset(top_11_8_reset),
    .write_en(top_11_8_write_en)
);
std_reg # (
    .WIDTH(32)
) left_11_8 (
    .clk(left_11_8_clk),
    .done(left_11_8_done),
    .in(left_11_8_in),
    .out(left_11_8_out),
    .reset(left_11_8_reset),
    .write_en(left_11_8_write_en)
);
mac_pe pe_11_9 (
    .clk(pe_11_9_clk),
    .done(pe_11_9_done),
    .go(pe_11_9_go),
    .left(pe_11_9_left),
    .mul_ready(pe_11_9_mul_ready),
    .out(pe_11_9_out),
    .reset(pe_11_9_reset),
    .top(pe_11_9_top)
);
std_reg # (
    .WIDTH(32)
) top_11_9 (
    .clk(top_11_9_clk),
    .done(top_11_9_done),
    .in(top_11_9_in),
    .out(top_11_9_out),
    .reset(top_11_9_reset),
    .write_en(top_11_9_write_en)
);
std_reg # (
    .WIDTH(32)
) left_11_9 (
    .clk(left_11_9_clk),
    .done(left_11_9_done),
    .in(left_11_9_in),
    .out(left_11_9_out),
    .reset(left_11_9_reset),
    .write_en(left_11_9_write_en)
);
mac_pe pe_11_10 (
    .clk(pe_11_10_clk),
    .done(pe_11_10_done),
    .go(pe_11_10_go),
    .left(pe_11_10_left),
    .mul_ready(pe_11_10_mul_ready),
    .out(pe_11_10_out),
    .reset(pe_11_10_reset),
    .top(pe_11_10_top)
);
std_reg # (
    .WIDTH(32)
) top_11_10 (
    .clk(top_11_10_clk),
    .done(top_11_10_done),
    .in(top_11_10_in),
    .out(top_11_10_out),
    .reset(top_11_10_reset),
    .write_en(top_11_10_write_en)
);
std_reg # (
    .WIDTH(32)
) left_11_10 (
    .clk(left_11_10_clk),
    .done(left_11_10_done),
    .in(left_11_10_in),
    .out(left_11_10_out),
    .reset(left_11_10_reset),
    .write_en(left_11_10_write_en)
);
mac_pe pe_11_11 (
    .clk(pe_11_11_clk),
    .done(pe_11_11_done),
    .go(pe_11_11_go),
    .left(pe_11_11_left),
    .mul_ready(pe_11_11_mul_ready),
    .out(pe_11_11_out),
    .reset(pe_11_11_reset),
    .top(pe_11_11_top)
);
std_reg # (
    .WIDTH(32)
) top_11_11 (
    .clk(top_11_11_clk),
    .done(top_11_11_done),
    .in(top_11_11_in),
    .out(top_11_11_out),
    .reset(top_11_11_reset),
    .write_en(top_11_11_write_en)
);
std_reg # (
    .WIDTH(32)
) left_11_11 (
    .clk(left_11_11_clk),
    .done(left_11_11_done),
    .in(left_11_11_in),
    .out(left_11_11_out),
    .reset(left_11_11_reset),
    .write_en(left_11_11_write_en)
);
mac_pe pe_11_12 (
    .clk(pe_11_12_clk),
    .done(pe_11_12_done),
    .go(pe_11_12_go),
    .left(pe_11_12_left),
    .mul_ready(pe_11_12_mul_ready),
    .out(pe_11_12_out),
    .reset(pe_11_12_reset),
    .top(pe_11_12_top)
);
std_reg # (
    .WIDTH(32)
) top_11_12 (
    .clk(top_11_12_clk),
    .done(top_11_12_done),
    .in(top_11_12_in),
    .out(top_11_12_out),
    .reset(top_11_12_reset),
    .write_en(top_11_12_write_en)
);
std_reg # (
    .WIDTH(32)
) left_11_12 (
    .clk(left_11_12_clk),
    .done(left_11_12_done),
    .in(left_11_12_in),
    .out(left_11_12_out),
    .reset(left_11_12_reset),
    .write_en(left_11_12_write_en)
);
mac_pe pe_11_13 (
    .clk(pe_11_13_clk),
    .done(pe_11_13_done),
    .go(pe_11_13_go),
    .left(pe_11_13_left),
    .mul_ready(pe_11_13_mul_ready),
    .out(pe_11_13_out),
    .reset(pe_11_13_reset),
    .top(pe_11_13_top)
);
std_reg # (
    .WIDTH(32)
) top_11_13 (
    .clk(top_11_13_clk),
    .done(top_11_13_done),
    .in(top_11_13_in),
    .out(top_11_13_out),
    .reset(top_11_13_reset),
    .write_en(top_11_13_write_en)
);
std_reg # (
    .WIDTH(32)
) left_11_13 (
    .clk(left_11_13_clk),
    .done(left_11_13_done),
    .in(left_11_13_in),
    .out(left_11_13_out),
    .reset(left_11_13_reset),
    .write_en(left_11_13_write_en)
);
mac_pe pe_11_14 (
    .clk(pe_11_14_clk),
    .done(pe_11_14_done),
    .go(pe_11_14_go),
    .left(pe_11_14_left),
    .mul_ready(pe_11_14_mul_ready),
    .out(pe_11_14_out),
    .reset(pe_11_14_reset),
    .top(pe_11_14_top)
);
std_reg # (
    .WIDTH(32)
) top_11_14 (
    .clk(top_11_14_clk),
    .done(top_11_14_done),
    .in(top_11_14_in),
    .out(top_11_14_out),
    .reset(top_11_14_reset),
    .write_en(top_11_14_write_en)
);
std_reg # (
    .WIDTH(32)
) left_11_14 (
    .clk(left_11_14_clk),
    .done(left_11_14_done),
    .in(left_11_14_in),
    .out(left_11_14_out),
    .reset(left_11_14_reset),
    .write_en(left_11_14_write_en)
);
mac_pe pe_11_15 (
    .clk(pe_11_15_clk),
    .done(pe_11_15_done),
    .go(pe_11_15_go),
    .left(pe_11_15_left),
    .mul_ready(pe_11_15_mul_ready),
    .out(pe_11_15_out),
    .reset(pe_11_15_reset),
    .top(pe_11_15_top)
);
std_reg # (
    .WIDTH(32)
) top_11_15 (
    .clk(top_11_15_clk),
    .done(top_11_15_done),
    .in(top_11_15_in),
    .out(top_11_15_out),
    .reset(top_11_15_reset),
    .write_en(top_11_15_write_en)
);
std_reg # (
    .WIDTH(32)
) left_11_15 (
    .clk(left_11_15_clk),
    .done(left_11_15_done),
    .in(left_11_15_in),
    .out(left_11_15_out),
    .reset(left_11_15_reset),
    .write_en(left_11_15_write_en)
);
mac_pe pe_12_0 (
    .clk(pe_12_0_clk),
    .done(pe_12_0_done),
    .go(pe_12_0_go),
    .left(pe_12_0_left),
    .mul_ready(pe_12_0_mul_ready),
    .out(pe_12_0_out),
    .reset(pe_12_0_reset),
    .top(pe_12_0_top)
);
std_reg # (
    .WIDTH(32)
) top_12_0 (
    .clk(top_12_0_clk),
    .done(top_12_0_done),
    .in(top_12_0_in),
    .out(top_12_0_out),
    .reset(top_12_0_reset),
    .write_en(top_12_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_12_0 (
    .clk(left_12_0_clk),
    .done(left_12_0_done),
    .in(left_12_0_in),
    .out(left_12_0_out),
    .reset(left_12_0_reset),
    .write_en(left_12_0_write_en)
);
mac_pe pe_12_1 (
    .clk(pe_12_1_clk),
    .done(pe_12_1_done),
    .go(pe_12_1_go),
    .left(pe_12_1_left),
    .mul_ready(pe_12_1_mul_ready),
    .out(pe_12_1_out),
    .reset(pe_12_1_reset),
    .top(pe_12_1_top)
);
std_reg # (
    .WIDTH(32)
) top_12_1 (
    .clk(top_12_1_clk),
    .done(top_12_1_done),
    .in(top_12_1_in),
    .out(top_12_1_out),
    .reset(top_12_1_reset),
    .write_en(top_12_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_12_1 (
    .clk(left_12_1_clk),
    .done(left_12_1_done),
    .in(left_12_1_in),
    .out(left_12_1_out),
    .reset(left_12_1_reset),
    .write_en(left_12_1_write_en)
);
mac_pe pe_12_2 (
    .clk(pe_12_2_clk),
    .done(pe_12_2_done),
    .go(pe_12_2_go),
    .left(pe_12_2_left),
    .mul_ready(pe_12_2_mul_ready),
    .out(pe_12_2_out),
    .reset(pe_12_2_reset),
    .top(pe_12_2_top)
);
std_reg # (
    .WIDTH(32)
) top_12_2 (
    .clk(top_12_2_clk),
    .done(top_12_2_done),
    .in(top_12_2_in),
    .out(top_12_2_out),
    .reset(top_12_2_reset),
    .write_en(top_12_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_12_2 (
    .clk(left_12_2_clk),
    .done(left_12_2_done),
    .in(left_12_2_in),
    .out(left_12_2_out),
    .reset(left_12_2_reset),
    .write_en(left_12_2_write_en)
);
mac_pe pe_12_3 (
    .clk(pe_12_3_clk),
    .done(pe_12_3_done),
    .go(pe_12_3_go),
    .left(pe_12_3_left),
    .mul_ready(pe_12_3_mul_ready),
    .out(pe_12_3_out),
    .reset(pe_12_3_reset),
    .top(pe_12_3_top)
);
std_reg # (
    .WIDTH(32)
) top_12_3 (
    .clk(top_12_3_clk),
    .done(top_12_3_done),
    .in(top_12_3_in),
    .out(top_12_3_out),
    .reset(top_12_3_reset),
    .write_en(top_12_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_12_3 (
    .clk(left_12_3_clk),
    .done(left_12_3_done),
    .in(left_12_3_in),
    .out(left_12_3_out),
    .reset(left_12_3_reset),
    .write_en(left_12_3_write_en)
);
mac_pe pe_12_4 (
    .clk(pe_12_4_clk),
    .done(pe_12_4_done),
    .go(pe_12_4_go),
    .left(pe_12_4_left),
    .mul_ready(pe_12_4_mul_ready),
    .out(pe_12_4_out),
    .reset(pe_12_4_reset),
    .top(pe_12_4_top)
);
std_reg # (
    .WIDTH(32)
) top_12_4 (
    .clk(top_12_4_clk),
    .done(top_12_4_done),
    .in(top_12_4_in),
    .out(top_12_4_out),
    .reset(top_12_4_reset),
    .write_en(top_12_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_12_4 (
    .clk(left_12_4_clk),
    .done(left_12_4_done),
    .in(left_12_4_in),
    .out(left_12_4_out),
    .reset(left_12_4_reset),
    .write_en(left_12_4_write_en)
);
mac_pe pe_12_5 (
    .clk(pe_12_5_clk),
    .done(pe_12_5_done),
    .go(pe_12_5_go),
    .left(pe_12_5_left),
    .mul_ready(pe_12_5_mul_ready),
    .out(pe_12_5_out),
    .reset(pe_12_5_reset),
    .top(pe_12_5_top)
);
std_reg # (
    .WIDTH(32)
) top_12_5 (
    .clk(top_12_5_clk),
    .done(top_12_5_done),
    .in(top_12_5_in),
    .out(top_12_5_out),
    .reset(top_12_5_reset),
    .write_en(top_12_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_12_5 (
    .clk(left_12_5_clk),
    .done(left_12_5_done),
    .in(left_12_5_in),
    .out(left_12_5_out),
    .reset(left_12_5_reset),
    .write_en(left_12_5_write_en)
);
mac_pe pe_12_6 (
    .clk(pe_12_6_clk),
    .done(pe_12_6_done),
    .go(pe_12_6_go),
    .left(pe_12_6_left),
    .mul_ready(pe_12_6_mul_ready),
    .out(pe_12_6_out),
    .reset(pe_12_6_reset),
    .top(pe_12_6_top)
);
std_reg # (
    .WIDTH(32)
) top_12_6 (
    .clk(top_12_6_clk),
    .done(top_12_6_done),
    .in(top_12_6_in),
    .out(top_12_6_out),
    .reset(top_12_6_reset),
    .write_en(top_12_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_12_6 (
    .clk(left_12_6_clk),
    .done(left_12_6_done),
    .in(left_12_6_in),
    .out(left_12_6_out),
    .reset(left_12_6_reset),
    .write_en(left_12_6_write_en)
);
mac_pe pe_12_7 (
    .clk(pe_12_7_clk),
    .done(pe_12_7_done),
    .go(pe_12_7_go),
    .left(pe_12_7_left),
    .mul_ready(pe_12_7_mul_ready),
    .out(pe_12_7_out),
    .reset(pe_12_7_reset),
    .top(pe_12_7_top)
);
std_reg # (
    .WIDTH(32)
) top_12_7 (
    .clk(top_12_7_clk),
    .done(top_12_7_done),
    .in(top_12_7_in),
    .out(top_12_7_out),
    .reset(top_12_7_reset),
    .write_en(top_12_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_12_7 (
    .clk(left_12_7_clk),
    .done(left_12_7_done),
    .in(left_12_7_in),
    .out(left_12_7_out),
    .reset(left_12_7_reset),
    .write_en(left_12_7_write_en)
);
mac_pe pe_12_8 (
    .clk(pe_12_8_clk),
    .done(pe_12_8_done),
    .go(pe_12_8_go),
    .left(pe_12_8_left),
    .mul_ready(pe_12_8_mul_ready),
    .out(pe_12_8_out),
    .reset(pe_12_8_reset),
    .top(pe_12_8_top)
);
std_reg # (
    .WIDTH(32)
) top_12_8 (
    .clk(top_12_8_clk),
    .done(top_12_8_done),
    .in(top_12_8_in),
    .out(top_12_8_out),
    .reset(top_12_8_reset),
    .write_en(top_12_8_write_en)
);
std_reg # (
    .WIDTH(32)
) left_12_8 (
    .clk(left_12_8_clk),
    .done(left_12_8_done),
    .in(left_12_8_in),
    .out(left_12_8_out),
    .reset(left_12_8_reset),
    .write_en(left_12_8_write_en)
);
mac_pe pe_12_9 (
    .clk(pe_12_9_clk),
    .done(pe_12_9_done),
    .go(pe_12_9_go),
    .left(pe_12_9_left),
    .mul_ready(pe_12_9_mul_ready),
    .out(pe_12_9_out),
    .reset(pe_12_9_reset),
    .top(pe_12_9_top)
);
std_reg # (
    .WIDTH(32)
) top_12_9 (
    .clk(top_12_9_clk),
    .done(top_12_9_done),
    .in(top_12_9_in),
    .out(top_12_9_out),
    .reset(top_12_9_reset),
    .write_en(top_12_9_write_en)
);
std_reg # (
    .WIDTH(32)
) left_12_9 (
    .clk(left_12_9_clk),
    .done(left_12_9_done),
    .in(left_12_9_in),
    .out(left_12_9_out),
    .reset(left_12_9_reset),
    .write_en(left_12_9_write_en)
);
mac_pe pe_12_10 (
    .clk(pe_12_10_clk),
    .done(pe_12_10_done),
    .go(pe_12_10_go),
    .left(pe_12_10_left),
    .mul_ready(pe_12_10_mul_ready),
    .out(pe_12_10_out),
    .reset(pe_12_10_reset),
    .top(pe_12_10_top)
);
std_reg # (
    .WIDTH(32)
) top_12_10 (
    .clk(top_12_10_clk),
    .done(top_12_10_done),
    .in(top_12_10_in),
    .out(top_12_10_out),
    .reset(top_12_10_reset),
    .write_en(top_12_10_write_en)
);
std_reg # (
    .WIDTH(32)
) left_12_10 (
    .clk(left_12_10_clk),
    .done(left_12_10_done),
    .in(left_12_10_in),
    .out(left_12_10_out),
    .reset(left_12_10_reset),
    .write_en(left_12_10_write_en)
);
mac_pe pe_12_11 (
    .clk(pe_12_11_clk),
    .done(pe_12_11_done),
    .go(pe_12_11_go),
    .left(pe_12_11_left),
    .mul_ready(pe_12_11_mul_ready),
    .out(pe_12_11_out),
    .reset(pe_12_11_reset),
    .top(pe_12_11_top)
);
std_reg # (
    .WIDTH(32)
) top_12_11 (
    .clk(top_12_11_clk),
    .done(top_12_11_done),
    .in(top_12_11_in),
    .out(top_12_11_out),
    .reset(top_12_11_reset),
    .write_en(top_12_11_write_en)
);
std_reg # (
    .WIDTH(32)
) left_12_11 (
    .clk(left_12_11_clk),
    .done(left_12_11_done),
    .in(left_12_11_in),
    .out(left_12_11_out),
    .reset(left_12_11_reset),
    .write_en(left_12_11_write_en)
);
mac_pe pe_12_12 (
    .clk(pe_12_12_clk),
    .done(pe_12_12_done),
    .go(pe_12_12_go),
    .left(pe_12_12_left),
    .mul_ready(pe_12_12_mul_ready),
    .out(pe_12_12_out),
    .reset(pe_12_12_reset),
    .top(pe_12_12_top)
);
std_reg # (
    .WIDTH(32)
) top_12_12 (
    .clk(top_12_12_clk),
    .done(top_12_12_done),
    .in(top_12_12_in),
    .out(top_12_12_out),
    .reset(top_12_12_reset),
    .write_en(top_12_12_write_en)
);
std_reg # (
    .WIDTH(32)
) left_12_12 (
    .clk(left_12_12_clk),
    .done(left_12_12_done),
    .in(left_12_12_in),
    .out(left_12_12_out),
    .reset(left_12_12_reset),
    .write_en(left_12_12_write_en)
);
mac_pe pe_12_13 (
    .clk(pe_12_13_clk),
    .done(pe_12_13_done),
    .go(pe_12_13_go),
    .left(pe_12_13_left),
    .mul_ready(pe_12_13_mul_ready),
    .out(pe_12_13_out),
    .reset(pe_12_13_reset),
    .top(pe_12_13_top)
);
std_reg # (
    .WIDTH(32)
) top_12_13 (
    .clk(top_12_13_clk),
    .done(top_12_13_done),
    .in(top_12_13_in),
    .out(top_12_13_out),
    .reset(top_12_13_reset),
    .write_en(top_12_13_write_en)
);
std_reg # (
    .WIDTH(32)
) left_12_13 (
    .clk(left_12_13_clk),
    .done(left_12_13_done),
    .in(left_12_13_in),
    .out(left_12_13_out),
    .reset(left_12_13_reset),
    .write_en(left_12_13_write_en)
);
mac_pe pe_12_14 (
    .clk(pe_12_14_clk),
    .done(pe_12_14_done),
    .go(pe_12_14_go),
    .left(pe_12_14_left),
    .mul_ready(pe_12_14_mul_ready),
    .out(pe_12_14_out),
    .reset(pe_12_14_reset),
    .top(pe_12_14_top)
);
std_reg # (
    .WIDTH(32)
) top_12_14 (
    .clk(top_12_14_clk),
    .done(top_12_14_done),
    .in(top_12_14_in),
    .out(top_12_14_out),
    .reset(top_12_14_reset),
    .write_en(top_12_14_write_en)
);
std_reg # (
    .WIDTH(32)
) left_12_14 (
    .clk(left_12_14_clk),
    .done(left_12_14_done),
    .in(left_12_14_in),
    .out(left_12_14_out),
    .reset(left_12_14_reset),
    .write_en(left_12_14_write_en)
);
mac_pe pe_12_15 (
    .clk(pe_12_15_clk),
    .done(pe_12_15_done),
    .go(pe_12_15_go),
    .left(pe_12_15_left),
    .mul_ready(pe_12_15_mul_ready),
    .out(pe_12_15_out),
    .reset(pe_12_15_reset),
    .top(pe_12_15_top)
);
std_reg # (
    .WIDTH(32)
) top_12_15 (
    .clk(top_12_15_clk),
    .done(top_12_15_done),
    .in(top_12_15_in),
    .out(top_12_15_out),
    .reset(top_12_15_reset),
    .write_en(top_12_15_write_en)
);
std_reg # (
    .WIDTH(32)
) left_12_15 (
    .clk(left_12_15_clk),
    .done(left_12_15_done),
    .in(left_12_15_in),
    .out(left_12_15_out),
    .reset(left_12_15_reset),
    .write_en(left_12_15_write_en)
);
mac_pe pe_13_0 (
    .clk(pe_13_0_clk),
    .done(pe_13_0_done),
    .go(pe_13_0_go),
    .left(pe_13_0_left),
    .mul_ready(pe_13_0_mul_ready),
    .out(pe_13_0_out),
    .reset(pe_13_0_reset),
    .top(pe_13_0_top)
);
std_reg # (
    .WIDTH(32)
) top_13_0 (
    .clk(top_13_0_clk),
    .done(top_13_0_done),
    .in(top_13_0_in),
    .out(top_13_0_out),
    .reset(top_13_0_reset),
    .write_en(top_13_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_13_0 (
    .clk(left_13_0_clk),
    .done(left_13_0_done),
    .in(left_13_0_in),
    .out(left_13_0_out),
    .reset(left_13_0_reset),
    .write_en(left_13_0_write_en)
);
mac_pe pe_13_1 (
    .clk(pe_13_1_clk),
    .done(pe_13_1_done),
    .go(pe_13_1_go),
    .left(pe_13_1_left),
    .mul_ready(pe_13_1_mul_ready),
    .out(pe_13_1_out),
    .reset(pe_13_1_reset),
    .top(pe_13_1_top)
);
std_reg # (
    .WIDTH(32)
) top_13_1 (
    .clk(top_13_1_clk),
    .done(top_13_1_done),
    .in(top_13_1_in),
    .out(top_13_1_out),
    .reset(top_13_1_reset),
    .write_en(top_13_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_13_1 (
    .clk(left_13_1_clk),
    .done(left_13_1_done),
    .in(left_13_1_in),
    .out(left_13_1_out),
    .reset(left_13_1_reset),
    .write_en(left_13_1_write_en)
);
mac_pe pe_13_2 (
    .clk(pe_13_2_clk),
    .done(pe_13_2_done),
    .go(pe_13_2_go),
    .left(pe_13_2_left),
    .mul_ready(pe_13_2_mul_ready),
    .out(pe_13_2_out),
    .reset(pe_13_2_reset),
    .top(pe_13_2_top)
);
std_reg # (
    .WIDTH(32)
) top_13_2 (
    .clk(top_13_2_clk),
    .done(top_13_2_done),
    .in(top_13_2_in),
    .out(top_13_2_out),
    .reset(top_13_2_reset),
    .write_en(top_13_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_13_2 (
    .clk(left_13_2_clk),
    .done(left_13_2_done),
    .in(left_13_2_in),
    .out(left_13_2_out),
    .reset(left_13_2_reset),
    .write_en(left_13_2_write_en)
);
mac_pe pe_13_3 (
    .clk(pe_13_3_clk),
    .done(pe_13_3_done),
    .go(pe_13_3_go),
    .left(pe_13_3_left),
    .mul_ready(pe_13_3_mul_ready),
    .out(pe_13_3_out),
    .reset(pe_13_3_reset),
    .top(pe_13_3_top)
);
std_reg # (
    .WIDTH(32)
) top_13_3 (
    .clk(top_13_3_clk),
    .done(top_13_3_done),
    .in(top_13_3_in),
    .out(top_13_3_out),
    .reset(top_13_3_reset),
    .write_en(top_13_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_13_3 (
    .clk(left_13_3_clk),
    .done(left_13_3_done),
    .in(left_13_3_in),
    .out(left_13_3_out),
    .reset(left_13_3_reset),
    .write_en(left_13_3_write_en)
);
mac_pe pe_13_4 (
    .clk(pe_13_4_clk),
    .done(pe_13_4_done),
    .go(pe_13_4_go),
    .left(pe_13_4_left),
    .mul_ready(pe_13_4_mul_ready),
    .out(pe_13_4_out),
    .reset(pe_13_4_reset),
    .top(pe_13_4_top)
);
std_reg # (
    .WIDTH(32)
) top_13_4 (
    .clk(top_13_4_clk),
    .done(top_13_4_done),
    .in(top_13_4_in),
    .out(top_13_4_out),
    .reset(top_13_4_reset),
    .write_en(top_13_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_13_4 (
    .clk(left_13_4_clk),
    .done(left_13_4_done),
    .in(left_13_4_in),
    .out(left_13_4_out),
    .reset(left_13_4_reset),
    .write_en(left_13_4_write_en)
);
mac_pe pe_13_5 (
    .clk(pe_13_5_clk),
    .done(pe_13_5_done),
    .go(pe_13_5_go),
    .left(pe_13_5_left),
    .mul_ready(pe_13_5_mul_ready),
    .out(pe_13_5_out),
    .reset(pe_13_5_reset),
    .top(pe_13_5_top)
);
std_reg # (
    .WIDTH(32)
) top_13_5 (
    .clk(top_13_5_clk),
    .done(top_13_5_done),
    .in(top_13_5_in),
    .out(top_13_5_out),
    .reset(top_13_5_reset),
    .write_en(top_13_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_13_5 (
    .clk(left_13_5_clk),
    .done(left_13_5_done),
    .in(left_13_5_in),
    .out(left_13_5_out),
    .reset(left_13_5_reset),
    .write_en(left_13_5_write_en)
);
mac_pe pe_13_6 (
    .clk(pe_13_6_clk),
    .done(pe_13_6_done),
    .go(pe_13_6_go),
    .left(pe_13_6_left),
    .mul_ready(pe_13_6_mul_ready),
    .out(pe_13_6_out),
    .reset(pe_13_6_reset),
    .top(pe_13_6_top)
);
std_reg # (
    .WIDTH(32)
) top_13_6 (
    .clk(top_13_6_clk),
    .done(top_13_6_done),
    .in(top_13_6_in),
    .out(top_13_6_out),
    .reset(top_13_6_reset),
    .write_en(top_13_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_13_6 (
    .clk(left_13_6_clk),
    .done(left_13_6_done),
    .in(left_13_6_in),
    .out(left_13_6_out),
    .reset(left_13_6_reset),
    .write_en(left_13_6_write_en)
);
mac_pe pe_13_7 (
    .clk(pe_13_7_clk),
    .done(pe_13_7_done),
    .go(pe_13_7_go),
    .left(pe_13_7_left),
    .mul_ready(pe_13_7_mul_ready),
    .out(pe_13_7_out),
    .reset(pe_13_7_reset),
    .top(pe_13_7_top)
);
std_reg # (
    .WIDTH(32)
) top_13_7 (
    .clk(top_13_7_clk),
    .done(top_13_7_done),
    .in(top_13_7_in),
    .out(top_13_7_out),
    .reset(top_13_7_reset),
    .write_en(top_13_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_13_7 (
    .clk(left_13_7_clk),
    .done(left_13_7_done),
    .in(left_13_7_in),
    .out(left_13_7_out),
    .reset(left_13_7_reset),
    .write_en(left_13_7_write_en)
);
mac_pe pe_13_8 (
    .clk(pe_13_8_clk),
    .done(pe_13_8_done),
    .go(pe_13_8_go),
    .left(pe_13_8_left),
    .mul_ready(pe_13_8_mul_ready),
    .out(pe_13_8_out),
    .reset(pe_13_8_reset),
    .top(pe_13_8_top)
);
std_reg # (
    .WIDTH(32)
) top_13_8 (
    .clk(top_13_8_clk),
    .done(top_13_8_done),
    .in(top_13_8_in),
    .out(top_13_8_out),
    .reset(top_13_8_reset),
    .write_en(top_13_8_write_en)
);
std_reg # (
    .WIDTH(32)
) left_13_8 (
    .clk(left_13_8_clk),
    .done(left_13_8_done),
    .in(left_13_8_in),
    .out(left_13_8_out),
    .reset(left_13_8_reset),
    .write_en(left_13_8_write_en)
);
mac_pe pe_13_9 (
    .clk(pe_13_9_clk),
    .done(pe_13_9_done),
    .go(pe_13_9_go),
    .left(pe_13_9_left),
    .mul_ready(pe_13_9_mul_ready),
    .out(pe_13_9_out),
    .reset(pe_13_9_reset),
    .top(pe_13_9_top)
);
std_reg # (
    .WIDTH(32)
) top_13_9 (
    .clk(top_13_9_clk),
    .done(top_13_9_done),
    .in(top_13_9_in),
    .out(top_13_9_out),
    .reset(top_13_9_reset),
    .write_en(top_13_9_write_en)
);
std_reg # (
    .WIDTH(32)
) left_13_9 (
    .clk(left_13_9_clk),
    .done(left_13_9_done),
    .in(left_13_9_in),
    .out(left_13_9_out),
    .reset(left_13_9_reset),
    .write_en(left_13_9_write_en)
);
mac_pe pe_13_10 (
    .clk(pe_13_10_clk),
    .done(pe_13_10_done),
    .go(pe_13_10_go),
    .left(pe_13_10_left),
    .mul_ready(pe_13_10_mul_ready),
    .out(pe_13_10_out),
    .reset(pe_13_10_reset),
    .top(pe_13_10_top)
);
std_reg # (
    .WIDTH(32)
) top_13_10 (
    .clk(top_13_10_clk),
    .done(top_13_10_done),
    .in(top_13_10_in),
    .out(top_13_10_out),
    .reset(top_13_10_reset),
    .write_en(top_13_10_write_en)
);
std_reg # (
    .WIDTH(32)
) left_13_10 (
    .clk(left_13_10_clk),
    .done(left_13_10_done),
    .in(left_13_10_in),
    .out(left_13_10_out),
    .reset(left_13_10_reset),
    .write_en(left_13_10_write_en)
);
mac_pe pe_13_11 (
    .clk(pe_13_11_clk),
    .done(pe_13_11_done),
    .go(pe_13_11_go),
    .left(pe_13_11_left),
    .mul_ready(pe_13_11_mul_ready),
    .out(pe_13_11_out),
    .reset(pe_13_11_reset),
    .top(pe_13_11_top)
);
std_reg # (
    .WIDTH(32)
) top_13_11 (
    .clk(top_13_11_clk),
    .done(top_13_11_done),
    .in(top_13_11_in),
    .out(top_13_11_out),
    .reset(top_13_11_reset),
    .write_en(top_13_11_write_en)
);
std_reg # (
    .WIDTH(32)
) left_13_11 (
    .clk(left_13_11_clk),
    .done(left_13_11_done),
    .in(left_13_11_in),
    .out(left_13_11_out),
    .reset(left_13_11_reset),
    .write_en(left_13_11_write_en)
);
mac_pe pe_13_12 (
    .clk(pe_13_12_clk),
    .done(pe_13_12_done),
    .go(pe_13_12_go),
    .left(pe_13_12_left),
    .mul_ready(pe_13_12_mul_ready),
    .out(pe_13_12_out),
    .reset(pe_13_12_reset),
    .top(pe_13_12_top)
);
std_reg # (
    .WIDTH(32)
) top_13_12 (
    .clk(top_13_12_clk),
    .done(top_13_12_done),
    .in(top_13_12_in),
    .out(top_13_12_out),
    .reset(top_13_12_reset),
    .write_en(top_13_12_write_en)
);
std_reg # (
    .WIDTH(32)
) left_13_12 (
    .clk(left_13_12_clk),
    .done(left_13_12_done),
    .in(left_13_12_in),
    .out(left_13_12_out),
    .reset(left_13_12_reset),
    .write_en(left_13_12_write_en)
);
mac_pe pe_13_13 (
    .clk(pe_13_13_clk),
    .done(pe_13_13_done),
    .go(pe_13_13_go),
    .left(pe_13_13_left),
    .mul_ready(pe_13_13_mul_ready),
    .out(pe_13_13_out),
    .reset(pe_13_13_reset),
    .top(pe_13_13_top)
);
std_reg # (
    .WIDTH(32)
) top_13_13 (
    .clk(top_13_13_clk),
    .done(top_13_13_done),
    .in(top_13_13_in),
    .out(top_13_13_out),
    .reset(top_13_13_reset),
    .write_en(top_13_13_write_en)
);
std_reg # (
    .WIDTH(32)
) left_13_13 (
    .clk(left_13_13_clk),
    .done(left_13_13_done),
    .in(left_13_13_in),
    .out(left_13_13_out),
    .reset(left_13_13_reset),
    .write_en(left_13_13_write_en)
);
mac_pe pe_13_14 (
    .clk(pe_13_14_clk),
    .done(pe_13_14_done),
    .go(pe_13_14_go),
    .left(pe_13_14_left),
    .mul_ready(pe_13_14_mul_ready),
    .out(pe_13_14_out),
    .reset(pe_13_14_reset),
    .top(pe_13_14_top)
);
std_reg # (
    .WIDTH(32)
) top_13_14 (
    .clk(top_13_14_clk),
    .done(top_13_14_done),
    .in(top_13_14_in),
    .out(top_13_14_out),
    .reset(top_13_14_reset),
    .write_en(top_13_14_write_en)
);
std_reg # (
    .WIDTH(32)
) left_13_14 (
    .clk(left_13_14_clk),
    .done(left_13_14_done),
    .in(left_13_14_in),
    .out(left_13_14_out),
    .reset(left_13_14_reset),
    .write_en(left_13_14_write_en)
);
mac_pe pe_13_15 (
    .clk(pe_13_15_clk),
    .done(pe_13_15_done),
    .go(pe_13_15_go),
    .left(pe_13_15_left),
    .mul_ready(pe_13_15_mul_ready),
    .out(pe_13_15_out),
    .reset(pe_13_15_reset),
    .top(pe_13_15_top)
);
std_reg # (
    .WIDTH(32)
) top_13_15 (
    .clk(top_13_15_clk),
    .done(top_13_15_done),
    .in(top_13_15_in),
    .out(top_13_15_out),
    .reset(top_13_15_reset),
    .write_en(top_13_15_write_en)
);
std_reg # (
    .WIDTH(32)
) left_13_15 (
    .clk(left_13_15_clk),
    .done(left_13_15_done),
    .in(left_13_15_in),
    .out(left_13_15_out),
    .reset(left_13_15_reset),
    .write_en(left_13_15_write_en)
);
mac_pe pe_14_0 (
    .clk(pe_14_0_clk),
    .done(pe_14_0_done),
    .go(pe_14_0_go),
    .left(pe_14_0_left),
    .mul_ready(pe_14_0_mul_ready),
    .out(pe_14_0_out),
    .reset(pe_14_0_reset),
    .top(pe_14_0_top)
);
std_reg # (
    .WIDTH(32)
) top_14_0 (
    .clk(top_14_0_clk),
    .done(top_14_0_done),
    .in(top_14_0_in),
    .out(top_14_0_out),
    .reset(top_14_0_reset),
    .write_en(top_14_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_14_0 (
    .clk(left_14_0_clk),
    .done(left_14_0_done),
    .in(left_14_0_in),
    .out(left_14_0_out),
    .reset(left_14_0_reset),
    .write_en(left_14_0_write_en)
);
mac_pe pe_14_1 (
    .clk(pe_14_1_clk),
    .done(pe_14_1_done),
    .go(pe_14_1_go),
    .left(pe_14_1_left),
    .mul_ready(pe_14_1_mul_ready),
    .out(pe_14_1_out),
    .reset(pe_14_1_reset),
    .top(pe_14_1_top)
);
std_reg # (
    .WIDTH(32)
) top_14_1 (
    .clk(top_14_1_clk),
    .done(top_14_1_done),
    .in(top_14_1_in),
    .out(top_14_1_out),
    .reset(top_14_1_reset),
    .write_en(top_14_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_14_1 (
    .clk(left_14_1_clk),
    .done(left_14_1_done),
    .in(left_14_1_in),
    .out(left_14_1_out),
    .reset(left_14_1_reset),
    .write_en(left_14_1_write_en)
);
mac_pe pe_14_2 (
    .clk(pe_14_2_clk),
    .done(pe_14_2_done),
    .go(pe_14_2_go),
    .left(pe_14_2_left),
    .mul_ready(pe_14_2_mul_ready),
    .out(pe_14_2_out),
    .reset(pe_14_2_reset),
    .top(pe_14_2_top)
);
std_reg # (
    .WIDTH(32)
) top_14_2 (
    .clk(top_14_2_clk),
    .done(top_14_2_done),
    .in(top_14_2_in),
    .out(top_14_2_out),
    .reset(top_14_2_reset),
    .write_en(top_14_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_14_2 (
    .clk(left_14_2_clk),
    .done(left_14_2_done),
    .in(left_14_2_in),
    .out(left_14_2_out),
    .reset(left_14_2_reset),
    .write_en(left_14_2_write_en)
);
mac_pe pe_14_3 (
    .clk(pe_14_3_clk),
    .done(pe_14_3_done),
    .go(pe_14_3_go),
    .left(pe_14_3_left),
    .mul_ready(pe_14_3_mul_ready),
    .out(pe_14_3_out),
    .reset(pe_14_3_reset),
    .top(pe_14_3_top)
);
std_reg # (
    .WIDTH(32)
) top_14_3 (
    .clk(top_14_3_clk),
    .done(top_14_3_done),
    .in(top_14_3_in),
    .out(top_14_3_out),
    .reset(top_14_3_reset),
    .write_en(top_14_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_14_3 (
    .clk(left_14_3_clk),
    .done(left_14_3_done),
    .in(left_14_3_in),
    .out(left_14_3_out),
    .reset(left_14_3_reset),
    .write_en(left_14_3_write_en)
);
mac_pe pe_14_4 (
    .clk(pe_14_4_clk),
    .done(pe_14_4_done),
    .go(pe_14_4_go),
    .left(pe_14_4_left),
    .mul_ready(pe_14_4_mul_ready),
    .out(pe_14_4_out),
    .reset(pe_14_4_reset),
    .top(pe_14_4_top)
);
std_reg # (
    .WIDTH(32)
) top_14_4 (
    .clk(top_14_4_clk),
    .done(top_14_4_done),
    .in(top_14_4_in),
    .out(top_14_4_out),
    .reset(top_14_4_reset),
    .write_en(top_14_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_14_4 (
    .clk(left_14_4_clk),
    .done(left_14_4_done),
    .in(left_14_4_in),
    .out(left_14_4_out),
    .reset(left_14_4_reset),
    .write_en(left_14_4_write_en)
);
mac_pe pe_14_5 (
    .clk(pe_14_5_clk),
    .done(pe_14_5_done),
    .go(pe_14_5_go),
    .left(pe_14_5_left),
    .mul_ready(pe_14_5_mul_ready),
    .out(pe_14_5_out),
    .reset(pe_14_5_reset),
    .top(pe_14_5_top)
);
std_reg # (
    .WIDTH(32)
) top_14_5 (
    .clk(top_14_5_clk),
    .done(top_14_5_done),
    .in(top_14_5_in),
    .out(top_14_5_out),
    .reset(top_14_5_reset),
    .write_en(top_14_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_14_5 (
    .clk(left_14_5_clk),
    .done(left_14_5_done),
    .in(left_14_5_in),
    .out(left_14_5_out),
    .reset(left_14_5_reset),
    .write_en(left_14_5_write_en)
);
mac_pe pe_14_6 (
    .clk(pe_14_6_clk),
    .done(pe_14_6_done),
    .go(pe_14_6_go),
    .left(pe_14_6_left),
    .mul_ready(pe_14_6_mul_ready),
    .out(pe_14_6_out),
    .reset(pe_14_6_reset),
    .top(pe_14_6_top)
);
std_reg # (
    .WIDTH(32)
) top_14_6 (
    .clk(top_14_6_clk),
    .done(top_14_6_done),
    .in(top_14_6_in),
    .out(top_14_6_out),
    .reset(top_14_6_reset),
    .write_en(top_14_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_14_6 (
    .clk(left_14_6_clk),
    .done(left_14_6_done),
    .in(left_14_6_in),
    .out(left_14_6_out),
    .reset(left_14_6_reset),
    .write_en(left_14_6_write_en)
);
mac_pe pe_14_7 (
    .clk(pe_14_7_clk),
    .done(pe_14_7_done),
    .go(pe_14_7_go),
    .left(pe_14_7_left),
    .mul_ready(pe_14_7_mul_ready),
    .out(pe_14_7_out),
    .reset(pe_14_7_reset),
    .top(pe_14_7_top)
);
std_reg # (
    .WIDTH(32)
) top_14_7 (
    .clk(top_14_7_clk),
    .done(top_14_7_done),
    .in(top_14_7_in),
    .out(top_14_7_out),
    .reset(top_14_7_reset),
    .write_en(top_14_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_14_7 (
    .clk(left_14_7_clk),
    .done(left_14_7_done),
    .in(left_14_7_in),
    .out(left_14_7_out),
    .reset(left_14_7_reset),
    .write_en(left_14_7_write_en)
);
mac_pe pe_14_8 (
    .clk(pe_14_8_clk),
    .done(pe_14_8_done),
    .go(pe_14_8_go),
    .left(pe_14_8_left),
    .mul_ready(pe_14_8_mul_ready),
    .out(pe_14_8_out),
    .reset(pe_14_8_reset),
    .top(pe_14_8_top)
);
std_reg # (
    .WIDTH(32)
) top_14_8 (
    .clk(top_14_8_clk),
    .done(top_14_8_done),
    .in(top_14_8_in),
    .out(top_14_8_out),
    .reset(top_14_8_reset),
    .write_en(top_14_8_write_en)
);
std_reg # (
    .WIDTH(32)
) left_14_8 (
    .clk(left_14_8_clk),
    .done(left_14_8_done),
    .in(left_14_8_in),
    .out(left_14_8_out),
    .reset(left_14_8_reset),
    .write_en(left_14_8_write_en)
);
mac_pe pe_14_9 (
    .clk(pe_14_9_clk),
    .done(pe_14_9_done),
    .go(pe_14_9_go),
    .left(pe_14_9_left),
    .mul_ready(pe_14_9_mul_ready),
    .out(pe_14_9_out),
    .reset(pe_14_9_reset),
    .top(pe_14_9_top)
);
std_reg # (
    .WIDTH(32)
) top_14_9 (
    .clk(top_14_9_clk),
    .done(top_14_9_done),
    .in(top_14_9_in),
    .out(top_14_9_out),
    .reset(top_14_9_reset),
    .write_en(top_14_9_write_en)
);
std_reg # (
    .WIDTH(32)
) left_14_9 (
    .clk(left_14_9_clk),
    .done(left_14_9_done),
    .in(left_14_9_in),
    .out(left_14_9_out),
    .reset(left_14_9_reset),
    .write_en(left_14_9_write_en)
);
mac_pe pe_14_10 (
    .clk(pe_14_10_clk),
    .done(pe_14_10_done),
    .go(pe_14_10_go),
    .left(pe_14_10_left),
    .mul_ready(pe_14_10_mul_ready),
    .out(pe_14_10_out),
    .reset(pe_14_10_reset),
    .top(pe_14_10_top)
);
std_reg # (
    .WIDTH(32)
) top_14_10 (
    .clk(top_14_10_clk),
    .done(top_14_10_done),
    .in(top_14_10_in),
    .out(top_14_10_out),
    .reset(top_14_10_reset),
    .write_en(top_14_10_write_en)
);
std_reg # (
    .WIDTH(32)
) left_14_10 (
    .clk(left_14_10_clk),
    .done(left_14_10_done),
    .in(left_14_10_in),
    .out(left_14_10_out),
    .reset(left_14_10_reset),
    .write_en(left_14_10_write_en)
);
mac_pe pe_14_11 (
    .clk(pe_14_11_clk),
    .done(pe_14_11_done),
    .go(pe_14_11_go),
    .left(pe_14_11_left),
    .mul_ready(pe_14_11_mul_ready),
    .out(pe_14_11_out),
    .reset(pe_14_11_reset),
    .top(pe_14_11_top)
);
std_reg # (
    .WIDTH(32)
) top_14_11 (
    .clk(top_14_11_clk),
    .done(top_14_11_done),
    .in(top_14_11_in),
    .out(top_14_11_out),
    .reset(top_14_11_reset),
    .write_en(top_14_11_write_en)
);
std_reg # (
    .WIDTH(32)
) left_14_11 (
    .clk(left_14_11_clk),
    .done(left_14_11_done),
    .in(left_14_11_in),
    .out(left_14_11_out),
    .reset(left_14_11_reset),
    .write_en(left_14_11_write_en)
);
mac_pe pe_14_12 (
    .clk(pe_14_12_clk),
    .done(pe_14_12_done),
    .go(pe_14_12_go),
    .left(pe_14_12_left),
    .mul_ready(pe_14_12_mul_ready),
    .out(pe_14_12_out),
    .reset(pe_14_12_reset),
    .top(pe_14_12_top)
);
std_reg # (
    .WIDTH(32)
) top_14_12 (
    .clk(top_14_12_clk),
    .done(top_14_12_done),
    .in(top_14_12_in),
    .out(top_14_12_out),
    .reset(top_14_12_reset),
    .write_en(top_14_12_write_en)
);
std_reg # (
    .WIDTH(32)
) left_14_12 (
    .clk(left_14_12_clk),
    .done(left_14_12_done),
    .in(left_14_12_in),
    .out(left_14_12_out),
    .reset(left_14_12_reset),
    .write_en(left_14_12_write_en)
);
mac_pe pe_14_13 (
    .clk(pe_14_13_clk),
    .done(pe_14_13_done),
    .go(pe_14_13_go),
    .left(pe_14_13_left),
    .mul_ready(pe_14_13_mul_ready),
    .out(pe_14_13_out),
    .reset(pe_14_13_reset),
    .top(pe_14_13_top)
);
std_reg # (
    .WIDTH(32)
) top_14_13 (
    .clk(top_14_13_clk),
    .done(top_14_13_done),
    .in(top_14_13_in),
    .out(top_14_13_out),
    .reset(top_14_13_reset),
    .write_en(top_14_13_write_en)
);
std_reg # (
    .WIDTH(32)
) left_14_13 (
    .clk(left_14_13_clk),
    .done(left_14_13_done),
    .in(left_14_13_in),
    .out(left_14_13_out),
    .reset(left_14_13_reset),
    .write_en(left_14_13_write_en)
);
mac_pe pe_14_14 (
    .clk(pe_14_14_clk),
    .done(pe_14_14_done),
    .go(pe_14_14_go),
    .left(pe_14_14_left),
    .mul_ready(pe_14_14_mul_ready),
    .out(pe_14_14_out),
    .reset(pe_14_14_reset),
    .top(pe_14_14_top)
);
std_reg # (
    .WIDTH(32)
) top_14_14 (
    .clk(top_14_14_clk),
    .done(top_14_14_done),
    .in(top_14_14_in),
    .out(top_14_14_out),
    .reset(top_14_14_reset),
    .write_en(top_14_14_write_en)
);
std_reg # (
    .WIDTH(32)
) left_14_14 (
    .clk(left_14_14_clk),
    .done(left_14_14_done),
    .in(left_14_14_in),
    .out(left_14_14_out),
    .reset(left_14_14_reset),
    .write_en(left_14_14_write_en)
);
mac_pe pe_14_15 (
    .clk(pe_14_15_clk),
    .done(pe_14_15_done),
    .go(pe_14_15_go),
    .left(pe_14_15_left),
    .mul_ready(pe_14_15_mul_ready),
    .out(pe_14_15_out),
    .reset(pe_14_15_reset),
    .top(pe_14_15_top)
);
std_reg # (
    .WIDTH(32)
) top_14_15 (
    .clk(top_14_15_clk),
    .done(top_14_15_done),
    .in(top_14_15_in),
    .out(top_14_15_out),
    .reset(top_14_15_reset),
    .write_en(top_14_15_write_en)
);
std_reg # (
    .WIDTH(32)
) left_14_15 (
    .clk(left_14_15_clk),
    .done(left_14_15_done),
    .in(left_14_15_in),
    .out(left_14_15_out),
    .reset(left_14_15_reset),
    .write_en(left_14_15_write_en)
);
mac_pe pe_15_0 (
    .clk(pe_15_0_clk),
    .done(pe_15_0_done),
    .go(pe_15_0_go),
    .left(pe_15_0_left),
    .mul_ready(pe_15_0_mul_ready),
    .out(pe_15_0_out),
    .reset(pe_15_0_reset),
    .top(pe_15_0_top)
);
std_reg # (
    .WIDTH(32)
) top_15_0 (
    .clk(top_15_0_clk),
    .done(top_15_0_done),
    .in(top_15_0_in),
    .out(top_15_0_out),
    .reset(top_15_0_reset),
    .write_en(top_15_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_15_0 (
    .clk(left_15_0_clk),
    .done(left_15_0_done),
    .in(left_15_0_in),
    .out(left_15_0_out),
    .reset(left_15_0_reset),
    .write_en(left_15_0_write_en)
);
mac_pe pe_15_1 (
    .clk(pe_15_1_clk),
    .done(pe_15_1_done),
    .go(pe_15_1_go),
    .left(pe_15_1_left),
    .mul_ready(pe_15_1_mul_ready),
    .out(pe_15_1_out),
    .reset(pe_15_1_reset),
    .top(pe_15_1_top)
);
std_reg # (
    .WIDTH(32)
) top_15_1 (
    .clk(top_15_1_clk),
    .done(top_15_1_done),
    .in(top_15_1_in),
    .out(top_15_1_out),
    .reset(top_15_1_reset),
    .write_en(top_15_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_15_1 (
    .clk(left_15_1_clk),
    .done(left_15_1_done),
    .in(left_15_1_in),
    .out(left_15_1_out),
    .reset(left_15_1_reset),
    .write_en(left_15_1_write_en)
);
mac_pe pe_15_2 (
    .clk(pe_15_2_clk),
    .done(pe_15_2_done),
    .go(pe_15_2_go),
    .left(pe_15_2_left),
    .mul_ready(pe_15_2_mul_ready),
    .out(pe_15_2_out),
    .reset(pe_15_2_reset),
    .top(pe_15_2_top)
);
std_reg # (
    .WIDTH(32)
) top_15_2 (
    .clk(top_15_2_clk),
    .done(top_15_2_done),
    .in(top_15_2_in),
    .out(top_15_2_out),
    .reset(top_15_2_reset),
    .write_en(top_15_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_15_2 (
    .clk(left_15_2_clk),
    .done(left_15_2_done),
    .in(left_15_2_in),
    .out(left_15_2_out),
    .reset(left_15_2_reset),
    .write_en(left_15_2_write_en)
);
mac_pe pe_15_3 (
    .clk(pe_15_3_clk),
    .done(pe_15_3_done),
    .go(pe_15_3_go),
    .left(pe_15_3_left),
    .mul_ready(pe_15_3_mul_ready),
    .out(pe_15_3_out),
    .reset(pe_15_3_reset),
    .top(pe_15_3_top)
);
std_reg # (
    .WIDTH(32)
) top_15_3 (
    .clk(top_15_3_clk),
    .done(top_15_3_done),
    .in(top_15_3_in),
    .out(top_15_3_out),
    .reset(top_15_3_reset),
    .write_en(top_15_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_15_3 (
    .clk(left_15_3_clk),
    .done(left_15_3_done),
    .in(left_15_3_in),
    .out(left_15_3_out),
    .reset(left_15_3_reset),
    .write_en(left_15_3_write_en)
);
mac_pe pe_15_4 (
    .clk(pe_15_4_clk),
    .done(pe_15_4_done),
    .go(pe_15_4_go),
    .left(pe_15_4_left),
    .mul_ready(pe_15_4_mul_ready),
    .out(pe_15_4_out),
    .reset(pe_15_4_reset),
    .top(pe_15_4_top)
);
std_reg # (
    .WIDTH(32)
) top_15_4 (
    .clk(top_15_4_clk),
    .done(top_15_4_done),
    .in(top_15_4_in),
    .out(top_15_4_out),
    .reset(top_15_4_reset),
    .write_en(top_15_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_15_4 (
    .clk(left_15_4_clk),
    .done(left_15_4_done),
    .in(left_15_4_in),
    .out(left_15_4_out),
    .reset(left_15_4_reset),
    .write_en(left_15_4_write_en)
);
mac_pe pe_15_5 (
    .clk(pe_15_5_clk),
    .done(pe_15_5_done),
    .go(pe_15_5_go),
    .left(pe_15_5_left),
    .mul_ready(pe_15_5_mul_ready),
    .out(pe_15_5_out),
    .reset(pe_15_5_reset),
    .top(pe_15_5_top)
);
std_reg # (
    .WIDTH(32)
) top_15_5 (
    .clk(top_15_5_clk),
    .done(top_15_5_done),
    .in(top_15_5_in),
    .out(top_15_5_out),
    .reset(top_15_5_reset),
    .write_en(top_15_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_15_5 (
    .clk(left_15_5_clk),
    .done(left_15_5_done),
    .in(left_15_5_in),
    .out(left_15_5_out),
    .reset(left_15_5_reset),
    .write_en(left_15_5_write_en)
);
mac_pe pe_15_6 (
    .clk(pe_15_6_clk),
    .done(pe_15_6_done),
    .go(pe_15_6_go),
    .left(pe_15_6_left),
    .mul_ready(pe_15_6_mul_ready),
    .out(pe_15_6_out),
    .reset(pe_15_6_reset),
    .top(pe_15_6_top)
);
std_reg # (
    .WIDTH(32)
) top_15_6 (
    .clk(top_15_6_clk),
    .done(top_15_6_done),
    .in(top_15_6_in),
    .out(top_15_6_out),
    .reset(top_15_6_reset),
    .write_en(top_15_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_15_6 (
    .clk(left_15_6_clk),
    .done(left_15_6_done),
    .in(left_15_6_in),
    .out(left_15_6_out),
    .reset(left_15_6_reset),
    .write_en(left_15_6_write_en)
);
mac_pe pe_15_7 (
    .clk(pe_15_7_clk),
    .done(pe_15_7_done),
    .go(pe_15_7_go),
    .left(pe_15_7_left),
    .mul_ready(pe_15_7_mul_ready),
    .out(pe_15_7_out),
    .reset(pe_15_7_reset),
    .top(pe_15_7_top)
);
std_reg # (
    .WIDTH(32)
) top_15_7 (
    .clk(top_15_7_clk),
    .done(top_15_7_done),
    .in(top_15_7_in),
    .out(top_15_7_out),
    .reset(top_15_7_reset),
    .write_en(top_15_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_15_7 (
    .clk(left_15_7_clk),
    .done(left_15_7_done),
    .in(left_15_7_in),
    .out(left_15_7_out),
    .reset(left_15_7_reset),
    .write_en(left_15_7_write_en)
);
mac_pe pe_15_8 (
    .clk(pe_15_8_clk),
    .done(pe_15_8_done),
    .go(pe_15_8_go),
    .left(pe_15_8_left),
    .mul_ready(pe_15_8_mul_ready),
    .out(pe_15_8_out),
    .reset(pe_15_8_reset),
    .top(pe_15_8_top)
);
std_reg # (
    .WIDTH(32)
) top_15_8 (
    .clk(top_15_8_clk),
    .done(top_15_8_done),
    .in(top_15_8_in),
    .out(top_15_8_out),
    .reset(top_15_8_reset),
    .write_en(top_15_8_write_en)
);
std_reg # (
    .WIDTH(32)
) left_15_8 (
    .clk(left_15_8_clk),
    .done(left_15_8_done),
    .in(left_15_8_in),
    .out(left_15_8_out),
    .reset(left_15_8_reset),
    .write_en(left_15_8_write_en)
);
mac_pe pe_15_9 (
    .clk(pe_15_9_clk),
    .done(pe_15_9_done),
    .go(pe_15_9_go),
    .left(pe_15_9_left),
    .mul_ready(pe_15_9_mul_ready),
    .out(pe_15_9_out),
    .reset(pe_15_9_reset),
    .top(pe_15_9_top)
);
std_reg # (
    .WIDTH(32)
) top_15_9 (
    .clk(top_15_9_clk),
    .done(top_15_9_done),
    .in(top_15_9_in),
    .out(top_15_9_out),
    .reset(top_15_9_reset),
    .write_en(top_15_9_write_en)
);
std_reg # (
    .WIDTH(32)
) left_15_9 (
    .clk(left_15_9_clk),
    .done(left_15_9_done),
    .in(left_15_9_in),
    .out(left_15_9_out),
    .reset(left_15_9_reset),
    .write_en(left_15_9_write_en)
);
mac_pe pe_15_10 (
    .clk(pe_15_10_clk),
    .done(pe_15_10_done),
    .go(pe_15_10_go),
    .left(pe_15_10_left),
    .mul_ready(pe_15_10_mul_ready),
    .out(pe_15_10_out),
    .reset(pe_15_10_reset),
    .top(pe_15_10_top)
);
std_reg # (
    .WIDTH(32)
) top_15_10 (
    .clk(top_15_10_clk),
    .done(top_15_10_done),
    .in(top_15_10_in),
    .out(top_15_10_out),
    .reset(top_15_10_reset),
    .write_en(top_15_10_write_en)
);
std_reg # (
    .WIDTH(32)
) left_15_10 (
    .clk(left_15_10_clk),
    .done(left_15_10_done),
    .in(left_15_10_in),
    .out(left_15_10_out),
    .reset(left_15_10_reset),
    .write_en(left_15_10_write_en)
);
mac_pe pe_15_11 (
    .clk(pe_15_11_clk),
    .done(pe_15_11_done),
    .go(pe_15_11_go),
    .left(pe_15_11_left),
    .mul_ready(pe_15_11_mul_ready),
    .out(pe_15_11_out),
    .reset(pe_15_11_reset),
    .top(pe_15_11_top)
);
std_reg # (
    .WIDTH(32)
) top_15_11 (
    .clk(top_15_11_clk),
    .done(top_15_11_done),
    .in(top_15_11_in),
    .out(top_15_11_out),
    .reset(top_15_11_reset),
    .write_en(top_15_11_write_en)
);
std_reg # (
    .WIDTH(32)
) left_15_11 (
    .clk(left_15_11_clk),
    .done(left_15_11_done),
    .in(left_15_11_in),
    .out(left_15_11_out),
    .reset(left_15_11_reset),
    .write_en(left_15_11_write_en)
);
mac_pe pe_15_12 (
    .clk(pe_15_12_clk),
    .done(pe_15_12_done),
    .go(pe_15_12_go),
    .left(pe_15_12_left),
    .mul_ready(pe_15_12_mul_ready),
    .out(pe_15_12_out),
    .reset(pe_15_12_reset),
    .top(pe_15_12_top)
);
std_reg # (
    .WIDTH(32)
) top_15_12 (
    .clk(top_15_12_clk),
    .done(top_15_12_done),
    .in(top_15_12_in),
    .out(top_15_12_out),
    .reset(top_15_12_reset),
    .write_en(top_15_12_write_en)
);
std_reg # (
    .WIDTH(32)
) left_15_12 (
    .clk(left_15_12_clk),
    .done(left_15_12_done),
    .in(left_15_12_in),
    .out(left_15_12_out),
    .reset(left_15_12_reset),
    .write_en(left_15_12_write_en)
);
mac_pe pe_15_13 (
    .clk(pe_15_13_clk),
    .done(pe_15_13_done),
    .go(pe_15_13_go),
    .left(pe_15_13_left),
    .mul_ready(pe_15_13_mul_ready),
    .out(pe_15_13_out),
    .reset(pe_15_13_reset),
    .top(pe_15_13_top)
);
std_reg # (
    .WIDTH(32)
) top_15_13 (
    .clk(top_15_13_clk),
    .done(top_15_13_done),
    .in(top_15_13_in),
    .out(top_15_13_out),
    .reset(top_15_13_reset),
    .write_en(top_15_13_write_en)
);
std_reg # (
    .WIDTH(32)
) left_15_13 (
    .clk(left_15_13_clk),
    .done(left_15_13_done),
    .in(left_15_13_in),
    .out(left_15_13_out),
    .reset(left_15_13_reset),
    .write_en(left_15_13_write_en)
);
mac_pe pe_15_14 (
    .clk(pe_15_14_clk),
    .done(pe_15_14_done),
    .go(pe_15_14_go),
    .left(pe_15_14_left),
    .mul_ready(pe_15_14_mul_ready),
    .out(pe_15_14_out),
    .reset(pe_15_14_reset),
    .top(pe_15_14_top)
);
std_reg # (
    .WIDTH(32)
) top_15_14 (
    .clk(top_15_14_clk),
    .done(top_15_14_done),
    .in(top_15_14_in),
    .out(top_15_14_out),
    .reset(top_15_14_reset),
    .write_en(top_15_14_write_en)
);
std_reg # (
    .WIDTH(32)
) left_15_14 (
    .clk(left_15_14_clk),
    .done(left_15_14_done),
    .in(left_15_14_in),
    .out(left_15_14_out),
    .reset(left_15_14_reset),
    .write_en(left_15_14_write_en)
);
mac_pe pe_15_15 (
    .clk(pe_15_15_clk),
    .done(pe_15_15_done),
    .go(pe_15_15_go),
    .left(pe_15_15_left),
    .mul_ready(pe_15_15_mul_ready),
    .out(pe_15_15_out),
    .reset(pe_15_15_reset),
    .top(pe_15_15_top)
);
std_reg # (
    .WIDTH(32)
) top_15_15 (
    .clk(top_15_15_clk),
    .done(top_15_15_done),
    .in(top_15_15_in),
    .out(top_15_15_out),
    .reset(top_15_15_reset),
    .write_en(top_15_15_write_en)
);
std_reg # (
    .WIDTH(32)
) left_15_15 (
    .clk(left_15_15_clk),
    .done(left_15_15_done),
    .in(left_15_15_in),
    .out(left_15_15_out),
    .reset(left_15_15_reset),
    .write_en(left_15_15_write_en)
);
std_reg # (
    .WIDTH(5)
) t0_idx (
    .clk(t0_idx_clk),
    .done(t0_idx_done),
    .in(t0_idx_in),
    .out(t0_idx_out),
    .reset(t0_idx_reset),
    .write_en(t0_idx_write_en)
);
std_add # (
    .WIDTH(5)
) t0_add (
    .left(t0_add_left),
    .out(t0_add_out),
    .right(t0_add_right)
);
std_reg # (
    .WIDTH(5)
) t1_idx (
    .clk(t1_idx_clk),
    .done(t1_idx_done),
    .in(t1_idx_in),
    .out(t1_idx_out),
    .reset(t1_idx_reset),
    .write_en(t1_idx_write_en)
);
std_add # (
    .WIDTH(5)
) t1_add (
    .left(t1_add_left),
    .out(t1_add_out),
    .right(t1_add_right)
);
std_reg # (
    .WIDTH(5)
) t2_idx (
    .clk(t2_idx_clk),
    .done(t2_idx_done),
    .in(t2_idx_in),
    .out(t2_idx_out),
    .reset(t2_idx_reset),
    .write_en(t2_idx_write_en)
);
std_add # (
    .WIDTH(5)
) t2_add (
    .left(t2_add_left),
    .out(t2_add_out),
    .right(t2_add_right)
);
std_reg # (
    .WIDTH(5)
) t3_idx (
    .clk(t3_idx_clk),
    .done(t3_idx_done),
    .in(t3_idx_in),
    .out(t3_idx_out),
    .reset(t3_idx_reset),
    .write_en(t3_idx_write_en)
);
std_add # (
    .WIDTH(5)
) t3_add (
    .left(t3_add_left),
    .out(t3_add_out),
    .right(t3_add_right)
);
std_reg # (
    .WIDTH(5)
) t4_idx (
    .clk(t4_idx_clk),
    .done(t4_idx_done),
    .in(t4_idx_in),
    .out(t4_idx_out),
    .reset(t4_idx_reset),
    .write_en(t4_idx_write_en)
);
std_add # (
    .WIDTH(5)
) t4_add (
    .left(t4_add_left),
    .out(t4_add_out),
    .right(t4_add_right)
);
std_reg # (
    .WIDTH(5)
) t5_idx (
    .clk(t5_idx_clk),
    .done(t5_idx_done),
    .in(t5_idx_in),
    .out(t5_idx_out),
    .reset(t5_idx_reset),
    .write_en(t5_idx_write_en)
);
std_add # (
    .WIDTH(5)
) t5_add (
    .left(t5_add_left),
    .out(t5_add_out),
    .right(t5_add_right)
);
std_reg # (
    .WIDTH(5)
) t6_idx (
    .clk(t6_idx_clk),
    .done(t6_idx_done),
    .in(t6_idx_in),
    .out(t6_idx_out),
    .reset(t6_idx_reset),
    .write_en(t6_idx_write_en)
);
std_add # (
    .WIDTH(5)
) t6_add (
    .left(t6_add_left),
    .out(t6_add_out),
    .right(t6_add_right)
);
std_reg # (
    .WIDTH(5)
) t7_idx (
    .clk(t7_idx_clk),
    .done(t7_idx_done),
    .in(t7_idx_in),
    .out(t7_idx_out),
    .reset(t7_idx_reset),
    .write_en(t7_idx_write_en)
);
std_add # (
    .WIDTH(5)
) t7_add (
    .left(t7_add_left),
    .out(t7_add_out),
    .right(t7_add_right)
);
std_reg # (
    .WIDTH(5)
) t8_idx (
    .clk(t8_idx_clk),
    .done(t8_idx_done),
    .in(t8_idx_in),
    .out(t8_idx_out),
    .reset(t8_idx_reset),
    .write_en(t8_idx_write_en)
);
std_add # (
    .WIDTH(5)
) t8_add (
    .left(t8_add_left),
    .out(t8_add_out),
    .right(t8_add_right)
);
std_reg # (
    .WIDTH(5)
) t9_idx (
    .clk(t9_idx_clk),
    .done(t9_idx_done),
    .in(t9_idx_in),
    .out(t9_idx_out),
    .reset(t9_idx_reset),
    .write_en(t9_idx_write_en)
);
std_add # (
    .WIDTH(5)
) t9_add (
    .left(t9_add_left),
    .out(t9_add_out),
    .right(t9_add_right)
);
std_reg # (
    .WIDTH(5)
) t10_idx (
    .clk(t10_idx_clk),
    .done(t10_idx_done),
    .in(t10_idx_in),
    .out(t10_idx_out),
    .reset(t10_idx_reset),
    .write_en(t10_idx_write_en)
);
std_add # (
    .WIDTH(5)
) t10_add (
    .left(t10_add_left),
    .out(t10_add_out),
    .right(t10_add_right)
);
std_reg # (
    .WIDTH(5)
) t11_idx (
    .clk(t11_idx_clk),
    .done(t11_idx_done),
    .in(t11_idx_in),
    .out(t11_idx_out),
    .reset(t11_idx_reset),
    .write_en(t11_idx_write_en)
);
std_add # (
    .WIDTH(5)
) t11_add (
    .left(t11_add_left),
    .out(t11_add_out),
    .right(t11_add_right)
);
std_reg # (
    .WIDTH(5)
) t12_idx (
    .clk(t12_idx_clk),
    .done(t12_idx_done),
    .in(t12_idx_in),
    .out(t12_idx_out),
    .reset(t12_idx_reset),
    .write_en(t12_idx_write_en)
);
std_add # (
    .WIDTH(5)
) t12_add (
    .left(t12_add_left),
    .out(t12_add_out),
    .right(t12_add_right)
);
std_reg # (
    .WIDTH(5)
) t13_idx (
    .clk(t13_idx_clk),
    .done(t13_idx_done),
    .in(t13_idx_in),
    .out(t13_idx_out),
    .reset(t13_idx_reset),
    .write_en(t13_idx_write_en)
);
std_add # (
    .WIDTH(5)
) t13_add (
    .left(t13_add_left),
    .out(t13_add_out),
    .right(t13_add_right)
);
std_reg # (
    .WIDTH(5)
) t14_idx (
    .clk(t14_idx_clk),
    .done(t14_idx_done),
    .in(t14_idx_in),
    .out(t14_idx_out),
    .reset(t14_idx_reset),
    .write_en(t14_idx_write_en)
);
std_add # (
    .WIDTH(5)
) t14_add (
    .left(t14_add_left),
    .out(t14_add_out),
    .right(t14_add_right)
);
std_reg # (
    .WIDTH(5)
) t15_idx (
    .clk(t15_idx_clk),
    .done(t15_idx_done),
    .in(t15_idx_in),
    .out(t15_idx_out),
    .reset(t15_idx_reset),
    .write_en(t15_idx_write_en)
);
std_add # (
    .WIDTH(5)
) t15_add (
    .left(t15_add_left),
    .out(t15_add_out),
    .right(t15_add_right)
);
std_reg # (
    .WIDTH(5)
) l0_idx (
    .clk(l0_idx_clk),
    .done(l0_idx_done),
    .in(l0_idx_in),
    .out(l0_idx_out),
    .reset(l0_idx_reset),
    .write_en(l0_idx_write_en)
);
std_add # (
    .WIDTH(5)
) l0_add (
    .left(l0_add_left),
    .out(l0_add_out),
    .right(l0_add_right)
);
std_reg # (
    .WIDTH(5)
) l1_idx (
    .clk(l1_idx_clk),
    .done(l1_idx_done),
    .in(l1_idx_in),
    .out(l1_idx_out),
    .reset(l1_idx_reset),
    .write_en(l1_idx_write_en)
);
std_add # (
    .WIDTH(5)
) l1_add (
    .left(l1_add_left),
    .out(l1_add_out),
    .right(l1_add_right)
);
std_reg # (
    .WIDTH(5)
) l2_idx (
    .clk(l2_idx_clk),
    .done(l2_idx_done),
    .in(l2_idx_in),
    .out(l2_idx_out),
    .reset(l2_idx_reset),
    .write_en(l2_idx_write_en)
);
std_add # (
    .WIDTH(5)
) l2_add (
    .left(l2_add_left),
    .out(l2_add_out),
    .right(l2_add_right)
);
std_reg # (
    .WIDTH(5)
) l3_idx (
    .clk(l3_idx_clk),
    .done(l3_idx_done),
    .in(l3_idx_in),
    .out(l3_idx_out),
    .reset(l3_idx_reset),
    .write_en(l3_idx_write_en)
);
std_add # (
    .WIDTH(5)
) l3_add (
    .left(l3_add_left),
    .out(l3_add_out),
    .right(l3_add_right)
);
std_reg # (
    .WIDTH(5)
) l4_idx (
    .clk(l4_idx_clk),
    .done(l4_idx_done),
    .in(l4_idx_in),
    .out(l4_idx_out),
    .reset(l4_idx_reset),
    .write_en(l4_idx_write_en)
);
std_add # (
    .WIDTH(5)
) l4_add (
    .left(l4_add_left),
    .out(l4_add_out),
    .right(l4_add_right)
);
std_reg # (
    .WIDTH(5)
) l5_idx (
    .clk(l5_idx_clk),
    .done(l5_idx_done),
    .in(l5_idx_in),
    .out(l5_idx_out),
    .reset(l5_idx_reset),
    .write_en(l5_idx_write_en)
);
std_add # (
    .WIDTH(5)
) l5_add (
    .left(l5_add_left),
    .out(l5_add_out),
    .right(l5_add_right)
);
std_reg # (
    .WIDTH(5)
) l6_idx (
    .clk(l6_idx_clk),
    .done(l6_idx_done),
    .in(l6_idx_in),
    .out(l6_idx_out),
    .reset(l6_idx_reset),
    .write_en(l6_idx_write_en)
);
std_add # (
    .WIDTH(5)
) l6_add (
    .left(l6_add_left),
    .out(l6_add_out),
    .right(l6_add_right)
);
std_reg # (
    .WIDTH(5)
) l7_idx (
    .clk(l7_idx_clk),
    .done(l7_idx_done),
    .in(l7_idx_in),
    .out(l7_idx_out),
    .reset(l7_idx_reset),
    .write_en(l7_idx_write_en)
);
std_add # (
    .WIDTH(5)
) l7_add (
    .left(l7_add_left),
    .out(l7_add_out),
    .right(l7_add_right)
);
std_reg # (
    .WIDTH(5)
) l8_idx (
    .clk(l8_idx_clk),
    .done(l8_idx_done),
    .in(l8_idx_in),
    .out(l8_idx_out),
    .reset(l8_idx_reset),
    .write_en(l8_idx_write_en)
);
std_add # (
    .WIDTH(5)
) l8_add (
    .left(l8_add_left),
    .out(l8_add_out),
    .right(l8_add_right)
);
std_reg # (
    .WIDTH(5)
) l9_idx (
    .clk(l9_idx_clk),
    .done(l9_idx_done),
    .in(l9_idx_in),
    .out(l9_idx_out),
    .reset(l9_idx_reset),
    .write_en(l9_idx_write_en)
);
std_add # (
    .WIDTH(5)
) l9_add (
    .left(l9_add_left),
    .out(l9_add_out),
    .right(l9_add_right)
);
std_reg # (
    .WIDTH(5)
) l10_idx (
    .clk(l10_idx_clk),
    .done(l10_idx_done),
    .in(l10_idx_in),
    .out(l10_idx_out),
    .reset(l10_idx_reset),
    .write_en(l10_idx_write_en)
);
std_add # (
    .WIDTH(5)
) l10_add (
    .left(l10_add_left),
    .out(l10_add_out),
    .right(l10_add_right)
);
std_reg # (
    .WIDTH(5)
) l11_idx (
    .clk(l11_idx_clk),
    .done(l11_idx_done),
    .in(l11_idx_in),
    .out(l11_idx_out),
    .reset(l11_idx_reset),
    .write_en(l11_idx_write_en)
);
std_add # (
    .WIDTH(5)
) l11_add (
    .left(l11_add_left),
    .out(l11_add_out),
    .right(l11_add_right)
);
std_reg # (
    .WIDTH(5)
) l12_idx (
    .clk(l12_idx_clk),
    .done(l12_idx_done),
    .in(l12_idx_in),
    .out(l12_idx_out),
    .reset(l12_idx_reset),
    .write_en(l12_idx_write_en)
);
std_add # (
    .WIDTH(5)
) l12_add (
    .left(l12_add_left),
    .out(l12_add_out),
    .right(l12_add_right)
);
std_reg # (
    .WIDTH(5)
) l13_idx (
    .clk(l13_idx_clk),
    .done(l13_idx_done),
    .in(l13_idx_in),
    .out(l13_idx_out),
    .reset(l13_idx_reset),
    .write_en(l13_idx_write_en)
);
std_add # (
    .WIDTH(5)
) l13_add (
    .left(l13_add_left),
    .out(l13_add_out),
    .right(l13_add_right)
);
std_reg # (
    .WIDTH(5)
) l14_idx (
    .clk(l14_idx_clk),
    .done(l14_idx_done),
    .in(l14_idx_in),
    .out(l14_idx_out),
    .reset(l14_idx_reset),
    .write_en(l14_idx_write_en)
);
std_add # (
    .WIDTH(5)
) l14_add (
    .left(l14_add_left),
    .out(l14_add_out),
    .right(l14_add_right)
);
std_reg # (
    .WIDTH(5)
) l15_idx (
    .clk(l15_idx_clk),
    .done(l15_idx_done),
    .in(l15_idx_in),
    .out(l15_idx_out),
    .reset(l15_idx_reset),
    .write_en(l15_idx_write_en)
);
std_add # (
    .WIDTH(5)
) l15_add (
    .left(l15_add_left),
    .out(l15_add_out),
    .right(l15_add_right)
);
std_reg # (
    .WIDTH(6)
) idx (
    .clk(idx_clk),
    .done(idx_done),
    .in(idx_in),
    .out(idx_out),
    .reset(idx_reset),
    .write_en(idx_write_en)
);
std_add # (
    .WIDTH(6)
) idx_add (
    .left(idx_add_left),
    .out(idx_add_out),
    .right(idx_add_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_16_20_reg (
    .clk(idx_between_16_20_reg_clk),
    .done(idx_between_16_20_reg_done),
    .in(idx_between_16_20_reg_in),
    .out(idx_between_16_20_reg_out),
    .reset(idx_between_16_20_reg_reset),
    .write_en(idx_between_16_20_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_20 (
    .left(index_lt_20_left),
    .out(index_lt_20_out),
    .right(index_lt_20_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_16 (
    .left(index_ge_16_left),
    .out(index_ge_16_out),
    .right(index_ge_16_right)
);
std_and # (
    .WIDTH(1)
) idx_between_16_20_comb (
    .left(idx_between_16_20_comb_left),
    .out(idx_between_16_20_comb_out),
    .right(idx_between_16_20_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_26_30_reg (
    .clk(idx_between_26_30_reg_clk),
    .done(idx_between_26_30_reg_done),
    .in(idx_between_26_30_reg_in),
    .out(idx_between_26_30_reg_out),
    .reset(idx_between_26_30_reg_reset),
    .write_en(idx_between_26_30_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_30 (
    .left(index_lt_30_left),
    .out(index_lt_30_out),
    .right(index_lt_30_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_26 (
    .left(index_ge_26_left),
    .out(index_ge_26_out),
    .right(index_ge_26_right)
);
std_and # (
    .WIDTH(1)
) idx_between_26_30_comb (
    .left(idx_between_26_30_comb_left),
    .out(idx_between_26_30_comb_out),
    .right(idx_between_26_30_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_30_46_reg (
    .clk(idx_between_30_46_reg_clk),
    .done(idx_between_30_46_reg_done),
    .in(idx_between_30_46_reg_in),
    .out(idx_between_30_46_reg_out),
    .reset(idx_between_30_46_reg_reset),
    .write_en(idx_between_30_46_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_46 (
    .left(index_lt_46_left),
    .out(index_lt_46_out),
    .right(index_lt_46_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_30 (
    .left(index_ge_30_left),
    .out(index_ge_30_out),
    .right(index_ge_30_right)
);
std_and # (
    .WIDTH(1)
) idx_between_30_46_comb (
    .left(idx_between_30_46_comb_left),
    .out(idx_between_30_46_comb_out),
    .right(idx_between_30_46_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_44_45_reg (
    .clk(idx_between_44_45_reg_clk),
    .done(idx_between_44_45_reg_done),
    .in(idx_between_44_45_reg_in),
    .out(idx_between_44_45_reg_out),
    .reset(idx_between_44_45_reg_reset),
    .write_en(idx_between_44_45_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_45 (
    .left(index_lt_45_left),
    .out(index_lt_45_out),
    .right(index_lt_45_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_44 (
    .left(index_ge_44_left),
    .out(index_ge_44_out),
    .right(index_ge_44_right)
);
std_and # (
    .WIDTH(1)
) idx_between_44_45_comb (
    .left(idx_between_44_45_comb_left),
    .out(idx_between_44_45_comb_out),
    .right(idx_between_44_45_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_25_41_reg (
    .clk(idx_between_25_41_reg_clk),
    .done(idx_between_25_41_reg_done),
    .in(idx_between_25_41_reg_in),
    .out(idx_between_25_41_reg_out),
    .reset(idx_between_25_41_reg_reset),
    .write_en(idx_between_25_41_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_41 (
    .left(index_lt_41_left),
    .out(index_lt_41_out),
    .right(index_lt_41_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_25 (
    .left(index_ge_25_left),
    .out(index_ge_25_out),
    .right(index_ge_25_right)
);
std_and # (
    .WIDTH(1)
) idx_between_25_41_comb (
    .left(idx_between_25_41_comb_left),
    .out(idx_between_25_41_comb_out),
    .right(idx_between_25_41_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_35_51_reg (
    .clk(idx_between_35_51_reg_clk),
    .done(idx_between_35_51_reg_done),
    .in(idx_between_35_51_reg_in),
    .out(idx_between_35_51_reg_out),
    .reset(idx_between_35_51_reg_reset),
    .write_en(idx_between_35_51_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_51 (
    .left(index_lt_51_left),
    .out(index_lt_51_out),
    .right(index_lt_51_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_35 (
    .left(index_ge_35_left),
    .out(index_ge_35_out),
    .right(index_ge_35_right)
);
std_and # (
    .WIDTH(1)
) idx_between_35_51_comb (
    .left(idx_between_35_51_comb_left),
    .out(idx_between_35_51_comb_out),
    .right(idx_between_35_51_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_22_26_reg (
    .clk(idx_between_22_26_reg_clk),
    .done(idx_between_22_26_reg_done),
    .in(idx_between_22_26_reg_in),
    .out(idx_between_22_26_reg_out),
    .reset(idx_between_22_26_reg_reset),
    .write_en(idx_between_22_26_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_26 (
    .left(index_lt_26_left),
    .out(index_lt_26_out),
    .right(index_lt_26_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_22 (
    .left(index_ge_22_left),
    .out(index_ge_22_out),
    .right(index_ge_22_right)
);
std_and # (
    .WIDTH(1)
) idx_between_22_26_comb (
    .left(idx_between_22_26_comb_left),
    .out(idx_between_22_26_comb_out),
    .right(idx_between_22_26_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_40_41_reg (
    .clk(idx_between_40_41_reg_clk),
    .done(idx_between_40_41_reg_done),
    .in(idx_between_40_41_reg_in),
    .out(idx_between_40_41_reg_out),
    .reset(idx_between_40_41_reg_reset),
    .write_en(idx_between_40_41_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_40 (
    .left(index_ge_40_left),
    .out(index_ge_40_out),
    .right(index_ge_40_right)
);
std_and # (
    .WIDTH(1)
) idx_between_40_41_comb (
    .left(idx_between_40_41_comb_left),
    .out(idx_between_40_41_comb_out),
    .right(idx_between_40_41_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_17_21_reg (
    .clk(idx_between_17_21_reg_clk),
    .done(idx_between_17_21_reg_done),
    .in(idx_between_17_21_reg_in),
    .out(idx_between_17_21_reg_out),
    .reset(idx_between_17_21_reg_reset),
    .write_en(idx_between_17_21_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_21 (
    .left(index_lt_21_left),
    .out(index_lt_21_out),
    .right(index_lt_21_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_17 (
    .left(index_ge_17_left),
    .out(index_ge_17_out),
    .right(index_ge_17_right)
);
std_and # (
    .WIDTH(1)
) idx_between_17_21_comb (
    .left(idx_between_17_21_comb_left),
    .out(idx_between_17_21_comb_out),
    .right(idx_between_17_21_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_21_37_reg (
    .clk(idx_between_21_37_reg_clk),
    .done(idx_between_21_37_reg_done),
    .in(idx_between_21_37_reg_in),
    .out(idx_between_21_37_reg_out),
    .reset(idx_between_21_37_reg_reset),
    .write_en(idx_between_21_37_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_37 (
    .left(index_lt_37_left),
    .out(index_lt_37_out),
    .right(index_lt_37_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_21 (
    .left(index_ge_21_left),
    .out(index_ge_21_out),
    .right(index_ge_21_right)
);
std_and # (
    .WIDTH(1)
) idx_between_21_37_comb (
    .left(idx_between_21_37_comb_left),
    .out(idx_between_21_37_comb_out),
    .right(idx_between_21_37_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_31_47_reg (
    .clk(idx_between_31_47_reg_clk),
    .done(idx_between_31_47_reg_done),
    .in(idx_between_31_47_reg_in),
    .out(idx_between_31_47_reg_out),
    .reset(idx_between_31_47_reg_reset),
    .write_en(idx_between_31_47_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_47 (
    .left(index_lt_47_left),
    .out(index_lt_47_out),
    .right(index_lt_47_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_31 (
    .left(index_ge_31_left),
    .out(index_ge_31_out),
    .right(index_ge_31_right)
);
std_and # (
    .WIDTH(1)
) idx_between_31_47_comb (
    .left(idx_between_31_47_comb_left),
    .out(idx_between_31_47_comb_out),
    .right(idx_between_31_47_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_13_17_reg (
    .clk(idx_between_13_17_reg_clk),
    .done(idx_between_13_17_reg_done),
    .in(idx_between_13_17_reg_in),
    .out(idx_between_13_17_reg_out),
    .reset(idx_between_13_17_reg_reset),
    .write_en(idx_between_13_17_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_17 (
    .left(index_lt_17_left),
    .out(index_lt_17_out),
    .right(index_lt_17_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_13 (
    .left(index_ge_13_left),
    .out(index_ge_13_out),
    .right(index_ge_13_right)
);
std_and # (
    .WIDTH(1)
) idx_between_13_17_comb (
    .left(idx_between_13_17_comb_left),
    .out(idx_between_13_17_comb_out),
    .right(idx_between_13_17_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_27_43_reg (
    .clk(idx_between_27_43_reg_clk),
    .done(idx_between_27_43_reg_done),
    .in(idx_between_27_43_reg_in),
    .out(idx_between_27_43_reg_out),
    .reset(idx_between_27_43_reg_reset),
    .write_en(idx_between_27_43_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_43 (
    .left(index_lt_43_left),
    .out(index_lt_43_out),
    .right(index_lt_43_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_27 (
    .left(index_ge_27_left),
    .out(index_ge_27_out),
    .right(index_ge_27_right)
);
std_and # (
    .WIDTH(1)
) idx_between_27_43_comb (
    .left(idx_between_27_43_comb_left),
    .out(idx_between_27_43_comb_out),
    .right(idx_between_27_43_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_41_42_reg (
    .clk(idx_between_41_42_reg_clk),
    .done(idx_between_41_42_reg_done),
    .in(idx_between_41_42_reg_in),
    .out(idx_between_41_42_reg_out),
    .reset(idx_between_41_42_reg_reset),
    .write_en(idx_between_41_42_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_42 (
    .left(index_lt_42_left),
    .out(index_lt_42_out),
    .right(index_lt_42_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_41 (
    .left(index_ge_41_left),
    .out(index_ge_41_out),
    .right(index_ge_41_right)
);
std_and # (
    .WIDTH(1)
) idx_between_41_42_comb (
    .left(idx_between_41_42_comb_left),
    .out(idx_between_41_42_comb_out),
    .right(idx_between_41_42_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_23_27_reg (
    .clk(idx_between_23_27_reg_clk),
    .done(idx_between_23_27_reg_done),
    .in(idx_between_23_27_reg_in),
    .out(idx_between_23_27_reg_out),
    .reset(idx_between_23_27_reg_reset),
    .write_en(idx_between_23_27_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_27 (
    .left(index_lt_27_left),
    .out(index_lt_27_out),
    .right(index_lt_27_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_23 (
    .left(index_ge_23_left),
    .out(index_ge_23_out),
    .right(index_ge_23_right)
);
std_and # (
    .WIDTH(1)
) idx_between_23_27_comb (
    .left(idx_between_23_27_comb_left),
    .out(idx_between_23_27_comb_out),
    .right(idx_between_23_27_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_5_21_reg (
    .clk(idx_between_5_21_reg_clk),
    .done(idx_between_5_21_reg_done),
    .in(idx_between_5_21_reg_in),
    .out(idx_between_5_21_reg_out),
    .reset(idx_between_5_21_reg_reset),
    .write_en(idx_between_5_21_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_5 (
    .left(index_ge_5_left),
    .out(index_ge_5_out),
    .right(index_ge_5_right)
);
std_and # (
    .WIDTH(1)
) idx_between_5_21_comb (
    .left(idx_between_5_21_comb_left),
    .out(idx_between_5_21_comb_out),
    .right(idx_between_5_21_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_0_16_reg (
    .clk(idx_between_0_16_reg_clk),
    .done(idx_between_0_16_reg_done),
    .in(idx_between_0_16_reg_in),
    .out(idx_between_0_16_reg_out),
    .reset(idx_between_0_16_reg_reset),
    .write_en(idx_between_0_16_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_16 (
    .left(index_lt_16_left),
    .out(index_lt_16_out),
    .right(index_lt_16_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_1_17_reg (
    .clk(idx_between_1_17_reg_clk),
    .done(idx_between_1_17_reg_done),
    .in(idx_between_1_17_reg_in),
    .out(idx_between_1_17_reg_out),
    .reset(idx_between_1_17_reg_reset),
    .write_en(idx_between_1_17_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_1 (
    .left(index_ge_1_left),
    .out(index_ge_1_out),
    .right(index_ge_1_right)
);
std_and # (
    .WIDTH(1)
) idx_between_1_17_comb (
    .left(idx_between_1_17_comb_left),
    .out(idx_between_1_17_comb_out),
    .right(idx_between_1_17_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_47_48_reg (
    .clk(idx_between_47_48_reg_clk),
    .done(idx_between_47_48_reg_done),
    .in(idx_between_47_48_reg_in),
    .out(idx_between_47_48_reg_out),
    .reset(idx_between_47_48_reg_reset),
    .write_en(idx_between_47_48_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_48 (
    .left(index_lt_48_left),
    .out(index_lt_48_out),
    .right(index_lt_48_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_47 (
    .left(index_ge_47_left),
    .out(index_ge_47_out),
    .right(index_ge_47_right)
);
std_and # (
    .WIDTH(1)
) idx_between_47_48_comb (
    .left(idx_between_47_48_comb_left),
    .out(idx_between_47_48_comb_out),
    .right(idx_between_47_48_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_24_28_reg (
    .clk(idx_between_24_28_reg_clk),
    .done(idx_between_24_28_reg_done),
    .in(idx_between_24_28_reg_in),
    .out(idx_between_24_28_reg_out),
    .reset(idx_between_24_28_reg_reset),
    .write_en(idx_between_24_28_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_28 (
    .left(index_lt_28_left),
    .out(index_lt_28_out),
    .right(index_lt_28_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_24 (
    .left(index_ge_24_left),
    .out(index_ge_24_out),
    .right(index_ge_24_right)
);
std_and # (
    .WIDTH(1)
) idx_between_24_28_comb (
    .left(idx_between_24_28_comb_left),
    .out(idx_between_24_28_comb_out),
    .right(idx_between_24_28_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_42_43_reg (
    .clk(idx_between_42_43_reg_clk),
    .done(idx_between_42_43_reg_done),
    .in(idx_between_42_43_reg_in),
    .out(idx_between_42_43_reg_out),
    .reset(idx_between_42_43_reg_reset),
    .write_en(idx_between_42_43_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_42 (
    .left(index_ge_42_left),
    .out(index_ge_42_out),
    .right(index_ge_42_right)
);
std_and # (
    .WIDTH(1)
) idx_between_42_43_comb (
    .left(idx_between_42_43_comb_left),
    .out(idx_between_42_43_comb_out),
    .right(idx_between_42_43_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_33_49_reg (
    .clk(idx_between_33_49_reg_clk),
    .done(idx_between_33_49_reg_done),
    .in(idx_between_33_49_reg_in),
    .out(idx_between_33_49_reg_out),
    .reset(idx_between_33_49_reg_reset),
    .write_en(idx_between_33_49_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_49 (
    .left(index_lt_49_left),
    .out(index_lt_49_out),
    .right(index_lt_49_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_33 (
    .left(index_ge_33_left),
    .out(index_ge_33_out),
    .right(index_ge_33_right)
);
std_and # (
    .WIDTH(1)
) idx_between_33_49_comb (
    .left(idx_between_33_49_comb_left),
    .out(idx_between_33_49_comb_out),
    .right(idx_between_33_49_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_20_24_reg (
    .clk(idx_between_20_24_reg_clk),
    .done(idx_between_20_24_reg_done),
    .in(idx_between_20_24_reg_in),
    .out(idx_between_20_24_reg_out),
    .reset(idx_between_20_24_reg_reset),
    .write_en(idx_between_20_24_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_24 (
    .left(index_lt_24_left),
    .out(index_lt_24_out),
    .right(index_lt_24_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_20 (
    .left(index_ge_20_left),
    .out(index_ge_20_out),
    .right(index_ge_20_right)
);
std_and # (
    .WIDTH(1)
) idx_between_20_24_comb (
    .left(idx_between_20_24_comb_left),
    .out(idx_between_20_24_comb_out),
    .right(idx_between_20_24_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_38_39_reg (
    .clk(idx_between_38_39_reg_clk),
    .done(idx_between_38_39_reg_done),
    .in(idx_between_38_39_reg_in),
    .out(idx_between_38_39_reg_out),
    .reset(idx_between_38_39_reg_reset),
    .write_en(idx_between_38_39_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_39 (
    .left(index_lt_39_left),
    .out(index_lt_39_out),
    .right(index_lt_39_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_38 (
    .left(index_ge_38_left),
    .out(index_ge_38_out),
    .right(index_ge_38_right)
);
std_and # (
    .WIDTH(1)
) idx_between_38_39_comb (
    .left(idx_between_38_39_comb_left),
    .out(idx_between_38_39_comb_out),
    .right(idx_between_38_39_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_48_49_reg (
    .clk(idx_between_48_49_reg_clk),
    .done(idx_between_48_49_reg_done),
    .in(idx_between_48_49_reg_in),
    .out(idx_between_48_49_reg_out),
    .reset(idx_between_48_49_reg_reset),
    .write_en(idx_between_48_49_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_48 (
    .left(index_ge_48_left),
    .out(index_ge_48_out),
    .right(index_ge_48_right)
);
std_and # (
    .WIDTH(1)
) idx_between_48_49_comb (
    .left(idx_between_48_49_comb_left),
    .out(idx_between_48_49_comb_out),
    .right(idx_between_48_49_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_29_45_reg (
    .clk(idx_between_29_45_reg_clk),
    .done(idx_between_29_45_reg_done),
    .in(idx_between_29_45_reg_in),
    .out(idx_between_29_45_reg_out),
    .reset(idx_between_29_45_reg_reset),
    .write_en(idx_between_29_45_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_29 (
    .left(index_ge_29_left),
    .out(index_ge_29_out),
    .right(index_ge_29_right)
);
std_and # (
    .WIDTH(1)
) idx_between_29_45_comb (
    .left(idx_between_29_45_comb_left),
    .out(idx_between_29_45_comb_out),
    .right(idx_between_29_45_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_30_34_reg (
    .clk(idx_between_30_34_reg_clk),
    .done(idx_between_30_34_reg_done),
    .in(idx_between_30_34_reg_in),
    .out(idx_between_30_34_reg_out),
    .reset(idx_between_30_34_reg_reset),
    .write_en(idx_between_30_34_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_34 (
    .left(index_lt_34_left),
    .out(index_lt_34_out),
    .right(index_lt_34_right)
);
std_and # (
    .WIDTH(1)
) idx_between_30_34_comb (
    .left(idx_between_30_34_comb_left),
    .out(idx_between_30_34_comb_out),
    .right(idx_between_30_34_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_25_29_reg (
    .clk(idx_between_25_29_reg_clk),
    .done(idx_between_25_29_reg_done),
    .in(idx_between_25_29_reg_in),
    .out(idx_between_25_29_reg_out),
    .reset(idx_between_25_29_reg_reset),
    .write_en(idx_between_25_29_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_29 (
    .left(index_lt_29_left),
    .out(index_lt_29_out),
    .right(index_lt_29_right)
);
std_and # (
    .WIDTH(1)
) idx_between_25_29_comb (
    .left(idx_between_25_29_comb_left),
    .out(idx_between_25_29_comb_out),
    .right(idx_between_25_29_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_7_23_reg (
    .clk(idx_between_7_23_reg_clk),
    .done(idx_between_7_23_reg_done),
    .in(idx_between_7_23_reg_in),
    .out(idx_between_7_23_reg_out),
    .reset(idx_between_7_23_reg_reset),
    .write_en(idx_between_7_23_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_23 (
    .left(index_lt_23_left),
    .out(index_lt_23_out),
    .right(index_lt_23_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_7 (
    .left(index_ge_7_left),
    .out(index_ge_7_out),
    .right(index_ge_7_right)
);
std_and # (
    .WIDTH(1)
) idx_between_7_23_comb (
    .left(idx_between_7_23_comb_left),
    .out(idx_between_7_23_comb_out),
    .right(idx_between_7_23_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_22_23_reg (
    .clk(idx_between_22_23_reg_clk),
    .done(idx_between_22_23_reg_done),
    .in(idx_between_22_23_reg_in),
    .out(idx_between_22_23_reg_out),
    .reset(idx_between_22_23_reg_reset),
    .write_en(idx_between_22_23_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_22_23_comb (
    .left(idx_between_22_23_comb_left),
    .out(idx_between_22_23_comb_out),
    .right(idx_between_22_23_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_21_25_reg (
    .clk(idx_between_21_25_reg_clk),
    .done(idx_between_21_25_reg_done),
    .in(idx_between_21_25_reg_in),
    .out(idx_between_21_25_reg_out),
    .reset(idx_between_21_25_reg_reset),
    .write_en(idx_between_21_25_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_25 (
    .left(index_lt_25_left),
    .out(index_lt_25_out),
    .right(index_lt_25_right)
);
std_and # (
    .WIDTH(1)
) idx_between_21_25_comb (
    .left(idx_between_21_25_comb_left),
    .out(idx_between_21_25_comb_out),
    .right(idx_between_21_25_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_3_19_reg (
    .clk(idx_between_3_19_reg_clk),
    .done(idx_between_3_19_reg_done),
    .in(idx_between_3_19_reg_in),
    .out(idx_between_3_19_reg_out),
    .reset(idx_between_3_19_reg_reset),
    .write_en(idx_between_3_19_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_19 (
    .left(index_lt_19_left),
    .out(index_lt_19_out),
    .right(index_lt_19_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_3 (
    .left(index_ge_3_left),
    .out(index_ge_3_out),
    .right(index_ge_3_right)
);
std_and # (
    .WIDTH(1)
) idx_between_3_19_comb (
    .left(idx_between_3_19_comb_left),
    .out(idx_between_3_19_comb_out),
    .right(idx_between_3_19_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_31_35_reg (
    .clk(idx_between_31_35_reg_clk),
    .done(idx_between_31_35_reg_done),
    .in(idx_between_31_35_reg_in),
    .out(idx_between_31_35_reg_out),
    .reset(idx_between_31_35_reg_reset),
    .write_en(idx_between_31_35_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_35 (
    .left(index_lt_35_left),
    .out(index_lt_35_out),
    .right(index_lt_35_right)
);
std_and # (
    .WIDTH(1)
) idx_between_31_35_comb (
    .left(idx_between_31_35_comb_left),
    .out(idx_between_31_35_comb_out),
    .right(idx_between_31_35_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_49_50_reg (
    .clk(idx_between_49_50_reg_clk),
    .done(idx_between_49_50_reg_done),
    .in(idx_between_49_50_reg_in),
    .out(idx_between_49_50_reg_out),
    .reset(idx_between_49_50_reg_reset),
    .write_en(idx_between_49_50_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_50 (
    .left(index_lt_50_left),
    .out(index_lt_50_out),
    .right(index_lt_50_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_49 (
    .left(index_ge_49_left),
    .out(index_ge_49_out),
    .right(index_ge_49_right)
);
std_and # (
    .WIDTH(1)
) idx_between_49_50_comb (
    .left(idx_between_49_50_comb_left),
    .out(idx_between_49_50_comb_out),
    .right(idx_between_49_50_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_27_31_reg (
    .clk(idx_between_27_31_reg_clk),
    .done(idx_between_27_31_reg_done),
    .in(idx_between_27_31_reg_in),
    .out(idx_between_27_31_reg_out),
    .reset(idx_between_27_31_reg_reset),
    .write_en(idx_between_27_31_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_31 (
    .left(index_lt_31_left),
    .out(index_lt_31_out),
    .right(index_lt_31_right)
);
std_and # (
    .WIDTH(1)
) idx_between_27_31_comb (
    .left(idx_between_27_31_comb_left),
    .out(idx_between_27_31_comb_out),
    .right(idx_between_27_31_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_45_46_reg (
    .clk(idx_between_45_46_reg_clk),
    .done(idx_between_45_46_reg_done),
    .in(idx_between_45_46_reg_in),
    .out(idx_between_45_46_reg_out),
    .reset(idx_between_45_46_reg_reset),
    .write_en(idx_between_45_46_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_45 (
    .left(index_ge_45_left),
    .out(index_ge_45_out),
    .right(index_ge_45_right)
);
std_and # (
    .WIDTH(1)
) idx_between_45_46_comb (
    .left(idx_between_45_46_comb_left),
    .out(idx_between_45_46_comb_out),
    .right(idx_between_45_46_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_50_51_reg (
    .clk(idx_between_50_51_reg_clk),
    .done(idx_between_50_51_reg_done),
    .in(idx_between_50_51_reg_in),
    .out(idx_between_50_51_reg_out),
    .reset(idx_between_50_51_reg_reset),
    .write_en(idx_between_50_51_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_50 (
    .left(index_ge_50_left),
    .out(index_ge_50_out),
    .right(index_ge_50_right)
);
std_and # (
    .WIDTH(1)
) idx_between_50_51_comb (
    .left(idx_between_50_51_comb_left),
    .out(idx_between_50_51_comb_out),
    .right(idx_between_50_51_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_51_52_reg (
    .clk(idx_between_51_52_reg_clk),
    .done(idx_between_51_52_reg_done),
    .in(idx_between_51_52_reg_in),
    .out(idx_between_51_52_reg_out),
    .reset(idx_between_51_52_reg_reset),
    .write_en(idx_between_51_52_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_52 (
    .left(index_lt_52_left),
    .out(index_lt_52_out),
    .right(index_lt_52_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_51 (
    .left(index_ge_51_left),
    .out(index_ge_51_out),
    .right(index_ge_51_right)
);
std_and # (
    .WIDTH(1)
) idx_between_51_52_comb (
    .left(idx_between_51_52_comb_left),
    .out(idx_between_51_52_comb_out),
    .right(idx_between_51_52_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_32_48_reg (
    .clk(idx_between_32_48_reg_clk),
    .done(idx_between_32_48_reg_done),
    .in(idx_between_32_48_reg_in),
    .out(idx_between_32_48_reg_out),
    .reset(idx_between_32_48_reg_reset),
    .write_en(idx_between_32_48_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_32 (
    .left(index_ge_32_left),
    .out(index_ge_32_out),
    .right(index_ge_32_right)
);
std_and # (
    .WIDTH(1)
) idx_between_32_48_comb (
    .left(idx_between_32_48_comb_left),
    .out(idx_between_32_48_comb_out),
    .right(idx_between_32_48_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_5_9_reg (
    .clk(idx_between_5_9_reg_clk),
    .done(idx_between_5_9_reg_done),
    .in(idx_between_5_9_reg_in),
    .out(idx_between_5_9_reg_out),
    .reset(idx_between_5_9_reg_reset),
    .write_en(idx_between_5_9_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_9 (
    .left(index_lt_9_left),
    .out(index_lt_9_out),
    .right(index_lt_9_right)
);
std_and # (
    .WIDTH(1)
) idx_between_5_9_comb (
    .left(idx_between_5_9_comb_left),
    .out(idx_between_5_9_comb_out),
    .right(idx_between_5_9_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_46_47_reg (
    .clk(idx_between_46_47_reg_clk),
    .done(idx_between_46_47_reg_done),
    .in(idx_between_46_47_reg_in),
    .out(idx_between_46_47_reg_out),
    .reset(idx_between_46_47_reg_reset),
    .write_en(idx_between_46_47_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_46 (
    .left(index_ge_46_left),
    .out(index_ge_46_out),
    .right(index_ge_46_right)
);
std_and # (
    .WIDTH(1)
) idx_between_46_47_comb (
    .left(idx_between_46_47_comb_left),
    .out(idx_between_46_47_comb_out),
    .right(idx_between_46_47_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_23_24_reg (
    .clk(idx_between_23_24_reg_clk),
    .done(idx_between_23_24_reg_done),
    .in(idx_between_23_24_reg_in),
    .out(idx_between_23_24_reg_out),
    .reset(idx_between_23_24_reg_reset),
    .write_en(idx_between_23_24_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_23_24_comb (
    .left(idx_between_23_24_comb_left),
    .out(idx_between_23_24_comb_out),
    .right(idx_between_23_24_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_4_20_reg (
    .clk(idx_between_4_20_reg_clk),
    .done(idx_between_4_20_reg_done),
    .in(idx_between_4_20_reg_in),
    .out(idx_between_4_20_reg_out),
    .reset(idx_between_4_20_reg_reset),
    .write_en(idx_between_4_20_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_4 (
    .left(index_ge_4_left),
    .out(index_ge_4_out),
    .right(index_ge_4_right)
);
std_and # (
    .WIDTH(1)
) idx_between_4_20_comb (
    .left(idx_between_4_20_comb_left),
    .out(idx_between_4_20_comb_out),
    .right(idx_between_4_20_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_14_30_reg (
    .clk(idx_between_14_30_reg_clk),
    .done(idx_between_14_30_reg_done),
    .in(idx_between_14_30_reg_in),
    .out(idx_between_14_30_reg_out),
    .reset(idx_between_14_30_reg_reset),
    .write_en(idx_between_14_30_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_14 (
    .left(index_ge_14_left),
    .out(index_ge_14_out),
    .right(index_ge_14_right)
);
std_and # (
    .WIDTH(1)
) idx_between_14_30_comb (
    .left(idx_between_14_30_comb_left),
    .out(idx_between_14_30_comb_out),
    .right(idx_between_14_30_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_1_5_reg (
    .clk(idx_between_1_5_reg_clk),
    .done(idx_between_1_5_reg_done),
    .in(idx_between_1_5_reg_in),
    .out(idx_between_1_5_reg_out),
    .reset(idx_between_1_5_reg_reset),
    .write_en(idx_between_1_5_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_5 (
    .left(index_lt_5_left),
    .out(index_lt_5_out),
    .right(index_lt_5_right)
);
std_and # (
    .WIDTH(1)
) idx_between_1_5_comb (
    .left(idx_between_1_5_comb_left),
    .out(idx_between_1_5_comb_out),
    .right(idx_between_1_5_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_28_32_reg (
    .clk(idx_between_28_32_reg_clk),
    .done(idx_between_28_32_reg_done),
    .in(idx_between_28_32_reg_in),
    .out(idx_between_28_32_reg_out),
    .reset(idx_between_28_32_reg_reset),
    .write_en(idx_between_28_32_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_32 (
    .left(index_lt_32_left),
    .out(index_lt_32_out),
    .right(index_lt_32_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_28 (
    .left(index_ge_28_left),
    .out(index_ge_28_out),
    .right(index_ge_28_right)
);
std_and # (
    .WIDTH(1)
) idx_between_28_32_comb (
    .left(idx_between_28_32_comb_left),
    .out(idx_between_28_32_comb_out),
    .right(idx_between_28_32_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_10_26_reg (
    .clk(idx_between_10_26_reg_clk),
    .done(idx_between_10_26_reg_done),
    .in(idx_between_10_26_reg_in),
    .out(idx_between_10_26_reg_out),
    .reset(idx_between_10_26_reg_reset),
    .write_en(idx_between_10_26_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_10 (
    .left(index_ge_10_left),
    .out(index_ge_10_out),
    .right(index_ge_10_right)
);
std_and # (
    .WIDTH(1)
) idx_between_10_26_comb (
    .left(idx_between_10_26_comb_left),
    .out(idx_between_10_26_comb_out),
    .right(idx_between_10_26_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_24_25_reg (
    .clk(idx_between_24_25_reg_clk),
    .done(idx_between_24_25_reg_done),
    .in(idx_between_24_25_reg_in),
    .out(idx_between_24_25_reg_out),
    .reset(idx_between_24_25_reg_reset),
    .write_en(idx_between_24_25_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_24_25_comb (
    .left(idx_between_24_25_comb_left),
    .out(idx_between_24_25_comb_out),
    .right(idx_between_24_25_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_6_22_reg (
    .clk(idx_between_6_22_reg_clk),
    .done(idx_between_6_22_reg_done),
    .in(idx_between_6_22_reg_in),
    .out(idx_between_6_22_reg_out),
    .reset(idx_between_6_22_reg_reset),
    .write_en(idx_between_6_22_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_22 (
    .left(index_lt_22_left),
    .out(index_lt_22_out),
    .right(index_lt_22_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_6 (
    .left(index_ge_6_left),
    .out(index_ge_6_out),
    .right(index_ge_6_right)
);
std_and # (
    .WIDTH(1)
) idx_between_6_22_comb (
    .left(idx_between_6_22_comb_left),
    .out(idx_between_6_22_comb_out),
    .right(idx_between_6_22_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_29_33_reg (
    .clk(idx_between_29_33_reg_clk),
    .done(idx_between_29_33_reg_done),
    .in(idx_between_29_33_reg_in),
    .out(idx_between_29_33_reg_out),
    .reset(idx_between_29_33_reg_reset),
    .write_en(idx_between_29_33_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_33 (
    .left(index_lt_33_left),
    .out(index_lt_33_out),
    .right(index_lt_33_right)
);
std_and # (
    .WIDTH(1)
) idx_between_29_33_comb (
    .left(idx_between_29_33_comb_left),
    .out(idx_between_29_33_comb_out),
    .right(idx_between_29_33_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_2_6_reg (
    .clk(idx_between_2_6_reg_clk),
    .done(idx_between_2_6_reg_done),
    .in(idx_between_2_6_reg_in),
    .out(idx_between_2_6_reg_out),
    .reset(idx_between_2_6_reg_reset),
    .write_en(idx_between_2_6_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_6 (
    .left(index_lt_6_left),
    .out(index_lt_6_out),
    .right(index_lt_6_right)
);
std_ge # (
    .WIDTH(6)
) index_ge_2 (
    .left(index_ge_2_left),
    .out(index_ge_2_out),
    .right(index_ge_2_right)
);
std_and # (
    .WIDTH(1)
) idx_between_2_6_comb (
    .left(idx_between_2_6_comb_left),
    .out(idx_between_2_6_comb_out),
    .right(idx_between_2_6_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_30_31_reg (
    .clk(idx_between_30_31_reg_clk),
    .done(idx_between_30_31_reg_done),
    .in(idx_between_30_31_reg_in),
    .out(idx_between_30_31_reg_out),
    .reset(idx_between_30_31_reg_reset),
    .write_en(idx_between_30_31_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_30_31_comb (
    .left(idx_between_30_31_comb_left),
    .out(idx_between_30_31_comb_out),
    .right(idx_between_30_31_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_34_50_reg (
    .clk(idx_between_34_50_reg_clk),
    .done(idx_between_34_50_reg_done),
    .in(idx_between_34_50_reg_in),
    .out(idx_between_34_50_reg_out),
    .reset(idx_between_34_50_reg_reset),
    .write_en(idx_between_34_50_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_34 (
    .left(index_ge_34_left),
    .out(index_ge_34_out),
    .right(index_ge_34_right)
);
std_and # (
    .WIDTH(1)
) idx_between_34_50_comb (
    .left(idx_between_34_50_comb_left),
    .out(idx_between_34_50_comb_out),
    .right(idx_between_34_50_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_7_11_reg (
    .clk(idx_between_7_11_reg_clk),
    .done(idx_between_7_11_reg_done),
    .in(idx_between_7_11_reg_in),
    .out(idx_between_7_11_reg_out),
    .reset(idx_between_7_11_reg_reset),
    .write_en(idx_between_7_11_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_11 (
    .left(index_lt_11_left),
    .out(index_lt_11_out),
    .right(index_lt_11_right)
);
std_and # (
    .WIDTH(1)
) idx_between_7_11_comb (
    .left(idx_between_7_11_comb_left),
    .out(idx_between_7_11_comb_out),
    .right(idx_between_7_11_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_11_27_reg (
    .clk(idx_between_11_27_reg_clk),
    .done(idx_between_11_27_reg_done),
    .in(idx_between_11_27_reg_in),
    .out(idx_between_11_27_reg_out),
    .reset(idx_between_11_27_reg_reset),
    .write_en(idx_between_11_27_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_11 (
    .left(index_ge_11_left),
    .out(index_ge_11_out),
    .right(index_ge_11_right)
);
std_and # (
    .WIDTH(1)
) idx_between_11_27_comb (
    .left(idx_between_11_27_comb_left),
    .out(idx_between_11_27_comb_out),
    .right(idx_between_11_27_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_25_26_reg (
    .clk(idx_between_25_26_reg_clk),
    .done(idx_between_25_26_reg_done),
    .in(idx_between_25_26_reg_in),
    .out(idx_between_25_26_reg_out),
    .reset(idx_between_25_26_reg_reset),
    .write_en(idx_between_25_26_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_25_26_comb (
    .left(idx_between_25_26_comb_left),
    .out(idx_between_25_26_comb_out),
    .right(idx_between_25_26_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_26_27_reg (
    .clk(idx_between_26_27_reg_clk),
    .done(idx_between_26_27_reg_done),
    .in(idx_between_26_27_reg_in),
    .out(idx_between_26_27_reg_out),
    .reset(idx_between_26_27_reg_reset),
    .write_en(idx_between_26_27_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_26_27_comb (
    .left(idx_between_26_27_comb_left),
    .out(idx_between_26_27_comb_out),
    .right(idx_between_26_27_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_3_7_reg (
    .clk(idx_between_3_7_reg_clk),
    .done(idx_between_3_7_reg_done),
    .in(idx_between_3_7_reg_in),
    .out(idx_between_3_7_reg_out),
    .reset(idx_between_3_7_reg_reset),
    .write_en(idx_between_3_7_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_7 (
    .left(index_lt_7_left),
    .out(index_lt_7_out),
    .right(index_lt_7_right)
);
std_and # (
    .WIDTH(1)
) idx_between_3_7_comb (
    .left(idx_between_3_7_comb_left),
    .out(idx_between_3_7_comb_out),
    .right(idx_between_3_7_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_21_22_reg (
    .clk(idx_between_21_22_reg_clk),
    .done(idx_between_21_22_reg_done),
    .in(idx_between_21_22_reg_in),
    .out(idx_between_21_22_reg_out),
    .reset(idx_between_21_22_reg_reset),
    .write_en(idx_between_21_22_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_21_22_comb (
    .left(idx_between_21_22_comb_left),
    .out(idx_between_21_22_comb_out),
    .right(idx_between_21_22_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_31_32_reg (
    .clk(idx_between_31_32_reg_clk),
    .done(idx_between_31_32_reg_done),
    .in(idx_between_31_32_reg_in),
    .out(idx_between_31_32_reg_out),
    .reset(idx_between_31_32_reg_reset),
    .write_en(idx_between_31_32_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_31_32_comb (
    .left(idx_between_31_32_comb_left),
    .out(idx_between_31_32_comb_out),
    .right(idx_between_31_32_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_12_28_reg (
    .clk(idx_between_12_28_reg_clk),
    .done(idx_between_12_28_reg_done),
    .in(idx_between_12_28_reg_in),
    .out(idx_between_12_28_reg_out),
    .reset(idx_between_12_28_reg_reset),
    .write_en(idx_between_12_28_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_12 (
    .left(index_ge_12_left),
    .out(index_ge_12_out),
    .right(index_ge_12_right)
);
std_and # (
    .WIDTH(1)
) idx_between_12_28_comb (
    .left(idx_between_12_28_comb_left),
    .out(idx_between_12_28_comb_out),
    .right(idx_between_12_28_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_27_28_reg (
    .clk(idx_between_27_28_reg_clk),
    .done(idx_between_27_28_reg_done),
    .in(idx_between_27_28_reg_in),
    .out(idx_between_27_28_reg_out),
    .reset(idx_between_27_28_reg_reset),
    .write_en(idx_between_27_28_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_27_28_comb (
    .left(idx_between_27_28_comb_left),
    .out(idx_between_27_28_comb_out),
    .right(idx_between_27_28_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_8_24_reg (
    .clk(idx_between_8_24_reg_clk),
    .done(idx_between_8_24_reg_done),
    .in(idx_between_8_24_reg_in),
    .out(idx_between_8_24_reg_out),
    .reset(idx_between_8_24_reg_reset),
    .write_en(idx_between_8_24_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_8 (
    .left(index_ge_8_left),
    .out(index_ge_8_out),
    .right(index_ge_8_right)
);
std_and # (
    .WIDTH(1)
) idx_between_8_24_comb (
    .left(idx_between_8_24_comb_left),
    .out(idx_between_8_24_comb_out),
    .right(idx_between_8_24_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_4_8_reg (
    .clk(idx_between_4_8_reg_clk),
    .done(idx_between_4_8_reg_done),
    .in(idx_between_4_8_reg_in),
    .out(idx_between_4_8_reg_out),
    .reset(idx_between_4_8_reg_reset),
    .write_en(idx_between_4_8_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_8 (
    .left(index_lt_8_left),
    .out(index_lt_8_out),
    .right(index_lt_8_right)
);
std_and # (
    .WIDTH(1)
) idx_between_4_8_comb (
    .left(idx_between_4_8_comb_left),
    .out(idx_between_4_8_comb_out),
    .right(idx_between_4_8_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_14_18_reg (
    .clk(idx_between_14_18_reg_clk),
    .done(idx_between_14_18_reg_done),
    .in(idx_between_14_18_reg_in),
    .out(idx_between_14_18_reg_out),
    .reset(idx_between_14_18_reg_reset),
    .write_en(idx_between_14_18_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_18 (
    .left(index_lt_18_left),
    .out(index_lt_18_out),
    .right(index_lt_18_right)
);
std_and # (
    .WIDTH(1)
) idx_between_14_18_comb (
    .left(idx_between_14_18_comb_left),
    .out(idx_between_14_18_comb_out),
    .right(idx_between_14_18_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_18_34_reg (
    .clk(idx_between_18_34_reg_clk),
    .done(idx_between_18_34_reg_done),
    .in(idx_between_18_34_reg_in),
    .out(idx_between_18_34_reg_out),
    .reset(idx_between_18_34_reg_reset),
    .write_en(idx_between_18_34_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_18 (
    .left(index_ge_18_left),
    .out(index_ge_18_out),
    .right(index_ge_18_right)
);
std_and # (
    .WIDTH(1)
) idx_between_18_34_comb (
    .left(idx_between_18_34_comb_left),
    .out(idx_between_18_34_comb_out),
    .right(idx_between_18_34_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_10_14_reg (
    .clk(idx_between_10_14_reg_clk),
    .done(idx_between_10_14_reg_done),
    .in(idx_between_10_14_reg_in),
    .out(idx_between_10_14_reg_out),
    .reset(idx_between_10_14_reg_reset),
    .write_en(idx_between_10_14_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_14 (
    .left(index_lt_14_left),
    .out(index_lt_14_out),
    .right(index_lt_14_right)
);
std_and # (
    .WIDTH(1)
) idx_between_10_14_comb (
    .left(idx_between_10_14_comb_left),
    .out(idx_between_10_14_comb_out),
    .right(idx_between_10_14_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_28_29_reg (
    .clk(idx_between_28_29_reg_clk),
    .done(idx_between_28_29_reg_done),
    .in(idx_between_28_29_reg_in),
    .out(idx_between_28_29_reg_out),
    .reset(idx_between_28_29_reg_reset),
    .write_en(idx_between_28_29_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_28_29_comb (
    .left(idx_between_28_29_comb_left),
    .out(idx_between_28_29_comb_out),
    .right(idx_between_28_29_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_9_25_reg (
    .clk(idx_between_9_25_reg_clk),
    .done(idx_between_9_25_reg_done),
    .in(idx_between_9_25_reg_in),
    .out(idx_between_9_25_reg_out),
    .reset(idx_between_9_25_reg_reset),
    .write_en(idx_between_9_25_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_9 (
    .left(index_ge_9_left),
    .out(index_ge_9_out),
    .right(index_ge_9_right)
);
std_and # (
    .WIDTH(1)
) idx_between_9_25_comb (
    .left(idx_between_9_25_comb_left),
    .out(idx_between_9_25_comb_out),
    .right(idx_between_9_25_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_19_35_reg (
    .clk(idx_between_19_35_reg_clk),
    .done(idx_between_19_35_reg_done),
    .in(idx_between_19_35_reg_in),
    .out(idx_between_19_35_reg_out),
    .reset(idx_between_19_35_reg_reset),
    .write_en(idx_between_19_35_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_19 (
    .left(index_ge_19_left),
    .out(index_ge_19_out),
    .right(index_ge_19_right)
);
std_and # (
    .WIDTH(1)
) idx_between_19_35_comb (
    .left(idx_between_19_35_comb_left),
    .out(idx_between_19_35_comb_out),
    .right(idx_between_19_35_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_6_10_reg (
    .clk(idx_between_6_10_reg_clk),
    .done(idx_between_6_10_reg_done),
    .in(idx_between_6_10_reg_in),
    .out(idx_between_6_10_reg_out),
    .reset(idx_between_6_10_reg_reset),
    .write_en(idx_between_6_10_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_10 (
    .left(index_lt_10_left),
    .out(index_lt_10_out),
    .right(index_lt_10_right)
);
std_and # (
    .WIDTH(1)
) idx_between_6_10_comb (
    .left(idx_between_6_10_comb_left),
    .out(idx_between_6_10_comb_out),
    .right(idx_between_6_10_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_15_31_reg (
    .clk(idx_between_15_31_reg_clk),
    .done(idx_between_15_31_reg_done),
    .in(idx_between_15_31_reg_in),
    .out(idx_between_15_31_reg_out),
    .reset(idx_between_15_31_reg_reset),
    .write_en(idx_between_15_31_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_15 (
    .left(index_ge_15_left),
    .out(index_ge_15_out),
    .right(index_ge_15_right)
);
std_and # (
    .WIDTH(1)
) idx_between_15_31_comb (
    .left(idx_between_15_31_comb_left),
    .out(idx_between_15_31_comb_out),
    .right(idx_between_15_31_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_29_30_reg (
    .clk(idx_between_29_30_reg_clk),
    .done(idx_between_29_30_reg_done),
    .in(idx_between_29_30_reg_in),
    .out(idx_between_29_30_reg_out),
    .reset(idx_between_29_30_reg_reset),
    .write_en(idx_between_29_30_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_29_30_comb (
    .left(idx_between_29_30_comb_left),
    .out(idx_between_29_30_comb_out),
    .right(idx_between_29_30_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_11_15_reg (
    .clk(idx_between_11_15_reg_clk),
    .done(idx_between_11_15_reg_done),
    .in(idx_between_11_15_reg_in),
    .out(idx_between_11_15_reg_out),
    .reset(idx_between_11_15_reg_reset),
    .write_en(idx_between_11_15_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_15 (
    .left(index_lt_15_left),
    .out(index_lt_15_out),
    .right(index_lt_15_right)
);
std_and # (
    .WIDTH(1)
) idx_between_11_15_comb (
    .left(idx_between_11_15_comb_left),
    .out(idx_between_11_15_comb_out),
    .right(idx_between_11_15_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_35_36_reg (
    .clk(idx_between_35_36_reg_clk),
    .done(idx_between_35_36_reg_done),
    .in(idx_between_35_36_reg_in),
    .out(idx_between_35_36_reg_out),
    .reset(idx_between_35_36_reg_reset),
    .write_en(idx_between_35_36_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_36 (
    .left(index_lt_36_left),
    .out(index_lt_36_out),
    .right(index_lt_36_right)
);
std_and # (
    .WIDTH(1)
) idx_between_35_36_comb (
    .left(idx_between_35_36_comb_left),
    .out(idx_between_35_36_comb_out),
    .right(idx_between_35_36_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_12_16_reg (
    .clk(idx_between_12_16_reg_clk),
    .done(idx_between_12_16_reg_done),
    .in(idx_between_12_16_reg_in),
    .out(idx_between_12_16_reg_out),
    .reset(idx_between_12_16_reg_reset),
    .write_en(idx_between_12_16_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_12_16_comb (
    .left(idx_between_12_16_comb_left),
    .out(idx_between_12_16_comb_out),
    .right(idx_between_12_16_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_16_32_reg (
    .clk(idx_between_16_32_reg_clk),
    .done(idx_between_16_32_reg_done),
    .in(idx_between_16_32_reg_in),
    .out(idx_between_16_32_reg_out),
    .reset(idx_between_16_32_reg_reset),
    .write_en(idx_between_16_32_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_16_32_comb (
    .left(idx_between_16_32_comb_left),
    .out(idx_between_16_32_comb_out),
    .right(idx_between_16_32_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_26_42_reg (
    .clk(idx_between_26_42_reg_clk),
    .done(idx_between_26_42_reg_done),
    .in(idx_between_26_42_reg_in),
    .out(idx_between_26_42_reg_out),
    .reset(idx_between_26_42_reg_reset),
    .write_en(idx_between_26_42_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_26_42_comb (
    .left(idx_between_26_42_comb_left),
    .out(idx_between_26_42_comb_out),
    .right(idx_between_26_42_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_8_12_reg (
    .clk(idx_between_8_12_reg_clk),
    .done(idx_between_8_12_reg_done),
    .in(idx_between_8_12_reg_in),
    .out(idx_between_8_12_reg_out),
    .reset(idx_between_8_12_reg_reset),
    .write_en(idx_between_8_12_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_12 (
    .left(index_lt_12_left),
    .out(index_lt_12_out),
    .right(index_lt_12_right)
);
std_and # (
    .WIDTH(1)
) idx_between_8_12_comb (
    .left(idx_between_8_12_comb_left),
    .out(idx_between_8_12_comb_out),
    .right(idx_between_8_12_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_22_38_reg (
    .clk(idx_between_22_38_reg_clk),
    .done(idx_between_22_38_reg_done),
    .in(idx_between_22_38_reg_in),
    .out(idx_between_22_38_reg_out),
    .reset(idx_between_22_38_reg_reset),
    .write_en(idx_between_22_38_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_38 (
    .left(index_lt_38_left),
    .out(index_lt_38_out),
    .right(index_lt_38_right)
);
std_and # (
    .WIDTH(1)
) idx_between_22_38_comb (
    .left(idx_between_22_38_comb_left),
    .out(idx_between_22_38_comb_out),
    .right(idx_between_22_38_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_36_37_reg (
    .clk(idx_between_36_37_reg_clk),
    .done(idx_between_36_37_reg_done),
    .in(idx_between_36_37_reg_in),
    .out(idx_between_36_37_reg_out),
    .reset(idx_between_36_37_reg_reset),
    .write_en(idx_between_36_37_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_36 (
    .left(index_ge_36_left),
    .out(index_ge_36_out),
    .right(index_ge_36_right)
);
std_and # (
    .WIDTH(1)
) idx_between_36_37_comb (
    .left(idx_between_36_37_comb_left),
    .out(idx_between_36_37_comb_out),
    .right(idx_between_36_37_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_17_33_reg (
    .clk(idx_between_17_33_reg_clk),
    .done(idx_between_17_33_reg_done),
    .in(idx_between_17_33_reg_in),
    .out(idx_between_17_33_reg_out),
    .reset(idx_between_17_33_reg_reset),
    .write_en(idx_between_17_33_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_17_33_comb (
    .left(idx_between_17_33_comb_left),
    .out(idx_between_17_33_comb_out),
    .right(idx_between_17_33_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_32_33_reg (
    .clk(idx_between_32_33_reg_clk),
    .done(idx_between_32_33_reg_done),
    .in(idx_between_32_33_reg_in),
    .out(idx_between_32_33_reg_out),
    .reset(idx_between_32_33_reg_reset),
    .write_en(idx_between_32_33_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_32_33_comb (
    .left(idx_between_32_33_comb_left),
    .out(idx_between_32_33_comb_out),
    .right(idx_between_32_33_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_13_29_reg (
    .clk(idx_between_13_29_reg_clk),
    .done(idx_between_13_29_reg_done),
    .in(idx_between_13_29_reg_in),
    .out(idx_between_13_29_reg_out),
    .reset(idx_between_13_29_reg_reset),
    .write_en(idx_between_13_29_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_13_29_comb (
    .left(idx_between_13_29_comb_left),
    .out(idx_between_13_29_comb_out),
    .right(idx_between_13_29_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_18_22_reg (
    .clk(idx_between_18_22_reg_clk),
    .done(idx_between_18_22_reg_done),
    .in(idx_between_18_22_reg_in),
    .out(idx_between_18_22_reg_out),
    .reset(idx_between_18_22_reg_reset),
    .write_en(idx_between_18_22_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_18_22_comb (
    .left(idx_between_18_22_comb_left),
    .out(idx_between_18_22_comb_out),
    .right(idx_between_18_22_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_9_13_reg (
    .clk(idx_between_9_13_reg_clk),
    .done(idx_between_9_13_reg_done),
    .in(idx_between_9_13_reg_in),
    .out(idx_between_9_13_reg_out),
    .reset(idx_between_9_13_reg_reset),
    .write_en(idx_between_9_13_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_13 (
    .left(index_lt_13_left),
    .out(index_lt_13_out),
    .right(index_lt_13_right)
);
std_and # (
    .WIDTH(1)
) idx_between_9_13_comb (
    .left(idx_between_9_13_comb_left),
    .out(idx_between_9_13_comb_out),
    .right(idx_between_9_13_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_19_23_reg (
    .clk(idx_between_19_23_reg_clk),
    .done(idx_between_19_23_reg_done),
    .in(idx_between_19_23_reg_in),
    .out(idx_between_19_23_reg_out),
    .reset(idx_between_19_23_reg_reset),
    .write_en(idx_between_19_23_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_19_23_comb (
    .left(idx_between_19_23_comb_left),
    .out(idx_between_19_23_comb_out),
    .right(idx_between_19_23_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_23_39_reg (
    .clk(idx_between_23_39_reg_clk),
    .done(idx_between_23_39_reg_done),
    .in(idx_between_23_39_reg_in),
    .out(idx_between_23_39_reg_out),
    .reset(idx_between_23_39_reg_reset),
    .write_en(idx_between_23_39_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_23_39_comb (
    .left(idx_between_23_39_comb_left),
    .out(idx_between_23_39_comb_out),
    .right(idx_between_23_39_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_37_38_reg (
    .clk(idx_between_37_38_reg_clk),
    .done(idx_between_37_38_reg_done),
    .in(idx_between_37_38_reg_in),
    .out(idx_between_37_38_reg_out),
    .reset(idx_between_37_38_reg_reset),
    .write_en(idx_between_37_38_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_37 (
    .left(index_ge_37_left),
    .out(index_ge_37_out),
    .right(index_ge_37_right)
);
std_and # (
    .WIDTH(1)
) idx_between_37_38_comb (
    .left(idx_between_37_38_comb_left),
    .out(idx_between_37_38_comb_out),
    .right(idx_between_37_38_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_28_44_reg (
    .clk(idx_between_28_44_reg_clk),
    .done(idx_between_28_44_reg_done),
    .in(idx_between_28_44_reg_in),
    .out(idx_between_28_44_reg_out),
    .reset(idx_between_28_44_reg_reset),
    .write_en(idx_between_28_44_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_44 (
    .left(index_lt_44_left),
    .out(index_lt_44_out),
    .right(index_lt_44_right)
);
std_and # (
    .WIDTH(1)
) idx_between_28_44_comb (
    .left(idx_between_28_44_comb_left),
    .out(idx_between_28_44_comb_out),
    .right(idx_between_28_44_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_15_19_reg (
    .clk(idx_between_15_19_reg_clk),
    .done(idx_between_15_19_reg_done),
    .in(idx_between_15_19_reg_in),
    .out(idx_between_15_19_reg_out),
    .reset(idx_between_15_19_reg_reset),
    .write_en(idx_between_15_19_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_15_19_comb (
    .left(idx_between_15_19_comb_left),
    .out(idx_between_15_19_comb_out),
    .right(idx_between_15_19_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_33_34_reg (
    .clk(idx_between_33_34_reg_clk),
    .done(idx_between_33_34_reg_done),
    .in(idx_between_33_34_reg_in),
    .out(idx_between_33_34_reg_out),
    .reset(idx_between_33_34_reg_reset),
    .write_en(idx_between_33_34_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_33_34_comb (
    .left(idx_between_33_34_comb_left),
    .out(idx_between_33_34_comb_out),
    .right(idx_between_33_34_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_43_44_reg (
    .clk(idx_between_43_44_reg_clk),
    .done(idx_between_43_44_reg_done),
    .in(idx_between_43_44_reg_in),
    .out(idx_between_43_44_reg_out),
    .reset(idx_between_43_44_reg_reset),
    .write_en(idx_between_43_44_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_43 (
    .left(index_ge_43_left),
    .out(index_ge_43_out),
    .right(index_ge_43_right)
);
std_and # (
    .WIDTH(1)
) idx_between_43_44_comb (
    .left(idx_between_43_44_comb_left),
    .out(idx_between_43_44_comb_out),
    .right(idx_between_43_44_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_24_40_reg (
    .clk(idx_between_24_40_reg_clk),
    .done(idx_between_24_40_reg_done),
    .in(idx_between_24_40_reg_in),
    .out(idx_between_24_40_reg_out),
    .reset(idx_between_24_40_reg_reset),
    .write_en(idx_between_24_40_reg_write_en)
);
std_lt # (
    .WIDTH(6)
) index_lt_40 (
    .left(index_lt_40_left),
    .out(index_lt_40_out),
    .right(index_lt_40_right)
);
std_and # (
    .WIDTH(1)
) idx_between_24_40_comb (
    .left(idx_between_24_40_comb_left),
    .out(idx_between_24_40_comb_out),
    .right(idx_between_24_40_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_39_40_reg (
    .clk(idx_between_39_40_reg_clk),
    .done(idx_between_39_40_reg_done),
    .in(idx_between_39_40_reg_in),
    .out(idx_between_39_40_reg_out),
    .reset(idx_between_39_40_reg_reset),
    .write_en(idx_between_39_40_reg_write_en)
);
std_ge # (
    .WIDTH(6)
) index_ge_39 (
    .left(index_ge_39_left),
    .out(index_ge_39_out),
    .right(index_ge_39_right)
);
std_and # (
    .WIDTH(1)
) idx_between_39_40_comb (
    .left(idx_between_39_40_comb_left),
    .out(idx_between_39_40_comb_out),
    .right(idx_between_39_40_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_20_36_reg (
    .clk(idx_between_20_36_reg_clk),
    .done(idx_between_20_36_reg_done),
    .in(idx_between_20_36_reg_in),
    .out(idx_between_20_36_reg_out),
    .reset(idx_between_20_36_reg_reset),
    .write_en(idx_between_20_36_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_20_36_comb (
    .left(idx_between_20_36_comb_left),
    .out(idx_between_20_36_comb_out),
    .right(idx_between_20_36_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_34_35_reg (
    .clk(idx_between_34_35_reg_clk),
    .done(idx_between_34_35_reg_done),
    .in(idx_between_34_35_reg_in),
    .out(idx_between_34_35_reg_out),
    .reset(idx_between_34_35_reg_reset),
    .write_en(idx_between_34_35_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_34_35_comb (
    .left(idx_between_34_35_comb_left),
    .out(idx_between_34_35_comb_out),
    .right(idx_between_34_35_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_2_18_reg (
    .clk(idx_between_2_18_reg_clk),
    .done(idx_between_2_18_reg_done),
    .in(idx_between_2_18_reg_in),
    .out(idx_between_2_18_reg_out),
    .reset(idx_between_2_18_reg_reset),
    .write_en(idx_between_2_18_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_2_18_comb (
    .left(idx_between_2_18_comb_left),
    .out(idx_between_2_18_comb_out),
    .right(idx_between_2_18_comb_right)
);
std_reg # (
    .WIDTH(1)
) cond (
    .clk(cond_clk),
    .done(cond_done),
    .in(cond_in),
    .out(cond_out),
    .reset(cond_reset),
    .write_en(cond_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire (
    .in(cond_wire_in),
    .out(cond_wire_out)
);
std_reg # (
    .WIDTH(1)
) cond0 (
    .clk(cond0_clk),
    .done(cond0_done),
    .in(cond0_in),
    .out(cond0_out),
    .reset(cond0_reset),
    .write_en(cond0_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire0 (
    .in(cond_wire0_in),
    .out(cond_wire0_out)
);
std_reg # (
    .WIDTH(1)
) cond1 (
    .clk(cond1_clk),
    .done(cond1_done),
    .in(cond1_in),
    .out(cond1_out),
    .reset(cond1_reset),
    .write_en(cond1_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1 (
    .in(cond_wire1_in),
    .out(cond_wire1_out)
);
std_reg # (
    .WIDTH(1)
) cond2 (
    .clk(cond2_clk),
    .done(cond2_done),
    .in(cond2_in),
    .out(cond2_out),
    .reset(cond2_reset),
    .write_en(cond2_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire2 (
    .in(cond_wire2_in),
    .out(cond_wire2_out)
);
std_reg # (
    .WIDTH(1)
) cond3 (
    .clk(cond3_clk),
    .done(cond3_done),
    .in(cond3_in),
    .out(cond3_out),
    .reset(cond3_reset),
    .write_en(cond3_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire3 (
    .in(cond_wire3_in),
    .out(cond_wire3_out)
);
std_reg # (
    .WIDTH(1)
) cond4 (
    .clk(cond4_clk),
    .done(cond4_done),
    .in(cond4_in),
    .out(cond4_out),
    .reset(cond4_reset),
    .write_en(cond4_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire4 (
    .in(cond_wire4_in),
    .out(cond_wire4_out)
);
std_reg # (
    .WIDTH(1)
) cond5 (
    .clk(cond5_clk),
    .done(cond5_done),
    .in(cond5_in),
    .out(cond5_out),
    .reset(cond5_reset),
    .write_en(cond5_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire5 (
    .in(cond_wire5_in),
    .out(cond_wire5_out)
);
std_reg # (
    .WIDTH(1)
) cond6 (
    .clk(cond6_clk),
    .done(cond6_done),
    .in(cond6_in),
    .out(cond6_out),
    .reset(cond6_reset),
    .write_en(cond6_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire6 (
    .in(cond_wire6_in),
    .out(cond_wire6_out)
);
std_reg # (
    .WIDTH(1)
) cond7 (
    .clk(cond7_clk),
    .done(cond7_done),
    .in(cond7_in),
    .out(cond7_out),
    .reset(cond7_reset),
    .write_en(cond7_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire7 (
    .in(cond_wire7_in),
    .out(cond_wire7_out)
);
std_reg # (
    .WIDTH(1)
) cond8 (
    .clk(cond8_clk),
    .done(cond8_done),
    .in(cond8_in),
    .out(cond8_out),
    .reset(cond8_reset),
    .write_en(cond8_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire8 (
    .in(cond_wire8_in),
    .out(cond_wire8_out)
);
std_reg # (
    .WIDTH(1)
) cond9 (
    .clk(cond9_clk),
    .done(cond9_done),
    .in(cond9_in),
    .out(cond9_out),
    .reset(cond9_reset),
    .write_en(cond9_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire9 (
    .in(cond_wire9_in),
    .out(cond_wire9_out)
);
std_reg # (
    .WIDTH(1)
) cond10 (
    .clk(cond10_clk),
    .done(cond10_done),
    .in(cond10_in),
    .out(cond10_out),
    .reset(cond10_reset),
    .write_en(cond10_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire10 (
    .in(cond_wire10_in),
    .out(cond_wire10_out)
);
std_reg # (
    .WIDTH(1)
) cond11 (
    .clk(cond11_clk),
    .done(cond11_done),
    .in(cond11_in),
    .out(cond11_out),
    .reset(cond11_reset),
    .write_en(cond11_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire11 (
    .in(cond_wire11_in),
    .out(cond_wire11_out)
);
std_reg # (
    .WIDTH(1)
) cond12 (
    .clk(cond12_clk),
    .done(cond12_done),
    .in(cond12_in),
    .out(cond12_out),
    .reset(cond12_reset),
    .write_en(cond12_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire12 (
    .in(cond_wire12_in),
    .out(cond_wire12_out)
);
std_reg # (
    .WIDTH(1)
) cond13 (
    .clk(cond13_clk),
    .done(cond13_done),
    .in(cond13_in),
    .out(cond13_out),
    .reset(cond13_reset),
    .write_en(cond13_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire13 (
    .in(cond_wire13_in),
    .out(cond_wire13_out)
);
std_reg # (
    .WIDTH(1)
) cond14 (
    .clk(cond14_clk),
    .done(cond14_done),
    .in(cond14_in),
    .out(cond14_out),
    .reset(cond14_reset),
    .write_en(cond14_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire14 (
    .in(cond_wire14_in),
    .out(cond_wire14_out)
);
std_reg # (
    .WIDTH(1)
) cond15 (
    .clk(cond15_clk),
    .done(cond15_done),
    .in(cond15_in),
    .out(cond15_out),
    .reset(cond15_reset),
    .write_en(cond15_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire15 (
    .in(cond_wire15_in),
    .out(cond_wire15_out)
);
std_reg # (
    .WIDTH(1)
) cond16 (
    .clk(cond16_clk),
    .done(cond16_done),
    .in(cond16_in),
    .out(cond16_out),
    .reset(cond16_reset),
    .write_en(cond16_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire16 (
    .in(cond_wire16_in),
    .out(cond_wire16_out)
);
std_reg # (
    .WIDTH(1)
) cond17 (
    .clk(cond17_clk),
    .done(cond17_done),
    .in(cond17_in),
    .out(cond17_out),
    .reset(cond17_reset),
    .write_en(cond17_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire17 (
    .in(cond_wire17_in),
    .out(cond_wire17_out)
);
std_reg # (
    .WIDTH(1)
) cond18 (
    .clk(cond18_clk),
    .done(cond18_done),
    .in(cond18_in),
    .out(cond18_out),
    .reset(cond18_reset),
    .write_en(cond18_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire18 (
    .in(cond_wire18_in),
    .out(cond_wire18_out)
);
std_reg # (
    .WIDTH(1)
) cond19 (
    .clk(cond19_clk),
    .done(cond19_done),
    .in(cond19_in),
    .out(cond19_out),
    .reset(cond19_reset),
    .write_en(cond19_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire19 (
    .in(cond_wire19_in),
    .out(cond_wire19_out)
);
std_reg # (
    .WIDTH(1)
) cond20 (
    .clk(cond20_clk),
    .done(cond20_done),
    .in(cond20_in),
    .out(cond20_out),
    .reset(cond20_reset),
    .write_en(cond20_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire20 (
    .in(cond_wire20_in),
    .out(cond_wire20_out)
);
std_reg # (
    .WIDTH(1)
) cond21 (
    .clk(cond21_clk),
    .done(cond21_done),
    .in(cond21_in),
    .out(cond21_out),
    .reset(cond21_reset),
    .write_en(cond21_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire21 (
    .in(cond_wire21_in),
    .out(cond_wire21_out)
);
std_reg # (
    .WIDTH(1)
) cond22 (
    .clk(cond22_clk),
    .done(cond22_done),
    .in(cond22_in),
    .out(cond22_out),
    .reset(cond22_reset),
    .write_en(cond22_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire22 (
    .in(cond_wire22_in),
    .out(cond_wire22_out)
);
std_reg # (
    .WIDTH(1)
) cond23 (
    .clk(cond23_clk),
    .done(cond23_done),
    .in(cond23_in),
    .out(cond23_out),
    .reset(cond23_reset),
    .write_en(cond23_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire23 (
    .in(cond_wire23_in),
    .out(cond_wire23_out)
);
std_reg # (
    .WIDTH(1)
) cond24 (
    .clk(cond24_clk),
    .done(cond24_done),
    .in(cond24_in),
    .out(cond24_out),
    .reset(cond24_reset),
    .write_en(cond24_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire24 (
    .in(cond_wire24_in),
    .out(cond_wire24_out)
);
std_reg # (
    .WIDTH(1)
) cond25 (
    .clk(cond25_clk),
    .done(cond25_done),
    .in(cond25_in),
    .out(cond25_out),
    .reset(cond25_reset),
    .write_en(cond25_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire25 (
    .in(cond_wire25_in),
    .out(cond_wire25_out)
);
std_reg # (
    .WIDTH(1)
) cond26 (
    .clk(cond26_clk),
    .done(cond26_done),
    .in(cond26_in),
    .out(cond26_out),
    .reset(cond26_reset),
    .write_en(cond26_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire26 (
    .in(cond_wire26_in),
    .out(cond_wire26_out)
);
std_reg # (
    .WIDTH(1)
) cond27 (
    .clk(cond27_clk),
    .done(cond27_done),
    .in(cond27_in),
    .out(cond27_out),
    .reset(cond27_reset),
    .write_en(cond27_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire27 (
    .in(cond_wire27_in),
    .out(cond_wire27_out)
);
std_reg # (
    .WIDTH(1)
) cond28 (
    .clk(cond28_clk),
    .done(cond28_done),
    .in(cond28_in),
    .out(cond28_out),
    .reset(cond28_reset),
    .write_en(cond28_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire28 (
    .in(cond_wire28_in),
    .out(cond_wire28_out)
);
std_reg # (
    .WIDTH(1)
) cond29 (
    .clk(cond29_clk),
    .done(cond29_done),
    .in(cond29_in),
    .out(cond29_out),
    .reset(cond29_reset),
    .write_en(cond29_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire29 (
    .in(cond_wire29_in),
    .out(cond_wire29_out)
);
std_reg # (
    .WIDTH(1)
) cond30 (
    .clk(cond30_clk),
    .done(cond30_done),
    .in(cond30_in),
    .out(cond30_out),
    .reset(cond30_reset),
    .write_en(cond30_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire30 (
    .in(cond_wire30_in),
    .out(cond_wire30_out)
);
std_reg # (
    .WIDTH(1)
) cond31 (
    .clk(cond31_clk),
    .done(cond31_done),
    .in(cond31_in),
    .out(cond31_out),
    .reset(cond31_reset),
    .write_en(cond31_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire31 (
    .in(cond_wire31_in),
    .out(cond_wire31_out)
);
std_reg # (
    .WIDTH(1)
) cond32 (
    .clk(cond32_clk),
    .done(cond32_done),
    .in(cond32_in),
    .out(cond32_out),
    .reset(cond32_reset),
    .write_en(cond32_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire32 (
    .in(cond_wire32_in),
    .out(cond_wire32_out)
);
std_reg # (
    .WIDTH(1)
) cond33 (
    .clk(cond33_clk),
    .done(cond33_done),
    .in(cond33_in),
    .out(cond33_out),
    .reset(cond33_reset),
    .write_en(cond33_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire33 (
    .in(cond_wire33_in),
    .out(cond_wire33_out)
);
std_reg # (
    .WIDTH(1)
) cond34 (
    .clk(cond34_clk),
    .done(cond34_done),
    .in(cond34_in),
    .out(cond34_out),
    .reset(cond34_reset),
    .write_en(cond34_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire34 (
    .in(cond_wire34_in),
    .out(cond_wire34_out)
);
std_reg # (
    .WIDTH(1)
) cond35 (
    .clk(cond35_clk),
    .done(cond35_done),
    .in(cond35_in),
    .out(cond35_out),
    .reset(cond35_reset),
    .write_en(cond35_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire35 (
    .in(cond_wire35_in),
    .out(cond_wire35_out)
);
std_reg # (
    .WIDTH(1)
) cond36 (
    .clk(cond36_clk),
    .done(cond36_done),
    .in(cond36_in),
    .out(cond36_out),
    .reset(cond36_reset),
    .write_en(cond36_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire36 (
    .in(cond_wire36_in),
    .out(cond_wire36_out)
);
std_reg # (
    .WIDTH(1)
) cond37 (
    .clk(cond37_clk),
    .done(cond37_done),
    .in(cond37_in),
    .out(cond37_out),
    .reset(cond37_reset),
    .write_en(cond37_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire37 (
    .in(cond_wire37_in),
    .out(cond_wire37_out)
);
std_reg # (
    .WIDTH(1)
) cond38 (
    .clk(cond38_clk),
    .done(cond38_done),
    .in(cond38_in),
    .out(cond38_out),
    .reset(cond38_reset),
    .write_en(cond38_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire38 (
    .in(cond_wire38_in),
    .out(cond_wire38_out)
);
std_reg # (
    .WIDTH(1)
) cond39 (
    .clk(cond39_clk),
    .done(cond39_done),
    .in(cond39_in),
    .out(cond39_out),
    .reset(cond39_reset),
    .write_en(cond39_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire39 (
    .in(cond_wire39_in),
    .out(cond_wire39_out)
);
std_reg # (
    .WIDTH(1)
) cond40 (
    .clk(cond40_clk),
    .done(cond40_done),
    .in(cond40_in),
    .out(cond40_out),
    .reset(cond40_reset),
    .write_en(cond40_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire40 (
    .in(cond_wire40_in),
    .out(cond_wire40_out)
);
std_reg # (
    .WIDTH(1)
) cond41 (
    .clk(cond41_clk),
    .done(cond41_done),
    .in(cond41_in),
    .out(cond41_out),
    .reset(cond41_reset),
    .write_en(cond41_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire41 (
    .in(cond_wire41_in),
    .out(cond_wire41_out)
);
std_reg # (
    .WIDTH(1)
) cond42 (
    .clk(cond42_clk),
    .done(cond42_done),
    .in(cond42_in),
    .out(cond42_out),
    .reset(cond42_reset),
    .write_en(cond42_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire42 (
    .in(cond_wire42_in),
    .out(cond_wire42_out)
);
std_reg # (
    .WIDTH(1)
) cond43 (
    .clk(cond43_clk),
    .done(cond43_done),
    .in(cond43_in),
    .out(cond43_out),
    .reset(cond43_reset),
    .write_en(cond43_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire43 (
    .in(cond_wire43_in),
    .out(cond_wire43_out)
);
std_reg # (
    .WIDTH(1)
) cond44 (
    .clk(cond44_clk),
    .done(cond44_done),
    .in(cond44_in),
    .out(cond44_out),
    .reset(cond44_reset),
    .write_en(cond44_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire44 (
    .in(cond_wire44_in),
    .out(cond_wire44_out)
);
std_reg # (
    .WIDTH(1)
) cond45 (
    .clk(cond45_clk),
    .done(cond45_done),
    .in(cond45_in),
    .out(cond45_out),
    .reset(cond45_reset),
    .write_en(cond45_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire45 (
    .in(cond_wire45_in),
    .out(cond_wire45_out)
);
std_reg # (
    .WIDTH(1)
) cond46 (
    .clk(cond46_clk),
    .done(cond46_done),
    .in(cond46_in),
    .out(cond46_out),
    .reset(cond46_reset),
    .write_en(cond46_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire46 (
    .in(cond_wire46_in),
    .out(cond_wire46_out)
);
std_reg # (
    .WIDTH(1)
) cond47 (
    .clk(cond47_clk),
    .done(cond47_done),
    .in(cond47_in),
    .out(cond47_out),
    .reset(cond47_reset),
    .write_en(cond47_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire47 (
    .in(cond_wire47_in),
    .out(cond_wire47_out)
);
std_reg # (
    .WIDTH(1)
) cond48 (
    .clk(cond48_clk),
    .done(cond48_done),
    .in(cond48_in),
    .out(cond48_out),
    .reset(cond48_reset),
    .write_en(cond48_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire48 (
    .in(cond_wire48_in),
    .out(cond_wire48_out)
);
std_reg # (
    .WIDTH(1)
) cond49 (
    .clk(cond49_clk),
    .done(cond49_done),
    .in(cond49_in),
    .out(cond49_out),
    .reset(cond49_reset),
    .write_en(cond49_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire49 (
    .in(cond_wire49_in),
    .out(cond_wire49_out)
);
std_reg # (
    .WIDTH(1)
) cond50 (
    .clk(cond50_clk),
    .done(cond50_done),
    .in(cond50_in),
    .out(cond50_out),
    .reset(cond50_reset),
    .write_en(cond50_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire50 (
    .in(cond_wire50_in),
    .out(cond_wire50_out)
);
std_reg # (
    .WIDTH(1)
) cond51 (
    .clk(cond51_clk),
    .done(cond51_done),
    .in(cond51_in),
    .out(cond51_out),
    .reset(cond51_reset),
    .write_en(cond51_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire51 (
    .in(cond_wire51_in),
    .out(cond_wire51_out)
);
std_reg # (
    .WIDTH(1)
) cond52 (
    .clk(cond52_clk),
    .done(cond52_done),
    .in(cond52_in),
    .out(cond52_out),
    .reset(cond52_reset),
    .write_en(cond52_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire52 (
    .in(cond_wire52_in),
    .out(cond_wire52_out)
);
std_reg # (
    .WIDTH(1)
) cond53 (
    .clk(cond53_clk),
    .done(cond53_done),
    .in(cond53_in),
    .out(cond53_out),
    .reset(cond53_reset),
    .write_en(cond53_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire53 (
    .in(cond_wire53_in),
    .out(cond_wire53_out)
);
std_reg # (
    .WIDTH(1)
) cond54 (
    .clk(cond54_clk),
    .done(cond54_done),
    .in(cond54_in),
    .out(cond54_out),
    .reset(cond54_reset),
    .write_en(cond54_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire54 (
    .in(cond_wire54_in),
    .out(cond_wire54_out)
);
std_reg # (
    .WIDTH(1)
) cond55 (
    .clk(cond55_clk),
    .done(cond55_done),
    .in(cond55_in),
    .out(cond55_out),
    .reset(cond55_reset),
    .write_en(cond55_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire55 (
    .in(cond_wire55_in),
    .out(cond_wire55_out)
);
std_reg # (
    .WIDTH(1)
) cond56 (
    .clk(cond56_clk),
    .done(cond56_done),
    .in(cond56_in),
    .out(cond56_out),
    .reset(cond56_reset),
    .write_en(cond56_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire56 (
    .in(cond_wire56_in),
    .out(cond_wire56_out)
);
std_reg # (
    .WIDTH(1)
) cond57 (
    .clk(cond57_clk),
    .done(cond57_done),
    .in(cond57_in),
    .out(cond57_out),
    .reset(cond57_reset),
    .write_en(cond57_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire57 (
    .in(cond_wire57_in),
    .out(cond_wire57_out)
);
std_reg # (
    .WIDTH(1)
) cond58 (
    .clk(cond58_clk),
    .done(cond58_done),
    .in(cond58_in),
    .out(cond58_out),
    .reset(cond58_reset),
    .write_en(cond58_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire58 (
    .in(cond_wire58_in),
    .out(cond_wire58_out)
);
std_reg # (
    .WIDTH(1)
) cond59 (
    .clk(cond59_clk),
    .done(cond59_done),
    .in(cond59_in),
    .out(cond59_out),
    .reset(cond59_reset),
    .write_en(cond59_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire59 (
    .in(cond_wire59_in),
    .out(cond_wire59_out)
);
std_reg # (
    .WIDTH(1)
) cond60 (
    .clk(cond60_clk),
    .done(cond60_done),
    .in(cond60_in),
    .out(cond60_out),
    .reset(cond60_reset),
    .write_en(cond60_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire60 (
    .in(cond_wire60_in),
    .out(cond_wire60_out)
);
std_reg # (
    .WIDTH(1)
) cond61 (
    .clk(cond61_clk),
    .done(cond61_done),
    .in(cond61_in),
    .out(cond61_out),
    .reset(cond61_reset),
    .write_en(cond61_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire61 (
    .in(cond_wire61_in),
    .out(cond_wire61_out)
);
std_reg # (
    .WIDTH(1)
) cond62 (
    .clk(cond62_clk),
    .done(cond62_done),
    .in(cond62_in),
    .out(cond62_out),
    .reset(cond62_reset),
    .write_en(cond62_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire62 (
    .in(cond_wire62_in),
    .out(cond_wire62_out)
);
std_reg # (
    .WIDTH(1)
) cond63 (
    .clk(cond63_clk),
    .done(cond63_done),
    .in(cond63_in),
    .out(cond63_out),
    .reset(cond63_reset),
    .write_en(cond63_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire63 (
    .in(cond_wire63_in),
    .out(cond_wire63_out)
);
std_reg # (
    .WIDTH(1)
) cond64 (
    .clk(cond64_clk),
    .done(cond64_done),
    .in(cond64_in),
    .out(cond64_out),
    .reset(cond64_reset),
    .write_en(cond64_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire64 (
    .in(cond_wire64_in),
    .out(cond_wire64_out)
);
std_reg # (
    .WIDTH(1)
) cond65 (
    .clk(cond65_clk),
    .done(cond65_done),
    .in(cond65_in),
    .out(cond65_out),
    .reset(cond65_reset),
    .write_en(cond65_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire65 (
    .in(cond_wire65_in),
    .out(cond_wire65_out)
);
std_reg # (
    .WIDTH(1)
) cond66 (
    .clk(cond66_clk),
    .done(cond66_done),
    .in(cond66_in),
    .out(cond66_out),
    .reset(cond66_reset),
    .write_en(cond66_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire66 (
    .in(cond_wire66_in),
    .out(cond_wire66_out)
);
std_reg # (
    .WIDTH(1)
) cond67 (
    .clk(cond67_clk),
    .done(cond67_done),
    .in(cond67_in),
    .out(cond67_out),
    .reset(cond67_reset),
    .write_en(cond67_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire67 (
    .in(cond_wire67_in),
    .out(cond_wire67_out)
);
std_reg # (
    .WIDTH(1)
) cond68 (
    .clk(cond68_clk),
    .done(cond68_done),
    .in(cond68_in),
    .out(cond68_out),
    .reset(cond68_reset),
    .write_en(cond68_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire68 (
    .in(cond_wire68_in),
    .out(cond_wire68_out)
);
std_reg # (
    .WIDTH(1)
) cond69 (
    .clk(cond69_clk),
    .done(cond69_done),
    .in(cond69_in),
    .out(cond69_out),
    .reset(cond69_reset),
    .write_en(cond69_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire69 (
    .in(cond_wire69_in),
    .out(cond_wire69_out)
);
std_reg # (
    .WIDTH(1)
) cond70 (
    .clk(cond70_clk),
    .done(cond70_done),
    .in(cond70_in),
    .out(cond70_out),
    .reset(cond70_reset),
    .write_en(cond70_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire70 (
    .in(cond_wire70_in),
    .out(cond_wire70_out)
);
std_reg # (
    .WIDTH(1)
) cond71 (
    .clk(cond71_clk),
    .done(cond71_done),
    .in(cond71_in),
    .out(cond71_out),
    .reset(cond71_reset),
    .write_en(cond71_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire71 (
    .in(cond_wire71_in),
    .out(cond_wire71_out)
);
std_reg # (
    .WIDTH(1)
) cond72 (
    .clk(cond72_clk),
    .done(cond72_done),
    .in(cond72_in),
    .out(cond72_out),
    .reset(cond72_reset),
    .write_en(cond72_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire72 (
    .in(cond_wire72_in),
    .out(cond_wire72_out)
);
std_reg # (
    .WIDTH(1)
) cond73 (
    .clk(cond73_clk),
    .done(cond73_done),
    .in(cond73_in),
    .out(cond73_out),
    .reset(cond73_reset),
    .write_en(cond73_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire73 (
    .in(cond_wire73_in),
    .out(cond_wire73_out)
);
std_reg # (
    .WIDTH(1)
) cond74 (
    .clk(cond74_clk),
    .done(cond74_done),
    .in(cond74_in),
    .out(cond74_out),
    .reset(cond74_reset),
    .write_en(cond74_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire74 (
    .in(cond_wire74_in),
    .out(cond_wire74_out)
);
std_reg # (
    .WIDTH(1)
) cond75 (
    .clk(cond75_clk),
    .done(cond75_done),
    .in(cond75_in),
    .out(cond75_out),
    .reset(cond75_reset),
    .write_en(cond75_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire75 (
    .in(cond_wire75_in),
    .out(cond_wire75_out)
);
std_reg # (
    .WIDTH(1)
) cond76 (
    .clk(cond76_clk),
    .done(cond76_done),
    .in(cond76_in),
    .out(cond76_out),
    .reset(cond76_reset),
    .write_en(cond76_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire76 (
    .in(cond_wire76_in),
    .out(cond_wire76_out)
);
std_reg # (
    .WIDTH(1)
) cond77 (
    .clk(cond77_clk),
    .done(cond77_done),
    .in(cond77_in),
    .out(cond77_out),
    .reset(cond77_reset),
    .write_en(cond77_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire77 (
    .in(cond_wire77_in),
    .out(cond_wire77_out)
);
std_reg # (
    .WIDTH(1)
) cond78 (
    .clk(cond78_clk),
    .done(cond78_done),
    .in(cond78_in),
    .out(cond78_out),
    .reset(cond78_reset),
    .write_en(cond78_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire78 (
    .in(cond_wire78_in),
    .out(cond_wire78_out)
);
std_reg # (
    .WIDTH(1)
) cond79 (
    .clk(cond79_clk),
    .done(cond79_done),
    .in(cond79_in),
    .out(cond79_out),
    .reset(cond79_reset),
    .write_en(cond79_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire79 (
    .in(cond_wire79_in),
    .out(cond_wire79_out)
);
std_reg # (
    .WIDTH(1)
) cond80 (
    .clk(cond80_clk),
    .done(cond80_done),
    .in(cond80_in),
    .out(cond80_out),
    .reset(cond80_reset),
    .write_en(cond80_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire80 (
    .in(cond_wire80_in),
    .out(cond_wire80_out)
);
std_reg # (
    .WIDTH(1)
) cond81 (
    .clk(cond81_clk),
    .done(cond81_done),
    .in(cond81_in),
    .out(cond81_out),
    .reset(cond81_reset),
    .write_en(cond81_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire81 (
    .in(cond_wire81_in),
    .out(cond_wire81_out)
);
std_reg # (
    .WIDTH(1)
) cond82 (
    .clk(cond82_clk),
    .done(cond82_done),
    .in(cond82_in),
    .out(cond82_out),
    .reset(cond82_reset),
    .write_en(cond82_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire82 (
    .in(cond_wire82_in),
    .out(cond_wire82_out)
);
std_reg # (
    .WIDTH(1)
) cond83 (
    .clk(cond83_clk),
    .done(cond83_done),
    .in(cond83_in),
    .out(cond83_out),
    .reset(cond83_reset),
    .write_en(cond83_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire83 (
    .in(cond_wire83_in),
    .out(cond_wire83_out)
);
std_reg # (
    .WIDTH(1)
) cond84 (
    .clk(cond84_clk),
    .done(cond84_done),
    .in(cond84_in),
    .out(cond84_out),
    .reset(cond84_reset),
    .write_en(cond84_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire84 (
    .in(cond_wire84_in),
    .out(cond_wire84_out)
);
std_reg # (
    .WIDTH(1)
) cond85 (
    .clk(cond85_clk),
    .done(cond85_done),
    .in(cond85_in),
    .out(cond85_out),
    .reset(cond85_reset),
    .write_en(cond85_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire85 (
    .in(cond_wire85_in),
    .out(cond_wire85_out)
);
std_reg # (
    .WIDTH(1)
) cond86 (
    .clk(cond86_clk),
    .done(cond86_done),
    .in(cond86_in),
    .out(cond86_out),
    .reset(cond86_reset),
    .write_en(cond86_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire86 (
    .in(cond_wire86_in),
    .out(cond_wire86_out)
);
std_reg # (
    .WIDTH(1)
) cond87 (
    .clk(cond87_clk),
    .done(cond87_done),
    .in(cond87_in),
    .out(cond87_out),
    .reset(cond87_reset),
    .write_en(cond87_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire87 (
    .in(cond_wire87_in),
    .out(cond_wire87_out)
);
std_reg # (
    .WIDTH(1)
) cond88 (
    .clk(cond88_clk),
    .done(cond88_done),
    .in(cond88_in),
    .out(cond88_out),
    .reset(cond88_reset),
    .write_en(cond88_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire88 (
    .in(cond_wire88_in),
    .out(cond_wire88_out)
);
std_reg # (
    .WIDTH(1)
) cond89 (
    .clk(cond89_clk),
    .done(cond89_done),
    .in(cond89_in),
    .out(cond89_out),
    .reset(cond89_reset),
    .write_en(cond89_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire89 (
    .in(cond_wire89_in),
    .out(cond_wire89_out)
);
std_reg # (
    .WIDTH(1)
) cond90 (
    .clk(cond90_clk),
    .done(cond90_done),
    .in(cond90_in),
    .out(cond90_out),
    .reset(cond90_reset),
    .write_en(cond90_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire90 (
    .in(cond_wire90_in),
    .out(cond_wire90_out)
);
std_reg # (
    .WIDTH(1)
) cond91 (
    .clk(cond91_clk),
    .done(cond91_done),
    .in(cond91_in),
    .out(cond91_out),
    .reset(cond91_reset),
    .write_en(cond91_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire91 (
    .in(cond_wire91_in),
    .out(cond_wire91_out)
);
std_reg # (
    .WIDTH(1)
) cond92 (
    .clk(cond92_clk),
    .done(cond92_done),
    .in(cond92_in),
    .out(cond92_out),
    .reset(cond92_reset),
    .write_en(cond92_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire92 (
    .in(cond_wire92_in),
    .out(cond_wire92_out)
);
std_reg # (
    .WIDTH(1)
) cond93 (
    .clk(cond93_clk),
    .done(cond93_done),
    .in(cond93_in),
    .out(cond93_out),
    .reset(cond93_reset),
    .write_en(cond93_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire93 (
    .in(cond_wire93_in),
    .out(cond_wire93_out)
);
std_reg # (
    .WIDTH(1)
) cond94 (
    .clk(cond94_clk),
    .done(cond94_done),
    .in(cond94_in),
    .out(cond94_out),
    .reset(cond94_reset),
    .write_en(cond94_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire94 (
    .in(cond_wire94_in),
    .out(cond_wire94_out)
);
std_reg # (
    .WIDTH(1)
) cond95 (
    .clk(cond95_clk),
    .done(cond95_done),
    .in(cond95_in),
    .out(cond95_out),
    .reset(cond95_reset),
    .write_en(cond95_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire95 (
    .in(cond_wire95_in),
    .out(cond_wire95_out)
);
std_reg # (
    .WIDTH(1)
) cond96 (
    .clk(cond96_clk),
    .done(cond96_done),
    .in(cond96_in),
    .out(cond96_out),
    .reset(cond96_reset),
    .write_en(cond96_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire96 (
    .in(cond_wire96_in),
    .out(cond_wire96_out)
);
std_reg # (
    .WIDTH(1)
) cond97 (
    .clk(cond97_clk),
    .done(cond97_done),
    .in(cond97_in),
    .out(cond97_out),
    .reset(cond97_reset),
    .write_en(cond97_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire97 (
    .in(cond_wire97_in),
    .out(cond_wire97_out)
);
std_reg # (
    .WIDTH(1)
) cond98 (
    .clk(cond98_clk),
    .done(cond98_done),
    .in(cond98_in),
    .out(cond98_out),
    .reset(cond98_reset),
    .write_en(cond98_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire98 (
    .in(cond_wire98_in),
    .out(cond_wire98_out)
);
std_reg # (
    .WIDTH(1)
) cond99 (
    .clk(cond99_clk),
    .done(cond99_done),
    .in(cond99_in),
    .out(cond99_out),
    .reset(cond99_reset),
    .write_en(cond99_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire99 (
    .in(cond_wire99_in),
    .out(cond_wire99_out)
);
std_reg # (
    .WIDTH(1)
) cond100 (
    .clk(cond100_clk),
    .done(cond100_done),
    .in(cond100_in),
    .out(cond100_out),
    .reset(cond100_reset),
    .write_en(cond100_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire100 (
    .in(cond_wire100_in),
    .out(cond_wire100_out)
);
std_reg # (
    .WIDTH(1)
) cond101 (
    .clk(cond101_clk),
    .done(cond101_done),
    .in(cond101_in),
    .out(cond101_out),
    .reset(cond101_reset),
    .write_en(cond101_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire101 (
    .in(cond_wire101_in),
    .out(cond_wire101_out)
);
std_reg # (
    .WIDTH(1)
) cond102 (
    .clk(cond102_clk),
    .done(cond102_done),
    .in(cond102_in),
    .out(cond102_out),
    .reset(cond102_reset),
    .write_en(cond102_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire102 (
    .in(cond_wire102_in),
    .out(cond_wire102_out)
);
std_reg # (
    .WIDTH(1)
) cond103 (
    .clk(cond103_clk),
    .done(cond103_done),
    .in(cond103_in),
    .out(cond103_out),
    .reset(cond103_reset),
    .write_en(cond103_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire103 (
    .in(cond_wire103_in),
    .out(cond_wire103_out)
);
std_reg # (
    .WIDTH(1)
) cond104 (
    .clk(cond104_clk),
    .done(cond104_done),
    .in(cond104_in),
    .out(cond104_out),
    .reset(cond104_reset),
    .write_en(cond104_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire104 (
    .in(cond_wire104_in),
    .out(cond_wire104_out)
);
std_reg # (
    .WIDTH(1)
) cond105 (
    .clk(cond105_clk),
    .done(cond105_done),
    .in(cond105_in),
    .out(cond105_out),
    .reset(cond105_reset),
    .write_en(cond105_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire105 (
    .in(cond_wire105_in),
    .out(cond_wire105_out)
);
std_reg # (
    .WIDTH(1)
) cond106 (
    .clk(cond106_clk),
    .done(cond106_done),
    .in(cond106_in),
    .out(cond106_out),
    .reset(cond106_reset),
    .write_en(cond106_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire106 (
    .in(cond_wire106_in),
    .out(cond_wire106_out)
);
std_reg # (
    .WIDTH(1)
) cond107 (
    .clk(cond107_clk),
    .done(cond107_done),
    .in(cond107_in),
    .out(cond107_out),
    .reset(cond107_reset),
    .write_en(cond107_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire107 (
    .in(cond_wire107_in),
    .out(cond_wire107_out)
);
std_reg # (
    .WIDTH(1)
) cond108 (
    .clk(cond108_clk),
    .done(cond108_done),
    .in(cond108_in),
    .out(cond108_out),
    .reset(cond108_reset),
    .write_en(cond108_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire108 (
    .in(cond_wire108_in),
    .out(cond_wire108_out)
);
std_reg # (
    .WIDTH(1)
) cond109 (
    .clk(cond109_clk),
    .done(cond109_done),
    .in(cond109_in),
    .out(cond109_out),
    .reset(cond109_reset),
    .write_en(cond109_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire109 (
    .in(cond_wire109_in),
    .out(cond_wire109_out)
);
std_reg # (
    .WIDTH(1)
) cond110 (
    .clk(cond110_clk),
    .done(cond110_done),
    .in(cond110_in),
    .out(cond110_out),
    .reset(cond110_reset),
    .write_en(cond110_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire110 (
    .in(cond_wire110_in),
    .out(cond_wire110_out)
);
std_reg # (
    .WIDTH(1)
) cond111 (
    .clk(cond111_clk),
    .done(cond111_done),
    .in(cond111_in),
    .out(cond111_out),
    .reset(cond111_reset),
    .write_en(cond111_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire111 (
    .in(cond_wire111_in),
    .out(cond_wire111_out)
);
std_reg # (
    .WIDTH(1)
) cond112 (
    .clk(cond112_clk),
    .done(cond112_done),
    .in(cond112_in),
    .out(cond112_out),
    .reset(cond112_reset),
    .write_en(cond112_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire112 (
    .in(cond_wire112_in),
    .out(cond_wire112_out)
);
std_reg # (
    .WIDTH(1)
) cond113 (
    .clk(cond113_clk),
    .done(cond113_done),
    .in(cond113_in),
    .out(cond113_out),
    .reset(cond113_reset),
    .write_en(cond113_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire113 (
    .in(cond_wire113_in),
    .out(cond_wire113_out)
);
std_reg # (
    .WIDTH(1)
) cond114 (
    .clk(cond114_clk),
    .done(cond114_done),
    .in(cond114_in),
    .out(cond114_out),
    .reset(cond114_reset),
    .write_en(cond114_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire114 (
    .in(cond_wire114_in),
    .out(cond_wire114_out)
);
std_reg # (
    .WIDTH(1)
) cond115 (
    .clk(cond115_clk),
    .done(cond115_done),
    .in(cond115_in),
    .out(cond115_out),
    .reset(cond115_reset),
    .write_en(cond115_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire115 (
    .in(cond_wire115_in),
    .out(cond_wire115_out)
);
std_reg # (
    .WIDTH(1)
) cond116 (
    .clk(cond116_clk),
    .done(cond116_done),
    .in(cond116_in),
    .out(cond116_out),
    .reset(cond116_reset),
    .write_en(cond116_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire116 (
    .in(cond_wire116_in),
    .out(cond_wire116_out)
);
std_reg # (
    .WIDTH(1)
) cond117 (
    .clk(cond117_clk),
    .done(cond117_done),
    .in(cond117_in),
    .out(cond117_out),
    .reset(cond117_reset),
    .write_en(cond117_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire117 (
    .in(cond_wire117_in),
    .out(cond_wire117_out)
);
std_reg # (
    .WIDTH(1)
) cond118 (
    .clk(cond118_clk),
    .done(cond118_done),
    .in(cond118_in),
    .out(cond118_out),
    .reset(cond118_reset),
    .write_en(cond118_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire118 (
    .in(cond_wire118_in),
    .out(cond_wire118_out)
);
std_reg # (
    .WIDTH(1)
) cond119 (
    .clk(cond119_clk),
    .done(cond119_done),
    .in(cond119_in),
    .out(cond119_out),
    .reset(cond119_reset),
    .write_en(cond119_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire119 (
    .in(cond_wire119_in),
    .out(cond_wire119_out)
);
std_reg # (
    .WIDTH(1)
) cond120 (
    .clk(cond120_clk),
    .done(cond120_done),
    .in(cond120_in),
    .out(cond120_out),
    .reset(cond120_reset),
    .write_en(cond120_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire120 (
    .in(cond_wire120_in),
    .out(cond_wire120_out)
);
std_reg # (
    .WIDTH(1)
) cond121 (
    .clk(cond121_clk),
    .done(cond121_done),
    .in(cond121_in),
    .out(cond121_out),
    .reset(cond121_reset),
    .write_en(cond121_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire121 (
    .in(cond_wire121_in),
    .out(cond_wire121_out)
);
std_reg # (
    .WIDTH(1)
) cond122 (
    .clk(cond122_clk),
    .done(cond122_done),
    .in(cond122_in),
    .out(cond122_out),
    .reset(cond122_reset),
    .write_en(cond122_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire122 (
    .in(cond_wire122_in),
    .out(cond_wire122_out)
);
std_reg # (
    .WIDTH(1)
) cond123 (
    .clk(cond123_clk),
    .done(cond123_done),
    .in(cond123_in),
    .out(cond123_out),
    .reset(cond123_reset),
    .write_en(cond123_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire123 (
    .in(cond_wire123_in),
    .out(cond_wire123_out)
);
std_reg # (
    .WIDTH(1)
) cond124 (
    .clk(cond124_clk),
    .done(cond124_done),
    .in(cond124_in),
    .out(cond124_out),
    .reset(cond124_reset),
    .write_en(cond124_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire124 (
    .in(cond_wire124_in),
    .out(cond_wire124_out)
);
std_reg # (
    .WIDTH(1)
) cond125 (
    .clk(cond125_clk),
    .done(cond125_done),
    .in(cond125_in),
    .out(cond125_out),
    .reset(cond125_reset),
    .write_en(cond125_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire125 (
    .in(cond_wire125_in),
    .out(cond_wire125_out)
);
std_reg # (
    .WIDTH(1)
) cond126 (
    .clk(cond126_clk),
    .done(cond126_done),
    .in(cond126_in),
    .out(cond126_out),
    .reset(cond126_reset),
    .write_en(cond126_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire126 (
    .in(cond_wire126_in),
    .out(cond_wire126_out)
);
std_reg # (
    .WIDTH(1)
) cond127 (
    .clk(cond127_clk),
    .done(cond127_done),
    .in(cond127_in),
    .out(cond127_out),
    .reset(cond127_reset),
    .write_en(cond127_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire127 (
    .in(cond_wire127_in),
    .out(cond_wire127_out)
);
std_reg # (
    .WIDTH(1)
) cond128 (
    .clk(cond128_clk),
    .done(cond128_done),
    .in(cond128_in),
    .out(cond128_out),
    .reset(cond128_reset),
    .write_en(cond128_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire128 (
    .in(cond_wire128_in),
    .out(cond_wire128_out)
);
std_reg # (
    .WIDTH(1)
) cond129 (
    .clk(cond129_clk),
    .done(cond129_done),
    .in(cond129_in),
    .out(cond129_out),
    .reset(cond129_reset),
    .write_en(cond129_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire129 (
    .in(cond_wire129_in),
    .out(cond_wire129_out)
);
std_reg # (
    .WIDTH(1)
) cond130 (
    .clk(cond130_clk),
    .done(cond130_done),
    .in(cond130_in),
    .out(cond130_out),
    .reset(cond130_reset),
    .write_en(cond130_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire130 (
    .in(cond_wire130_in),
    .out(cond_wire130_out)
);
std_reg # (
    .WIDTH(1)
) cond131 (
    .clk(cond131_clk),
    .done(cond131_done),
    .in(cond131_in),
    .out(cond131_out),
    .reset(cond131_reset),
    .write_en(cond131_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire131 (
    .in(cond_wire131_in),
    .out(cond_wire131_out)
);
std_reg # (
    .WIDTH(1)
) cond132 (
    .clk(cond132_clk),
    .done(cond132_done),
    .in(cond132_in),
    .out(cond132_out),
    .reset(cond132_reset),
    .write_en(cond132_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire132 (
    .in(cond_wire132_in),
    .out(cond_wire132_out)
);
std_reg # (
    .WIDTH(1)
) cond133 (
    .clk(cond133_clk),
    .done(cond133_done),
    .in(cond133_in),
    .out(cond133_out),
    .reset(cond133_reset),
    .write_en(cond133_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire133 (
    .in(cond_wire133_in),
    .out(cond_wire133_out)
);
std_reg # (
    .WIDTH(1)
) cond134 (
    .clk(cond134_clk),
    .done(cond134_done),
    .in(cond134_in),
    .out(cond134_out),
    .reset(cond134_reset),
    .write_en(cond134_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire134 (
    .in(cond_wire134_in),
    .out(cond_wire134_out)
);
std_reg # (
    .WIDTH(1)
) cond135 (
    .clk(cond135_clk),
    .done(cond135_done),
    .in(cond135_in),
    .out(cond135_out),
    .reset(cond135_reset),
    .write_en(cond135_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire135 (
    .in(cond_wire135_in),
    .out(cond_wire135_out)
);
std_reg # (
    .WIDTH(1)
) cond136 (
    .clk(cond136_clk),
    .done(cond136_done),
    .in(cond136_in),
    .out(cond136_out),
    .reset(cond136_reset),
    .write_en(cond136_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire136 (
    .in(cond_wire136_in),
    .out(cond_wire136_out)
);
std_reg # (
    .WIDTH(1)
) cond137 (
    .clk(cond137_clk),
    .done(cond137_done),
    .in(cond137_in),
    .out(cond137_out),
    .reset(cond137_reset),
    .write_en(cond137_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire137 (
    .in(cond_wire137_in),
    .out(cond_wire137_out)
);
std_reg # (
    .WIDTH(1)
) cond138 (
    .clk(cond138_clk),
    .done(cond138_done),
    .in(cond138_in),
    .out(cond138_out),
    .reset(cond138_reset),
    .write_en(cond138_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire138 (
    .in(cond_wire138_in),
    .out(cond_wire138_out)
);
std_reg # (
    .WIDTH(1)
) cond139 (
    .clk(cond139_clk),
    .done(cond139_done),
    .in(cond139_in),
    .out(cond139_out),
    .reset(cond139_reset),
    .write_en(cond139_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire139 (
    .in(cond_wire139_in),
    .out(cond_wire139_out)
);
std_reg # (
    .WIDTH(1)
) cond140 (
    .clk(cond140_clk),
    .done(cond140_done),
    .in(cond140_in),
    .out(cond140_out),
    .reset(cond140_reset),
    .write_en(cond140_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire140 (
    .in(cond_wire140_in),
    .out(cond_wire140_out)
);
std_reg # (
    .WIDTH(1)
) cond141 (
    .clk(cond141_clk),
    .done(cond141_done),
    .in(cond141_in),
    .out(cond141_out),
    .reset(cond141_reset),
    .write_en(cond141_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire141 (
    .in(cond_wire141_in),
    .out(cond_wire141_out)
);
std_reg # (
    .WIDTH(1)
) cond142 (
    .clk(cond142_clk),
    .done(cond142_done),
    .in(cond142_in),
    .out(cond142_out),
    .reset(cond142_reset),
    .write_en(cond142_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire142 (
    .in(cond_wire142_in),
    .out(cond_wire142_out)
);
std_reg # (
    .WIDTH(1)
) cond143 (
    .clk(cond143_clk),
    .done(cond143_done),
    .in(cond143_in),
    .out(cond143_out),
    .reset(cond143_reset),
    .write_en(cond143_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire143 (
    .in(cond_wire143_in),
    .out(cond_wire143_out)
);
std_reg # (
    .WIDTH(1)
) cond144 (
    .clk(cond144_clk),
    .done(cond144_done),
    .in(cond144_in),
    .out(cond144_out),
    .reset(cond144_reset),
    .write_en(cond144_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire144 (
    .in(cond_wire144_in),
    .out(cond_wire144_out)
);
std_reg # (
    .WIDTH(1)
) cond145 (
    .clk(cond145_clk),
    .done(cond145_done),
    .in(cond145_in),
    .out(cond145_out),
    .reset(cond145_reset),
    .write_en(cond145_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire145 (
    .in(cond_wire145_in),
    .out(cond_wire145_out)
);
std_reg # (
    .WIDTH(1)
) cond146 (
    .clk(cond146_clk),
    .done(cond146_done),
    .in(cond146_in),
    .out(cond146_out),
    .reset(cond146_reset),
    .write_en(cond146_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire146 (
    .in(cond_wire146_in),
    .out(cond_wire146_out)
);
std_reg # (
    .WIDTH(1)
) cond147 (
    .clk(cond147_clk),
    .done(cond147_done),
    .in(cond147_in),
    .out(cond147_out),
    .reset(cond147_reset),
    .write_en(cond147_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire147 (
    .in(cond_wire147_in),
    .out(cond_wire147_out)
);
std_reg # (
    .WIDTH(1)
) cond148 (
    .clk(cond148_clk),
    .done(cond148_done),
    .in(cond148_in),
    .out(cond148_out),
    .reset(cond148_reset),
    .write_en(cond148_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire148 (
    .in(cond_wire148_in),
    .out(cond_wire148_out)
);
std_reg # (
    .WIDTH(1)
) cond149 (
    .clk(cond149_clk),
    .done(cond149_done),
    .in(cond149_in),
    .out(cond149_out),
    .reset(cond149_reset),
    .write_en(cond149_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire149 (
    .in(cond_wire149_in),
    .out(cond_wire149_out)
);
std_reg # (
    .WIDTH(1)
) cond150 (
    .clk(cond150_clk),
    .done(cond150_done),
    .in(cond150_in),
    .out(cond150_out),
    .reset(cond150_reset),
    .write_en(cond150_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire150 (
    .in(cond_wire150_in),
    .out(cond_wire150_out)
);
std_reg # (
    .WIDTH(1)
) cond151 (
    .clk(cond151_clk),
    .done(cond151_done),
    .in(cond151_in),
    .out(cond151_out),
    .reset(cond151_reset),
    .write_en(cond151_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire151 (
    .in(cond_wire151_in),
    .out(cond_wire151_out)
);
std_reg # (
    .WIDTH(1)
) cond152 (
    .clk(cond152_clk),
    .done(cond152_done),
    .in(cond152_in),
    .out(cond152_out),
    .reset(cond152_reset),
    .write_en(cond152_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire152 (
    .in(cond_wire152_in),
    .out(cond_wire152_out)
);
std_reg # (
    .WIDTH(1)
) cond153 (
    .clk(cond153_clk),
    .done(cond153_done),
    .in(cond153_in),
    .out(cond153_out),
    .reset(cond153_reset),
    .write_en(cond153_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire153 (
    .in(cond_wire153_in),
    .out(cond_wire153_out)
);
std_reg # (
    .WIDTH(1)
) cond154 (
    .clk(cond154_clk),
    .done(cond154_done),
    .in(cond154_in),
    .out(cond154_out),
    .reset(cond154_reset),
    .write_en(cond154_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire154 (
    .in(cond_wire154_in),
    .out(cond_wire154_out)
);
std_reg # (
    .WIDTH(1)
) cond155 (
    .clk(cond155_clk),
    .done(cond155_done),
    .in(cond155_in),
    .out(cond155_out),
    .reset(cond155_reset),
    .write_en(cond155_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire155 (
    .in(cond_wire155_in),
    .out(cond_wire155_out)
);
std_reg # (
    .WIDTH(1)
) cond156 (
    .clk(cond156_clk),
    .done(cond156_done),
    .in(cond156_in),
    .out(cond156_out),
    .reset(cond156_reset),
    .write_en(cond156_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire156 (
    .in(cond_wire156_in),
    .out(cond_wire156_out)
);
std_reg # (
    .WIDTH(1)
) cond157 (
    .clk(cond157_clk),
    .done(cond157_done),
    .in(cond157_in),
    .out(cond157_out),
    .reset(cond157_reset),
    .write_en(cond157_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire157 (
    .in(cond_wire157_in),
    .out(cond_wire157_out)
);
std_reg # (
    .WIDTH(1)
) cond158 (
    .clk(cond158_clk),
    .done(cond158_done),
    .in(cond158_in),
    .out(cond158_out),
    .reset(cond158_reset),
    .write_en(cond158_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire158 (
    .in(cond_wire158_in),
    .out(cond_wire158_out)
);
std_reg # (
    .WIDTH(1)
) cond159 (
    .clk(cond159_clk),
    .done(cond159_done),
    .in(cond159_in),
    .out(cond159_out),
    .reset(cond159_reset),
    .write_en(cond159_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire159 (
    .in(cond_wire159_in),
    .out(cond_wire159_out)
);
std_reg # (
    .WIDTH(1)
) cond160 (
    .clk(cond160_clk),
    .done(cond160_done),
    .in(cond160_in),
    .out(cond160_out),
    .reset(cond160_reset),
    .write_en(cond160_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire160 (
    .in(cond_wire160_in),
    .out(cond_wire160_out)
);
std_reg # (
    .WIDTH(1)
) cond161 (
    .clk(cond161_clk),
    .done(cond161_done),
    .in(cond161_in),
    .out(cond161_out),
    .reset(cond161_reset),
    .write_en(cond161_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire161 (
    .in(cond_wire161_in),
    .out(cond_wire161_out)
);
std_reg # (
    .WIDTH(1)
) cond162 (
    .clk(cond162_clk),
    .done(cond162_done),
    .in(cond162_in),
    .out(cond162_out),
    .reset(cond162_reset),
    .write_en(cond162_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire162 (
    .in(cond_wire162_in),
    .out(cond_wire162_out)
);
std_reg # (
    .WIDTH(1)
) cond163 (
    .clk(cond163_clk),
    .done(cond163_done),
    .in(cond163_in),
    .out(cond163_out),
    .reset(cond163_reset),
    .write_en(cond163_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire163 (
    .in(cond_wire163_in),
    .out(cond_wire163_out)
);
std_reg # (
    .WIDTH(1)
) cond164 (
    .clk(cond164_clk),
    .done(cond164_done),
    .in(cond164_in),
    .out(cond164_out),
    .reset(cond164_reset),
    .write_en(cond164_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire164 (
    .in(cond_wire164_in),
    .out(cond_wire164_out)
);
std_reg # (
    .WIDTH(1)
) cond165 (
    .clk(cond165_clk),
    .done(cond165_done),
    .in(cond165_in),
    .out(cond165_out),
    .reset(cond165_reset),
    .write_en(cond165_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire165 (
    .in(cond_wire165_in),
    .out(cond_wire165_out)
);
std_reg # (
    .WIDTH(1)
) cond166 (
    .clk(cond166_clk),
    .done(cond166_done),
    .in(cond166_in),
    .out(cond166_out),
    .reset(cond166_reset),
    .write_en(cond166_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire166 (
    .in(cond_wire166_in),
    .out(cond_wire166_out)
);
std_reg # (
    .WIDTH(1)
) cond167 (
    .clk(cond167_clk),
    .done(cond167_done),
    .in(cond167_in),
    .out(cond167_out),
    .reset(cond167_reset),
    .write_en(cond167_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire167 (
    .in(cond_wire167_in),
    .out(cond_wire167_out)
);
std_reg # (
    .WIDTH(1)
) cond168 (
    .clk(cond168_clk),
    .done(cond168_done),
    .in(cond168_in),
    .out(cond168_out),
    .reset(cond168_reset),
    .write_en(cond168_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire168 (
    .in(cond_wire168_in),
    .out(cond_wire168_out)
);
std_reg # (
    .WIDTH(1)
) cond169 (
    .clk(cond169_clk),
    .done(cond169_done),
    .in(cond169_in),
    .out(cond169_out),
    .reset(cond169_reset),
    .write_en(cond169_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire169 (
    .in(cond_wire169_in),
    .out(cond_wire169_out)
);
std_reg # (
    .WIDTH(1)
) cond170 (
    .clk(cond170_clk),
    .done(cond170_done),
    .in(cond170_in),
    .out(cond170_out),
    .reset(cond170_reset),
    .write_en(cond170_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire170 (
    .in(cond_wire170_in),
    .out(cond_wire170_out)
);
std_reg # (
    .WIDTH(1)
) cond171 (
    .clk(cond171_clk),
    .done(cond171_done),
    .in(cond171_in),
    .out(cond171_out),
    .reset(cond171_reset),
    .write_en(cond171_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire171 (
    .in(cond_wire171_in),
    .out(cond_wire171_out)
);
std_reg # (
    .WIDTH(1)
) cond172 (
    .clk(cond172_clk),
    .done(cond172_done),
    .in(cond172_in),
    .out(cond172_out),
    .reset(cond172_reset),
    .write_en(cond172_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire172 (
    .in(cond_wire172_in),
    .out(cond_wire172_out)
);
std_reg # (
    .WIDTH(1)
) cond173 (
    .clk(cond173_clk),
    .done(cond173_done),
    .in(cond173_in),
    .out(cond173_out),
    .reset(cond173_reset),
    .write_en(cond173_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire173 (
    .in(cond_wire173_in),
    .out(cond_wire173_out)
);
std_reg # (
    .WIDTH(1)
) cond174 (
    .clk(cond174_clk),
    .done(cond174_done),
    .in(cond174_in),
    .out(cond174_out),
    .reset(cond174_reset),
    .write_en(cond174_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire174 (
    .in(cond_wire174_in),
    .out(cond_wire174_out)
);
std_reg # (
    .WIDTH(1)
) cond175 (
    .clk(cond175_clk),
    .done(cond175_done),
    .in(cond175_in),
    .out(cond175_out),
    .reset(cond175_reset),
    .write_en(cond175_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire175 (
    .in(cond_wire175_in),
    .out(cond_wire175_out)
);
std_reg # (
    .WIDTH(1)
) cond176 (
    .clk(cond176_clk),
    .done(cond176_done),
    .in(cond176_in),
    .out(cond176_out),
    .reset(cond176_reset),
    .write_en(cond176_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire176 (
    .in(cond_wire176_in),
    .out(cond_wire176_out)
);
std_reg # (
    .WIDTH(1)
) cond177 (
    .clk(cond177_clk),
    .done(cond177_done),
    .in(cond177_in),
    .out(cond177_out),
    .reset(cond177_reset),
    .write_en(cond177_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire177 (
    .in(cond_wire177_in),
    .out(cond_wire177_out)
);
std_reg # (
    .WIDTH(1)
) cond178 (
    .clk(cond178_clk),
    .done(cond178_done),
    .in(cond178_in),
    .out(cond178_out),
    .reset(cond178_reset),
    .write_en(cond178_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire178 (
    .in(cond_wire178_in),
    .out(cond_wire178_out)
);
std_reg # (
    .WIDTH(1)
) cond179 (
    .clk(cond179_clk),
    .done(cond179_done),
    .in(cond179_in),
    .out(cond179_out),
    .reset(cond179_reset),
    .write_en(cond179_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire179 (
    .in(cond_wire179_in),
    .out(cond_wire179_out)
);
std_reg # (
    .WIDTH(1)
) cond180 (
    .clk(cond180_clk),
    .done(cond180_done),
    .in(cond180_in),
    .out(cond180_out),
    .reset(cond180_reset),
    .write_en(cond180_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire180 (
    .in(cond_wire180_in),
    .out(cond_wire180_out)
);
std_reg # (
    .WIDTH(1)
) cond181 (
    .clk(cond181_clk),
    .done(cond181_done),
    .in(cond181_in),
    .out(cond181_out),
    .reset(cond181_reset),
    .write_en(cond181_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire181 (
    .in(cond_wire181_in),
    .out(cond_wire181_out)
);
std_reg # (
    .WIDTH(1)
) cond182 (
    .clk(cond182_clk),
    .done(cond182_done),
    .in(cond182_in),
    .out(cond182_out),
    .reset(cond182_reset),
    .write_en(cond182_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire182 (
    .in(cond_wire182_in),
    .out(cond_wire182_out)
);
std_reg # (
    .WIDTH(1)
) cond183 (
    .clk(cond183_clk),
    .done(cond183_done),
    .in(cond183_in),
    .out(cond183_out),
    .reset(cond183_reset),
    .write_en(cond183_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire183 (
    .in(cond_wire183_in),
    .out(cond_wire183_out)
);
std_reg # (
    .WIDTH(1)
) cond184 (
    .clk(cond184_clk),
    .done(cond184_done),
    .in(cond184_in),
    .out(cond184_out),
    .reset(cond184_reset),
    .write_en(cond184_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire184 (
    .in(cond_wire184_in),
    .out(cond_wire184_out)
);
std_reg # (
    .WIDTH(1)
) cond185 (
    .clk(cond185_clk),
    .done(cond185_done),
    .in(cond185_in),
    .out(cond185_out),
    .reset(cond185_reset),
    .write_en(cond185_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire185 (
    .in(cond_wire185_in),
    .out(cond_wire185_out)
);
std_reg # (
    .WIDTH(1)
) cond186 (
    .clk(cond186_clk),
    .done(cond186_done),
    .in(cond186_in),
    .out(cond186_out),
    .reset(cond186_reset),
    .write_en(cond186_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire186 (
    .in(cond_wire186_in),
    .out(cond_wire186_out)
);
std_reg # (
    .WIDTH(1)
) cond187 (
    .clk(cond187_clk),
    .done(cond187_done),
    .in(cond187_in),
    .out(cond187_out),
    .reset(cond187_reset),
    .write_en(cond187_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire187 (
    .in(cond_wire187_in),
    .out(cond_wire187_out)
);
std_reg # (
    .WIDTH(1)
) cond188 (
    .clk(cond188_clk),
    .done(cond188_done),
    .in(cond188_in),
    .out(cond188_out),
    .reset(cond188_reset),
    .write_en(cond188_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire188 (
    .in(cond_wire188_in),
    .out(cond_wire188_out)
);
std_reg # (
    .WIDTH(1)
) cond189 (
    .clk(cond189_clk),
    .done(cond189_done),
    .in(cond189_in),
    .out(cond189_out),
    .reset(cond189_reset),
    .write_en(cond189_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire189 (
    .in(cond_wire189_in),
    .out(cond_wire189_out)
);
std_reg # (
    .WIDTH(1)
) cond190 (
    .clk(cond190_clk),
    .done(cond190_done),
    .in(cond190_in),
    .out(cond190_out),
    .reset(cond190_reset),
    .write_en(cond190_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire190 (
    .in(cond_wire190_in),
    .out(cond_wire190_out)
);
std_reg # (
    .WIDTH(1)
) cond191 (
    .clk(cond191_clk),
    .done(cond191_done),
    .in(cond191_in),
    .out(cond191_out),
    .reset(cond191_reset),
    .write_en(cond191_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire191 (
    .in(cond_wire191_in),
    .out(cond_wire191_out)
);
std_reg # (
    .WIDTH(1)
) cond192 (
    .clk(cond192_clk),
    .done(cond192_done),
    .in(cond192_in),
    .out(cond192_out),
    .reset(cond192_reset),
    .write_en(cond192_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire192 (
    .in(cond_wire192_in),
    .out(cond_wire192_out)
);
std_reg # (
    .WIDTH(1)
) cond193 (
    .clk(cond193_clk),
    .done(cond193_done),
    .in(cond193_in),
    .out(cond193_out),
    .reset(cond193_reset),
    .write_en(cond193_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire193 (
    .in(cond_wire193_in),
    .out(cond_wire193_out)
);
std_reg # (
    .WIDTH(1)
) cond194 (
    .clk(cond194_clk),
    .done(cond194_done),
    .in(cond194_in),
    .out(cond194_out),
    .reset(cond194_reset),
    .write_en(cond194_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire194 (
    .in(cond_wire194_in),
    .out(cond_wire194_out)
);
std_reg # (
    .WIDTH(1)
) cond195 (
    .clk(cond195_clk),
    .done(cond195_done),
    .in(cond195_in),
    .out(cond195_out),
    .reset(cond195_reset),
    .write_en(cond195_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire195 (
    .in(cond_wire195_in),
    .out(cond_wire195_out)
);
std_reg # (
    .WIDTH(1)
) cond196 (
    .clk(cond196_clk),
    .done(cond196_done),
    .in(cond196_in),
    .out(cond196_out),
    .reset(cond196_reset),
    .write_en(cond196_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire196 (
    .in(cond_wire196_in),
    .out(cond_wire196_out)
);
std_reg # (
    .WIDTH(1)
) cond197 (
    .clk(cond197_clk),
    .done(cond197_done),
    .in(cond197_in),
    .out(cond197_out),
    .reset(cond197_reset),
    .write_en(cond197_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire197 (
    .in(cond_wire197_in),
    .out(cond_wire197_out)
);
std_reg # (
    .WIDTH(1)
) cond198 (
    .clk(cond198_clk),
    .done(cond198_done),
    .in(cond198_in),
    .out(cond198_out),
    .reset(cond198_reset),
    .write_en(cond198_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire198 (
    .in(cond_wire198_in),
    .out(cond_wire198_out)
);
std_reg # (
    .WIDTH(1)
) cond199 (
    .clk(cond199_clk),
    .done(cond199_done),
    .in(cond199_in),
    .out(cond199_out),
    .reset(cond199_reset),
    .write_en(cond199_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire199 (
    .in(cond_wire199_in),
    .out(cond_wire199_out)
);
std_reg # (
    .WIDTH(1)
) cond200 (
    .clk(cond200_clk),
    .done(cond200_done),
    .in(cond200_in),
    .out(cond200_out),
    .reset(cond200_reset),
    .write_en(cond200_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire200 (
    .in(cond_wire200_in),
    .out(cond_wire200_out)
);
std_reg # (
    .WIDTH(1)
) cond201 (
    .clk(cond201_clk),
    .done(cond201_done),
    .in(cond201_in),
    .out(cond201_out),
    .reset(cond201_reset),
    .write_en(cond201_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire201 (
    .in(cond_wire201_in),
    .out(cond_wire201_out)
);
std_reg # (
    .WIDTH(1)
) cond202 (
    .clk(cond202_clk),
    .done(cond202_done),
    .in(cond202_in),
    .out(cond202_out),
    .reset(cond202_reset),
    .write_en(cond202_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire202 (
    .in(cond_wire202_in),
    .out(cond_wire202_out)
);
std_reg # (
    .WIDTH(1)
) cond203 (
    .clk(cond203_clk),
    .done(cond203_done),
    .in(cond203_in),
    .out(cond203_out),
    .reset(cond203_reset),
    .write_en(cond203_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire203 (
    .in(cond_wire203_in),
    .out(cond_wire203_out)
);
std_reg # (
    .WIDTH(1)
) cond204 (
    .clk(cond204_clk),
    .done(cond204_done),
    .in(cond204_in),
    .out(cond204_out),
    .reset(cond204_reset),
    .write_en(cond204_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire204 (
    .in(cond_wire204_in),
    .out(cond_wire204_out)
);
std_reg # (
    .WIDTH(1)
) cond205 (
    .clk(cond205_clk),
    .done(cond205_done),
    .in(cond205_in),
    .out(cond205_out),
    .reset(cond205_reset),
    .write_en(cond205_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire205 (
    .in(cond_wire205_in),
    .out(cond_wire205_out)
);
std_reg # (
    .WIDTH(1)
) cond206 (
    .clk(cond206_clk),
    .done(cond206_done),
    .in(cond206_in),
    .out(cond206_out),
    .reset(cond206_reset),
    .write_en(cond206_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire206 (
    .in(cond_wire206_in),
    .out(cond_wire206_out)
);
std_reg # (
    .WIDTH(1)
) cond207 (
    .clk(cond207_clk),
    .done(cond207_done),
    .in(cond207_in),
    .out(cond207_out),
    .reset(cond207_reset),
    .write_en(cond207_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire207 (
    .in(cond_wire207_in),
    .out(cond_wire207_out)
);
std_reg # (
    .WIDTH(1)
) cond208 (
    .clk(cond208_clk),
    .done(cond208_done),
    .in(cond208_in),
    .out(cond208_out),
    .reset(cond208_reset),
    .write_en(cond208_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire208 (
    .in(cond_wire208_in),
    .out(cond_wire208_out)
);
std_reg # (
    .WIDTH(1)
) cond209 (
    .clk(cond209_clk),
    .done(cond209_done),
    .in(cond209_in),
    .out(cond209_out),
    .reset(cond209_reset),
    .write_en(cond209_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire209 (
    .in(cond_wire209_in),
    .out(cond_wire209_out)
);
std_reg # (
    .WIDTH(1)
) cond210 (
    .clk(cond210_clk),
    .done(cond210_done),
    .in(cond210_in),
    .out(cond210_out),
    .reset(cond210_reset),
    .write_en(cond210_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire210 (
    .in(cond_wire210_in),
    .out(cond_wire210_out)
);
std_reg # (
    .WIDTH(1)
) cond211 (
    .clk(cond211_clk),
    .done(cond211_done),
    .in(cond211_in),
    .out(cond211_out),
    .reset(cond211_reset),
    .write_en(cond211_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire211 (
    .in(cond_wire211_in),
    .out(cond_wire211_out)
);
std_reg # (
    .WIDTH(1)
) cond212 (
    .clk(cond212_clk),
    .done(cond212_done),
    .in(cond212_in),
    .out(cond212_out),
    .reset(cond212_reset),
    .write_en(cond212_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire212 (
    .in(cond_wire212_in),
    .out(cond_wire212_out)
);
std_reg # (
    .WIDTH(1)
) cond213 (
    .clk(cond213_clk),
    .done(cond213_done),
    .in(cond213_in),
    .out(cond213_out),
    .reset(cond213_reset),
    .write_en(cond213_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire213 (
    .in(cond_wire213_in),
    .out(cond_wire213_out)
);
std_reg # (
    .WIDTH(1)
) cond214 (
    .clk(cond214_clk),
    .done(cond214_done),
    .in(cond214_in),
    .out(cond214_out),
    .reset(cond214_reset),
    .write_en(cond214_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire214 (
    .in(cond_wire214_in),
    .out(cond_wire214_out)
);
std_reg # (
    .WIDTH(1)
) cond215 (
    .clk(cond215_clk),
    .done(cond215_done),
    .in(cond215_in),
    .out(cond215_out),
    .reset(cond215_reset),
    .write_en(cond215_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire215 (
    .in(cond_wire215_in),
    .out(cond_wire215_out)
);
std_reg # (
    .WIDTH(1)
) cond216 (
    .clk(cond216_clk),
    .done(cond216_done),
    .in(cond216_in),
    .out(cond216_out),
    .reset(cond216_reset),
    .write_en(cond216_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire216 (
    .in(cond_wire216_in),
    .out(cond_wire216_out)
);
std_reg # (
    .WIDTH(1)
) cond217 (
    .clk(cond217_clk),
    .done(cond217_done),
    .in(cond217_in),
    .out(cond217_out),
    .reset(cond217_reset),
    .write_en(cond217_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire217 (
    .in(cond_wire217_in),
    .out(cond_wire217_out)
);
std_reg # (
    .WIDTH(1)
) cond218 (
    .clk(cond218_clk),
    .done(cond218_done),
    .in(cond218_in),
    .out(cond218_out),
    .reset(cond218_reset),
    .write_en(cond218_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire218 (
    .in(cond_wire218_in),
    .out(cond_wire218_out)
);
std_reg # (
    .WIDTH(1)
) cond219 (
    .clk(cond219_clk),
    .done(cond219_done),
    .in(cond219_in),
    .out(cond219_out),
    .reset(cond219_reset),
    .write_en(cond219_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire219 (
    .in(cond_wire219_in),
    .out(cond_wire219_out)
);
std_reg # (
    .WIDTH(1)
) cond220 (
    .clk(cond220_clk),
    .done(cond220_done),
    .in(cond220_in),
    .out(cond220_out),
    .reset(cond220_reset),
    .write_en(cond220_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire220 (
    .in(cond_wire220_in),
    .out(cond_wire220_out)
);
std_reg # (
    .WIDTH(1)
) cond221 (
    .clk(cond221_clk),
    .done(cond221_done),
    .in(cond221_in),
    .out(cond221_out),
    .reset(cond221_reset),
    .write_en(cond221_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire221 (
    .in(cond_wire221_in),
    .out(cond_wire221_out)
);
std_reg # (
    .WIDTH(1)
) cond222 (
    .clk(cond222_clk),
    .done(cond222_done),
    .in(cond222_in),
    .out(cond222_out),
    .reset(cond222_reset),
    .write_en(cond222_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire222 (
    .in(cond_wire222_in),
    .out(cond_wire222_out)
);
std_reg # (
    .WIDTH(1)
) cond223 (
    .clk(cond223_clk),
    .done(cond223_done),
    .in(cond223_in),
    .out(cond223_out),
    .reset(cond223_reset),
    .write_en(cond223_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire223 (
    .in(cond_wire223_in),
    .out(cond_wire223_out)
);
std_reg # (
    .WIDTH(1)
) cond224 (
    .clk(cond224_clk),
    .done(cond224_done),
    .in(cond224_in),
    .out(cond224_out),
    .reset(cond224_reset),
    .write_en(cond224_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire224 (
    .in(cond_wire224_in),
    .out(cond_wire224_out)
);
std_reg # (
    .WIDTH(1)
) cond225 (
    .clk(cond225_clk),
    .done(cond225_done),
    .in(cond225_in),
    .out(cond225_out),
    .reset(cond225_reset),
    .write_en(cond225_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire225 (
    .in(cond_wire225_in),
    .out(cond_wire225_out)
);
std_reg # (
    .WIDTH(1)
) cond226 (
    .clk(cond226_clk),
    .done(cond226_done),
    .in(cond226_in),
    .out(cond226_out),
    .reset(cond226_reset),
    .write_en(cond226_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire226 (
    .in(cond_wire226_in),
    .out(cond_wire226_out)
);
std_reg # (
    .WIDTH(1)
) cond227 (
    .clk(cond227_clk),
    .done(cond227_done),
    .in(cond227_in),
    .out(cond227_out),
    .reset(cond227_reset),
    .write_en(cond227_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire227 (
    .in(cond_wire227_in),
    .out(cond_wire227_out)
);
std_reg # (
    .WIDTH(1)
) cond228 (
    .clk(cond228_clk),
    .done(cond228_done),
    .in(cond228_in),
    .out(cond228_out),
    .reset(cond228_reset),
    .write_en(cond228_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire228 (
    .in(cond_wire228_in),
    .out(cond_wire228_out)
);
std_reg # (
    .WIDTH(1)
) cond229 (
    .clk(cond229_clk),
    .done(cond229_done),
    .in(cond229_in),
    .out(cond229_out),
    .reset(cond229_reset),
    .write_en(cond229_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire229 (
    .in(cond_wire229_in),
    .out(cond_wire229_out)
);
std_reg # (
    .WIDTH(1)
) cond230 (
    .clk(cond230_clk),
    .done(cond230_done),
    .in(cond230_in),
    .out(cond230_out),
    .reset(cond230_reset),
    .write_en(cond230_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire230 (
    .in(cond_wire230_in),
    .out(cond_wire230_out)
);
std_reg # (
    .WIDTH(1)
) cond231 (
    .clk(cond231_clk),
    .done(cond231_done),
    .in(cond231_in),
    .out(cond231_out),
    .reset(cond231_reset),
    .write_en(cond231_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire231 (
    .in(cond_wire231_in),
    .out(cond_wire231_out)
);
std_reg # (
    .WIDTH(1)
) cond232 (
    .clk(cond232_clk),
    .done(cond232_done),
    .in(cond232_in),
    .out(cond232_out),
    .reset(cond232_reset),
    .write_en(cond232_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire232 (
    .in(cond_wire232_in),
    .out(cond_wire232_out)
);
std_reg # (
    .WIDTH(1)
) cond233 (
    .clk(cond233_clk),
    .done(cond233_done),
    .in(cond233_in),
    .out(cond233_out),
    .reset(cond233_reset),
    .write_en(cond233_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire233 (
    .in(cond_wire233_in),
    .out(cond_wire233_out)
);
std_reg # (
    .WIDTH(1)
) cond234 (
    .clk(cond234_clk),
    .done(cond234_done),
    .in(cond234_in),
    .out(cond234_out),
    .reset(cond234_reset),
    .write_en(cond234_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire234 (
    .in(cond_wire234_in),
    .out(cond_wire234_out)
);
std_reg # (
    .WIDTH(1)
) cond235 (
    .clk(cond235_clk),
    .done(cond235_done),
    .in(cond235_in),
    .out(cond235_out),
    .reset(cond235_reset),
    .write_en(cond235_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire235 (
    .in(cond_wire235_in),
    .out(cond_wire235_out)
);
std_reg # (
    .WIDTH(1)
) cond236 (
    .clk(cond236_clk),
    .done(cond236_done),
    .in(cond236_in),
    .out(cond236_out),
    .reset(cond236_reset),
    .write_en(cond236_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire236 (
    .in(cond_wire236_in),
    .out(cond_wire236_out)
);
std_reg # (
    .WIDTH(1)
) cond237 (
    .clk(cond237_clk),
    .done(cond237_done),
    .in(cond237_in),
    .out(cond237_out),
    .reset(cond237_reset),
    .write_en(cond237_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire237 (
    .in(cond_wire237_in),
    .out(cond_wire237_out)
);
std_reg # (
    .WIDTH(1)
) cond238 (
    .clk(cond238_clk),
    .done(cond238_done),
    .in(cond238_in),
    .out(cond238_out),
    .reset(cond238_reset),
    .write_en(cond238_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire238 (
    .in(cond_wire238_in),
    .out(cond_wire238_out)
);
std_reg # (
    .WIDTH(1)
) cond239 (
    .clk(cond239_clk),
    .done(cond239_done),
    .in(cond239_in),
    .out(cond239_out),
    .reset(cond239_reset),
    .write_en(cond239_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire239 (
    .in(cond_wire239_in),
    .out(cond_wire239_out)
);
std_reg # (
    .WIDTH(1)
) cond240 (
    .clk(cond240_clk),
    .done(cond240_done),
    .in(cond240_in),
    .out(cond240_out),
    .reset(cond240_reset),
    .write_en(cond240_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire240 (
    .in(cond_wire240_in),
    .out(cond_wire240_out)
);
std_reg # (
    .WIDTH(1)
) cond241 (
    .clk(cond241_clk),
    .done(cond241_done),
    .in(cond241_in),
    .out(cond241_out),
    .reset(cond241_reset),
    .write_en(cond241_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire241 (
    .in(cond_wire241_in),
    .out(cond_wire241_out)
);
std_reg # (
    .WIDTH(1)
) cond242 (
    .clk(cond242_clk),
    .done(cond242_done),
    .in(cond242_in),
    .out(cond242_out),
    .reset(cond242_reset),
    .write_en(cond242_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire242 (
    .in(cond_wire242_in),
    .out(cond_wire242_out)
);
std_reg # (
    .WIDTH(1)
) cond243 (
    .clk(cond243_clk),
    .done(cond243_done),
    .in(cond243_in),
    .out(cond243_out),
    .reset(cond243_reset),
    .write_en(cond243_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire243 (
    .in(cond_wire243_in),
    .out(cond_wire243_out)
);
std_reg # (
    .WIDTH(1)
) cond244 (
    .clk(cond244_clk),
    .done(cond244_done),
    .in(cond244_in),
    .out(cond244_out),
    .reset(cond244_reset),
    .write_en(cond244_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire244 (
    .in(cond_wire244_in),
    .out(cond_wire244_out)
);
std_reg # (
    .WIDTH(1)
) cond245 (
    .clk(cond245_clk),
    .done(cond245_done),
    .in(cond245_in),
    .out(cond245_out),
    .reset(cond245_reset),
    .write_en(cond245_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire245 (
    .in(cond_wire245_in),
    .out(cond_wire245_out)
);
std_reg # (
    .WIDTH(1)
) cond246 (
    .clk(cond246_clk),
    .done(cond246_done),
    .in(cond246_in),
    .out(cond246_out),
    .reset(cond246_reset),
    .write_en(cond246_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire246 (
    .in(cond_wire246_in),
    .out(cond_wire246_out)
);
std_reg # (
    .WIDTH(1)
) cond247 (
    .clk(cond247_clk),
    .done(cond247_done),
    .in(cond247_in),
    .out(cond247_out),
    .reset(cond247_reset),
    .write_en(cond247_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire247 (
    .in(cond_wire247_in),
    .out(cond_wire247_out)
);
std_reg # (
    .WIDTH(1)
) cond248 (
    .clk(cond248_clk),
    .done(cond248_done),
    .in(cond248_in),
    .out(cond248_out),
    .reset(cond248_reset),
    .write_en(cond248_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire248 (
    .in(cond_wire248_in),
    .out(cond_wire248_out)
);
std_reg # (
    .WIDTH(1)
) cond249 (
    .clk(cond249_clk),
    .done(cond249_done),
    .in(cond249_in),
    .out(cond249_out),
    .reset(cond249_reset),
    .write_en(cond249_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire249 (
    .in(cond_wire249_in),
    .out(cond_wire249_out)
);
std_reg # (
    .WIDTH(1)
) cond250 (
    .clk(cond250_clk),
    .done(cond250_done),
    .in(cond250_in),
    .out(cond250_out),
    .reset(cond250_reset),
    .write_en(cond250_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire250 (
    .in(cond_wire250_in),
    .out(cond_wire250_out)
);
std_reg # (
    .WIDTH(1)
) cond251 (
    .clk(cond251_clk),
    .done(cond251_done),
    .in(cond251_in),
    .out(cond251_out),
    .reset(cond251_reset),
    .write_en(cond251_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire251 (
    .in(cond_wire251_in),
    .out(cond_wire251_out)
);
std_reg # (
    .WIDTH(1)
) cond252 (
    .clk(cond252_clk),
    .done(cond252_done),
    .in(cond252_in),
    .out(cond252_out),
    .reset(cond252_reset),
    .write_en(cond252_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire252 (
    .in(cond_wire252_in),
    .out(cond_wire252_out)
);
std_reg # (
    .WIDTH(1)
) cond253 (
    .clk(cond253_clk),
    .done(cond253_done),
    .in(cond253_in),
    .out(cond253_out),
    .reset(cond253_reset),
    .write_en(cond253_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire253 (
    .in(cond_wire253_in),
    .out(cond_wire253_out)
);
std_reg # (
    .WIDTH(1)
) cond254 (
    .clk(cond254_clk),
    .done(cond254_done),
    .in(cond254_in),
    .out(cond254_out),
    .reset(cond254_reset),
    .write_en(cond254_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire254 (
    .in(cond_wire254_in),
    .out(cond_wire254_out)
);
std_reg # (
    .WIDTH(1)
) cond255 (
    .clk(cond255_clk),
    .done(cond255_done),
    .in(cond255_in),
    .out(cond255_out),
    .reset(cond255_reset),
    .write_en(cond255_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire255 (
    .in(cond_wire255_in),
    .out(cond_wire255_out)
);
std_reg # (
    .WIDTH(1)
) cond256 (
    .clk(cond256_clk),
    .done(cond256_done),
    .in(cond256_in),
    .out(cond256_out),
    .reset(cond256_reset),
    .write_en(cond256_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire256 (
    .in(cond_wire256_in),
    .out(cond_wire256_out)
);
std_reg # (
    .WIDTH(1)
) cond257 (
    .clk(cond257_clk),
    .done(cond257_done),
    .in(cond257_in),
    .out(cond257_out),
    .reset(cond257_reset),
    .write_en(cond257_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire257 (
    .in(cond_wire257_in),
    .out(cond_wire257_out)
);
std_reg # (
    .WIDTH(1)
) cond258 (
    .clk(cond258_clk),
    .done(cond258_done),
    .in(cond258_in),
    .out(cond258_out),
    .reset(cond258_reset),
    .write_en(cond258_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire258 (
    .in(cond_wire258_in),
    .out(cond_wire258_out)
);
std_reg # (
    .WIDTH(1)
) cond259 (
    .clk(cond259_clk),
    .done(cond259_done),
    .in(cond259_in),
    .out(cond259_out),
    .reset(cond259_reset),
    .write_en(cond259_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire259 (
    .in(cond_wire259_in),
    .out(cond_wire259_out)
);
std_reg # (
    .WIDTH(1)
) cond260 (
    .clk(cond260_clk),
    .done(cond260_done),
    .in(cond260_in),
    .out(cond260_out),
    .reset(cond260_reset),
    .write_en(cond260_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire260 (
    .in(cond_wire260_in),
    .out(cond_wire260_out)
);
std_reg # (
    .WIDTH(1)
) cond261 (
    .clk(cond261_clk),
    .done(cond261_done),
    .in(cond261_in),
    .out(cond261_out),
    .reset(cond261_reset),
    .write_en(cond261_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire261 (
    .in(cond_wire261_in),
    .out(cond_wire261_out)
);
std_reg # (
    .WIDTH(1)
) cond262 (
    .clk(cond262_clk),
    .done(cond262_done),
    .in(cond262_in),
    .out(cond262_out),
    .reset(cond262_reset),
    .write_en(cond262_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire262 (
    .in(cond_wire262_in),
    .out(cond_wire262_out)
);
std_reg # (
    .WIDTH(1)
) cond263 (
    .clk(cond263_clk),
    .done(cond263_done),
    .in(cond263_in),
    .out(cond263_out),
    .reset(cond263_reset),
    .write_en(cond263_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire263 (
    .in(cond_wire263_in),
    .out(cond_wire263_out)
);
std_reg # (
    .WIDTH(1)
) cond264 (
    .clk(cond264_clk),
    .done(cond264_done),
    .in(cond264_in),
    .out(cond264_out),
    .reset(cond264_reset),
    .write_en(cond264_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire264 (
    .in(cond_wire264_in),
    .out(cond_wire264_out)
);
std_reg # (
    .WIDTH(1)
) cond265 (
    .clk(cond265_clk),
    .done(cond265_done),
    .in(cond265_in),
    .out(cond265_out),
    .reset(cond265_reset),
    .write_en(cond265_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire265 (
    .in(cond_wire265_in),
    .out(cond_wire265_out)
);
std_reg # (
    .WIDTH(1)
) cond266 (
    .clk(cond266_clk),
    .done(cond266_done),
    .in(cond266_in),
    .out(cond266_out),
    .reset(cond266_reset),
    .write_en(cond266_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire266 (
    .in(cond_wire266_in),
    .out(cond_wire266_out)
);
std_reg # (
    .WIDTH(1)
) cond267 (
    .clk(cond267_clk),
    .done(cond267_done),
    .in(cond267_in),
    .out(cond267_out),
    .reset(cond267_reset),
    .write_en(cond267_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire267 (
    .in(cond_wire267_in),
    .out(cond_wire267_out)
);
std_reg # (
    .WIDTH(1)
) cond268 (
    .clk(cond268_clk),
    .done(cond268_done),
    .in(cond268_in),
    .out(cond268_out),
    .reset(cond268_reset),
    .write_en(cond268_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire268 (
    .in(cond_wire268_in),
    .out(cond_wire268_out)
);
std_reg # (
    .WIDTH(1)
) cond269 (
    .clk(cond269_clk),
    .done(cond269_done),
    .in(cond269_in),
    .out(cond269_out),
    .reset(cond269_reset),
    .write_en(cond269_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire269 (
    .in(cond_wire269_in),
    .out(cond_wire269_out)
);
std_reg # (
    .WIDTH(1)
) cond270 (
    .clk(cond270_clk),
    .done(cond270_done),
    .in(cond270_in),
    .out(cond270_out),
    .reset(cond270_reset),
    .write_en(cond270_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire270 (
    .in(cond_wire270_in),
    .out(cond_wire270_out)
);
std_reg # (
    .WIDTH(1)
) cond271 (
    .clk(cond271_clk),
    .done(cond271_done),
    .in(cond271_in),
    .out(cond271_out),
    .reset(cond271_reset),
    .write_en(cond271_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire271 (
    .in(cond_wire271_in),
    .out(cond_wire271_out)
);
std_reg # (
    .WIDTH(1)
) cond272 (
    .clk(cond272_clk),
    .done(cond272_done),
    .in(cond272_in),
    .out(cond272_out),
    .reset(cond272_reset),
    .write_en(cond272_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire272 (
    .in(cond_wire272_in),
    .out(cond_wire272_out)
);
std_reg # (
    .WIDTH(1)
) cond273 (
    .clk(cond273_clk),
    .done(cond273_done),
    .in(cond273_in),
    .out(cond273_out),
    .reset(cond273_reset),
    .write_en(cond273_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire273 (
    .in(cond_wire273_in),
    .out(cond_wire273_out)
);
std_reg # (
    .WIDTH(1)
) cond274 (
    .clk(cond274_clk),
    .done(cond274_done),
    .in(cond274_in),
    .out(cond274_out),
    .reset(cond274_reset),
    .write_en(cond274_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire274 (
    .in(cond_wire274_in),
    .out(cond_wire274_out)
);
std_reg # (
    .WIDTH(1)
) cond275 (
    .clk(cond275_clk),
    .done(cond275_done),
    .in(cond275_in),
    .out(cond275_out),
    .reset(cond275_reset),
    .write_en(cond275_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire275 (
    .in(cond_wire275_in),
    .out(cond_wire275_out)
);
std_reg # (
    .WIDTH(1)
) cond276 (
    .clk(cond276_clk),
    .done(cond276_done),
    .in(cond276_in),
    .out(cond276_out),
    .reset(cond276_reset),
    .write_en(cond276_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire276 (
    .in(cond_wire276_in),
    .out(cond_wire276_out)
);
std_reg # (
    .WIDTH(1)
) cond277 (
    .clk(cond277_clk),
    .done(cond277_done),
    .in(cond277_in),
    .out(cond277_out),
    .reset(cond277_reset),
    .write_en(cond277_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire277 (
    .in(cond_wire277_in),
    .out(cond_wire277_out)
);
std_reg # (
    .WIDTH(1)
) cond278 (
    .clk(cond278_clk),
    .done(cond278_done),
    .in(cond278_in),
    .out(cond278_out),
    .reset(cond278_reset),
    .write_en(cond278_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire278 (
    .in(cond_wire278_in),
    .out(cond_wire278_out)
);
std_reg # (
    .WIDTH(1)
) cond279 (
    .clk(cond279_clk),
    .done(cond279_done),
    .in(cond279_in),
    .out(cond279_out),
    .reset(cond279_reset),
    .write_en(cond279_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire279 (
    .in(cond_wire279_in),
    .out(cond_wire279_out)
);
std_reg # (
    .WIDTH(1)
) cond280 (
    .clk(cond280_clk),
    .done(cond280_done),
    .in(cond280_in),
    .out(cond280_out),
    .reset(cond280_reset),
    .write_en(cond280_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire280 (
    .in(cond_wire280_in),
    .out(cond_wire280_out)
);
std_reg # (
    .WIDTH(1)
) cond281 (
    .clk(cond281_clk),
    .done(cond281_done),
    .in(cond281_in),
    .out(cond281_out),
    .reset(cond281_reset),
    .write_en(cond281_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire281 (
    .in(cond_wire281_in),
    .out(cond_wire281_out)
);
std_reg # (
    .WIDTH(1)
) cond282 (
    .clk(cond282_clk),
    .done(cond282_done),
    .in(cond282_in),
    .out(cond282_out),
    .reset(cond282_reset),
    .write_en(cond282_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire282 (
    .in(cond_wire282_in),
    .out(cond_wire282_out)
);
std_reg # (
    .WIDTH(1)
) cond283 (
    .clk(cond283_clk),
    .done(cond283_done),
    .in(cond283_in),
    .out(cond283_out),
    .reset(cond283_reset),
    .write_en(cond283_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire283 (
    .in(cond_wire283_in),
    .out(cond_wire283_out)
);
std_reg # (
    .WIDTH(1)
) cond284 (
    .clk(cond284_clk),
    .done(cond284_done),
    .in(cond284_in),
    .out(cond284_out),
    .reset(cond284_reset),
    .write_en(cond284_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire284 (
    .in(cond_wire284_in),
    .out(cond_wire284_out)
);
std_reg # (
    .WIDTH(1)
) cond285 (
    .clk(cond285_clk),
    .done(cond285_done),
    .in(cond285_in),
    .out(cond285_out),
    .reset(cond285_reset),
    .write_en(cond285_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire285 (
    .in(cond_wire285_in),
    .out(cond_wire285_out)
);
std_reg # (
    .WIDTH(1)
) cond286 (
    .clk(cond286_clk),
    .done(cond286_done),
    .in(cond286_in),
    .out(cond286_out),
    .reset(cond286_reset),
    .write_en(cond286_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire286 (
    .in(cond_wire286_in),
    .out(cond_wire286_out)
);
std_reg # (
    .WIDTH(1)
) cond287 (
    .clk(cond287_clk),
    .done(cond287_done),
    .in(cond287_in),
    .out(cond287_out),
    .reset(cond287_reset),
    .write_en(cond287_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire287 (
    .in(cond_wire287_in),
    .out(cond_wire287_out)
);
std_reg # (
    .WIDTH(1)
) cond288 (
    .clk(cond288_clk),
    .done(cond288_done),
    .in(cond288_in),
    .out(cond288_out),
    .reset(cond288_reset),
    .write_en(cond288_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire288 (
    .in(cond_wire288_in),
    .out(cond_wire288_out)
);
std_reg # (
    .WIDTH(1)
) cond289 (
    .clk(cond289_clk),
    .done(cond289_done),
    .in(cond289_in),
    .out(cond289_out),
    .reset(cond289_reset),
    .write_en(cond289_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire289 (
    .in(cond_wire289_in),
    .out(cond_wire289_out)
);
std_reg # (
    .WIDTH(1)
) cond290 (
    .clk(cond290_clk),
    .done(cond290_done),
    .in(cond290_in),
    .out(cond290_out),
    .reset(cond290_reset),
    .write_en(cond290_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire290 (
    .in(cond_wire290_in),
    .out(cond_wire290_out)
);
std_reg # (
    .WIDTH(1)
) cond291 (
    .clk(cond291_clk),
    .done(cond291_done),
    .in(cond291_in),
    .out(cond291_out),
    .reset(cond291_reset),
    .write_en(cond291_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire291 (
    .in(cond_wire291_in),
    .out(cond_wire291_out)
);
std_reg # (
    .WIDTH(1)
) cond292 (
    .clk(cond292_clk),
    .done(cond292_done),
    .in(cond292_in),
    .out(cond292_out),
    .reset(cond292_reset),
    .write_en(cond292_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire292 (
    .in(cond_wire292_in),
    .out(cond_wire292_out)
);
std_reg # (
    .WIDTH(1)
) cond293 (
    .clk(cond293_clk),
    .done(cond293_done),
    .in(cond293_in),
    .out(cond293_out),
    .reset(cond293_reset),
    .write_en(cond293_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire293 (
    .in(cond_wire293_in),
    .out(cond_wire293_out)
);
std_reg # (
    .WIDTH(1)
) cond294 (
    .clk(cond294_clk),
    .done(cond294_done),
    .in(cond294_in),
    .out(cond294_out),
    .reset(cond294_reset),
    .write_en(cond294_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire294 (
    .in(cond_wire294_in),
    .out(cond_wire294_out)
);
std_reg # (
    .WIDTH(1)
) cond295 (
    .clk(cond295_clk),
    .done(cond295_done),
    .in(cond295_in),
    .out(cond295_out),
    .reset(cond295_reset),
    .write_en(cond295_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire295 (
    .in(cond_wire295_in),
    .out(cond_wire295_out)
);
std_reg # (
    .WIDTH(1)
) cond296 (
    .clk(cond296_clk),
    .done(cond296_done),
    .in(cond296_in),
    .out(cond296_out),
    .reset(cond296_reset),
    .write_en(cond296_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire296 (
    .in(cond_wire296_in),
    .out(cond_wire296_out)
);
std_reg # (
    .WIDTH(1)
) cond297 (
    .clk(cond297_clk),
    .done(cond297_done),
    .in(cond297_in),
    .out(cond297_out),
    .reset(cond297_reset),
    .write_en(cond297_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire297 (
    .in(cond_wire297_in),
    .out(cond_wire297_out)
);
std_reg # (
    .WIDTH(1)
) cond298 (
    .clk(cond298_clk),
    .done(cond298_done),
    .in(cond298_in),
    .out(cond298_out),
    .reset(cond298_reset),
    .write_en(cond298_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire298 (
    .in(cond_wire298_in),
    .out(cond_wire298_out)
);
std_reg # (
    .WIDTH(1)
) cond299 (
    .clk(cond299_clk),
    .done(cond299_done),
    .in(cond299_in),
    .out(cond299_out),
    .reset(cond299_reset),
    .write_en(cond299_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire299 (
    .in(cond_wire299_in),
    .out(cond_wire299_out)
);
std_reg # (
    .WIDTH(1)
) cond300 (
    .clk(cond300_clk),
    .done(cond300_done),
    .in(cond300_in),
    .out(cond300_out),
    .reset(cond300_reset),
    .write_en(cond300_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire300 (
    .in(cond_wire300_in),
    .out(cond_wire300_out)
);
std_reg # (
    .WIDTH(1)
) cond301 (
    .clk(cond301_clk),
    .done(cond301_done),
    .in(cond301_in),
    .out(cond301_out),
    .reset(cond301_reset),
    .write_en(cond301_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire301 (
    .in(cond_wire301_in),
    .out(cond_wire301_out)
);
std_reg # (
    .WIDTH(1)
) cond302 (
    .clk(cond302_clk),
    .done(cond302_done),
    .in(cond302_in),
    .out(cond302_out),
    .reset(cond302_reset),
    .write_en(cond302_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire302 (
    .in(cond_wire302_in),
    .out(cond_wire302_out)
);
std_reg # (
    .WIDTH(1)
) cond303 (
    .clk(cond303_clk),
    .done(cond303_done),
    .in(cond303_in),
    .out(cond303_out),
    .reset(cond303_reset),
    .write_en(cond303_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire303 (
    .in(cond_wire303_in),
    .out(cond_wire303_out)
);
std_reg # (
    .WIDTH(1)
) cond304 (
    .clk(cond304_clk),
    .done(cond304_done),
    .in(cond304_in),
    .out(cond304_out),
    .reset(cond304_reset),
    .write_en(cond304_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire304 (
    .in(cond_wire304_in),
    .out(cond_wire304_out)
);
std_reg # (
    .WIDTH(1)
) cond305 (
    .clk(cond305_clk),
    .done(cond305_done),
    .in(cond305_in),
    .out(cond305_out),
    .reset(cond305_reset),
    .write_en(cond305_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire305 (
    .in(cond_wire305_in),
    .out(cond_wire305_out)
);
std_reg # (
    .WIDTH(1)
) cond306 (
    .clk(cond306_clk),
    .done(cond306_done),
    .in(cond306_in),
    .out(cond306_out),
    .reset(cond306_reset),
    .write_en(cond306_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire306 (
    .in(cond_wire306_in),
    .out(cond_wire306_out)
);
std_reg # (
    .WIDTH(1)
) cond307 (
    .clk(cond307_clk),
    .done(cond307_done),
    .in(cond307_in),
    .out(cond307_out),
    .reset(cond307_reset),
    .write_en(cond307_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire307 (
    .in(cond_wire307_in),
    .out(cond_wire307_out)
);
std_reg # (
    .WIDTH(1)
) cond308 (
    .clk(cond308_clk),
    .done(cond308_done),
    .in(cond308_in),
    .out(cond308_out),
    .reset(cond308_reset),
    .write_en(cond308_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire308 (
    .in(cond_wire308_in),
    .out(cond_wire308_out)
);
std_reg # (
    .WIDTH(1)
) cond309 (
    .clk(cond309_clk),
    .done(cond309_done),
    .in(cond309_in),
    .out(cond309_out),
    .reset(cond309_reset),
    .write_en(cond309_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire309 (
    .in(cond_wire309_in),
    .out(cond_wire309_out)
);
std_reg # (
    .WIDTH(1)
) cond310 (
    .clk(cond310_clk),
    .done(cond310_done),
    .in(cond310_in),
    .out(cond310_out),
    .reset(cond310_reset),
    .write_en(cond310_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire310 (
    .in(cond_wire310_in),
    .out(cond_wire310_out)
);
std_reg # (
    .WIDTH(1)
) cond311 (
    .clk(cond311_clk),
    .done(cond311_done),
    .in(cond311_in),
    .out(cond311_out),
    .reset(cond311_reset),
    .write_en(cond311_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire311 (
    .in(cond_wire311_in),
    .out(cond_wire311_out)
);
std_reg # (
    .WIDTH(1)
) cond312 (
    .clk(cond312_clk),
    .done(cond312_done),
    .in(cond312_in),
    .out(cond312_out),
    .reset(cond312_reset),
    .write_en(cond312_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire312 (
    .in(cond_wire312_in),
    .out(cond_wire312_out)
);
std_reg # (
    .WIDTH(1)
) cond313 (
    .clk(cond313_clk),
    .done(cond313_done),
    .in(cond313_in),
    .out(cond313_out),
    .reset(cond313_reset),
    .write_en(cond313_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire313 (
    .in(cond_wire313_in),
    .out(cond_wire313_out)
);
std_reg # (
    .WIDTH(1)
) cond314 (
    .clk(cond314_clk),
    .done(cond314_done),
    .in(cond314_in),
    .out(cond314_out),
    .reset(cond314_reset),
    .write_en(cond314_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire314 (
    .in(cond_wire314_in),
    .out(cond_wire314_out)
);
std_reg # (
    .WIDTH(1)
) cond315 (
    .clk(cond315_clk),
    .done(cond315_done),
    .in(cond315_in),
    .out(cond315_out),
    .reset(cond315_reset),
    .write_en(cond315_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire315 (
    .in(cond_wire315_in),
    .out(cond_wire315_out)
);
std_reg # (
    .WIDTH(1)
) cond316 (
    .clk(cond316_clk),
    .done(cond316_done),
    .in(cond316_in),
    .out(cond316_out),
    .reset(cond316_reset),
    .write_en(cond316_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire316 (
    .in(cond_wire316_in),
    .out(cond_wire316_out)
);
std_reg # (
    .WIDTH(1)
) cond317 (
    .clk(cond317_clk),
    .done(cond317_done),
    .in(cond317_in),
    .out(cond317_out),
    .reset(cond317_reset),
    .write_en(cond317_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire317 (
    .in(cond_wire317_in),
    .out(cond_wire317_out)
);
std_reg # (
    .WIDTH(1)
) cond318 (
    .clk(cond318_clk),
    .done(cond318_done),
    .in(cond318_in),
    .out(cond318_out),
    .reset(cond318_reset),
    .write_en(cond318_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire318 (
    .in(cond_wire318_in),
    .out(cond_wire318_out)
);
std_reg # (
    .WIDTH(1)
) cond319 (
    .clk(cond319_clk),
    .done(cond319_done),
    .in(cond319_in),
    .out(cond319_out),
    .reset(cond319_reset),
    .write_en(cond319_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire319 (
    .in(cond_wire319_in),
    .out(cond_wire319_out)
);
std_reg # (
    .WIDTH(1)
) cond320 (
    .clk(cond320_clk),
    .done(cond320_done),
    .in(cond320_in),
    .out(cond320_out),
    .reset(cond320_reset),
    .write_en(cond320_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire320 (
    .in(cond_wire320_in),
    .out(cond_wire320_out)
);
std_reg # (
    .WIDTH(1)
) cond321 (
    .clk(cond321_clk),
    .done(cond321_done),
    .in(cond321_in),
    .out(cond321_out),
    .reset(cond321_reset),
    .write_en(cond321_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire321 (
    .in(cond_wire321_in),
    .out(cond_wire321_out)
);
std_reg # (
    .WIDTH(1)
) cond322 (
    .clk(cond322_clk),
    .done(cond322_done),
    .in(cond322_in),
    .out(cond322_out),
    .reset(cond322_reset),
    .write_en(cond322_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire322 (
    .in(cond_wire322_in),
    .out(cond_wire322_out)
);
std_reg # (
    .WIDTH(1)
) cond323 (
    .clk(cond323_clk),
    .done(cond323_done),
    .in(cond323_in),
    .out(cond323_out),
    .reset(cond323_reset),
    .write_en(cond323_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire323 (
    .in(cond_wire323_in),
    .out(cond_wire323_out)
);
std_reg # (
    .WIDTH(1)
) cond324 (
    .clk(cond324_clk),
    .done(cond324_done),
    .in(cond324_in),
    .out(cond324_out),
    .reset(cond324_reset),
    .write_en(cond324_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire324 (
    .in(cond_wire324_in),
    .out(cond_wire324_out)
);
std_reg # (
    .WIDTH(1)
) cond325 (
    .clk(cond325_clk),
    .done(cond325_done),
    .in(cond325_in),
    .out(cond325_out),
    .reset(cond325_reset),
    .write_en(cond325_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire325 (
    .in(cond_wire325_in),
    .out(cond_wire325_out)
);
std_reg # (
    .WIDTH(1)
) cond326 (
    .clk(cond326_clk),
    .done(cond326_done),
    .in(cond326_in),
    .out(cond326_out),
    .reset(cond326_reset),
    .write_en(cond326_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire326 (
    .in(cond_wire326_in),
    .out(cond_wire326_out)
);
std_reg # (
    .WIDTH(1)
) cond327 (
    .clk(cond327_clk),
    .done(cond327_done),
    .in(cond327_in),
    .out(cond327_out),
    .reset(cond327_reset),
    .write_en(cond327_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire327 (
    .in(cond_wire327_in),
    .out(cond_wire327_out)
);
std_reg # (
    .WIDTH(1)
) cond328 (
    .clk(cond328_clk),
    .done(cond328_done),
    .in(cond328_in),
    .out(cond328_out),
    .reset(cond328_reset),
    .write_en(cond328_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire328 (
    .in(cond_wire328_in),
    .out(cond_wire328_out)
);
std_reg # (
    .WIDTH(1)
) cond329 (
    .clk(cond329_clk),
    .done(cond329_done),
    .in(cond329_in),
    .out(cond329_out),
    .reset(cond329_reset),
    .write_en(cond329_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire329 (
    .in(cond_wire329_in),
    .out(cond_wire329_out)
);
std_reg # (
    .WIDTH(1)
) cond330 (
    .clk(cond330_clk),
    .done(cond330_done),
    .in(cond330_in),
    .out(cond330_out),
    .reset(cond330_reset),
    .write_en(cond330_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire330 (
    .in(cond_wire330_in),
    .out(cond_wire330_out)
);
std_reg # (
    .WIDTH(1)
) cond331 (
    .clk(cond331_clk),
    .done(cond331_done),
    .in(cond331_in),
    .out(cond331_out),
    .reset(cond331_reset),
    .write_en(cond331_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire331 (
    .in(cond_wire331_in),
    .out(cond_wire331_out)
);
std_reg # (
    .WIDTH(1)
) cond332 (
    .clk(cond332_clk),
    .done(cond332_done),
    .in(cond332_in),
    .out(cond332_out),
    .reset(cond332_reset),
    .write_en(cond332_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire332 (
    .in(cond_wire332_in),
    .out(cond_wire332_out)
);
std_reg # (
    .WIDTH(1)
) cond333 (
    .clk(cond333_clk),
    .done(cond333_done),
    .in(cond333_in),
    .out(cond333_out),
    .reset(cond333_reset),
    .write_en(cond333_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire333 (
    .in(cond_wire333_in),
    .out(cond_wire333_out)
);
std_reg # (
    .WIDTH(1)
) cond334 (
    .clk(cond334_clk),
    .done(cond334_done),
    .in(cond334_in),
    .out(cond334_out),
    .reset(cond334_reset),
    .write_en(cond334_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire334 (
    .in(cond_wire334_in),
    .out(cond_wire334_out)
);
std_reg # (
    .WIDTH(1)
) cond335 (
    .clk(cond335_clk),
    .done(cond335_done),
    .in(cond335_in),
    .out(cond335_out),
    .reset(cond335_reset),
    .write_en(cond335_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire335 (
    .in(cond_wire335_in),
    .out(cond_wire335_out)
);
std_reg # (
    .WIDTH(1)
) cond336 (
    .clk(cond336_clk),
    .done(cond336_done),
    .in(cond336_in),
    .out(cond336_out),
    .reset(cond336_reset),
    .write_en(cond336_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire336 (
    .in(cond_wire336_in),
    .out(cond_wire336_out)
);
std_reg # (
    .WIDTH(1)
) cond337 (
    .clk(cond337_clk),
    .done(cond337_done),
    .in(cond337_in),
    .out(cond337_out),
    .reset(cond337_reset),
    .write_en(cond337_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire337 (
    .in(cond_wire337_in),
    .out(cond_wire337_out)
);
std_reg # (
    .WIDTH(1)
) cond338 (
    .clk(cond338_clk),
    .done(cond338_done),
    .in(cond338_in),
    .out(cond338_out),
    .reset(cond338_reset),
    .write_en(cond338_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire338 (
    .in(cond_wire338_in),
    .out(cond_wire338_out)
);
std_reg # (
    .WIDTH(1)
) cond339 (
    .clk(cond339_clk),
    .done(cond339_done),
    .in(cond339_in),
    .out(cond339_out),
    .reset(cond339_reset),
    .write_en(cond339_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire339 (
    .in(cond_wire339_in),
    .out(cond_wire339_out)
);
std_reg # (
    .WIDTH(1)
) cond340 (
    .clk(cond340_clk),
    .done(cond340_done),
    .in(cond340_in),
    .out(cond340_out),
    .reset(cond340_reset),
    .write_en(cond340_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire340 (
    .in(cond_wire340_in),
    .out(cond_wire340_out)
);
std_reg # (
    .WIDTH(1)
) cond341 (
    .clk(cond341_clk),
    .done(cond341_done),
    .in(cond341_in),
    .out(cond341_out),
    .reset(cond341_reset),
    .write_en(cond341_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire341 (
    .in(cond_wire341_in),
    .out(cond_wire341_out)
);
std_reg # (
    .WIDTH(1)
) cond342 (
    .clk(cond342_clk),
    .done(cond342_done),
    .in(cond342_in),
    .out(cond342_out),
    .reset(cond342_reset),
    .write_en(cond342_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire342 (
    .in(cond_wire342_in),
    .out(cond_wire342_out)
);
std_reg # (
    .WIDTH(1)
) cond343 (
    .clk(cond343_clk),
    .done(cond343_done),
    .in(cond343_in),
    .out(cond343_out),
    .reset(cond343_reset),
    .write_en(cond343_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire343 (
    .in(cond_wire343_in),
    .out(cond_wire343_out)
);
std_reg # (
    .WIDTH(1)
) cond344 (
    .clk(cond344_clk),
    .done(cond344_done),
    .in(cond344_in),
    .out(cond344_out),
    .reset(cond344_reset),
    .write_en(cond344_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire344 (
    .in(cond_wire344_in),
    .out(cond_wire344_out)
);
std_reg # (
    .WIDTH(1)
) cond345 (
    .clk(cond345_clk),
    .done(cond345_done),
    .in(cond345_in),
    .out(cond345_out),
    .reset(cond345_reset),
    .write_en(cond345_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire345 (
    .in(cond_wire345_in),
    .out(cond_wire345_out)
);
std_reg # (
    .WIDTH(1)
) cond346 (
    .clk(cond346_clk),
    .done(cond346_done),
    .in(cond346_in),
    .out(cond346_out),
    .reset(cond346_reset),
    .write_en(cond346_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire346 (
    .in(cond_wire346_in),
    .out(cond_wire346_out)
);
std_reg # (
    .WIDTH(1)
) cond347 (
    .clk(cond347_clk),
    .done(cond347_done),
    .in(cond347_in),
    .out(cond347_out),
    .reset(cond347_reset),
    .write_en(cond347_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire347 (
    .in(cond_wire347_in),
    .out(cond_wire347_out)
);
std_reg # (
    .WIDTH(1)
) cond348 (
    .clk(cond348_clk),
    .done(cond348_done),
    .in(cond348_in),
    .out(cond348_out),
    .reset(cond348_reset),
    .write_en(cond348_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire348 (
    .in(cond_wire348_in),
    .out(cond_wire348_out)
);
std_reg # (
    .WIDTH(1)
) cond349 (
    .clk(cond349_clk),
    .done(cond349_done),
    .in(cond349_in),
    .out(cond349_out),
    .reset(cond349_reset),
    .write_en(cond349_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire349 (
    .in(cond_wire349_in),
    .out(cond_wire349_out)
);
std_reg # (
    .WIDTH(1)
) cond350 (
    .clk(cond350_clk),
    .done(cond350_done),
    .in(cond350_in),
    .out(cond350_out),
    .reset(cond350_reset),
    .write_en(cond350_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire350 (
    .in(cond_wire350_in),
    .out(cond_wire350_out)
);
std_reg # (
    .WIDTH(1)
) cond351 (
    .clk(cond351_clk),
    .done(cond351_done),
    .in(cond351_in),
    .out(cond351_out),
    .reset(cond351_reset),
    .write_en(cond351_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire351 (
    .in(cond_wire351_in),
    .out(cond_wire351_out)
);
std_reg # (
    .WIDTH(1)
) cond352 (
    .clk(cond352_clk),
    .done(cond352_done),
    .in(cond352_in),
    .out(cond352_out),
    .reset(cond352_reset),
    .write_en(cond352_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire352 (
    .in(cond_wire352_in),
    .out(cond_wire352_out)
);
std_reg # (
    .WIDTH(1)
) cond353 (
    .clk(cond353_clk),
    .done(cond353_done),
    .in(cond353_in),
    .out(cond353_out),
    .reset(cond353_reset),
    .write_en(cond353_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire353 (
    .in(cond_wire353_in),
    .out(cond_wire353_out)
);
std_reg # (
    .WIDTH(1)
) cond354 (
    .clk(cond354_clk),
    .done(cond354_done),
    .in(cond354_in),
    .out(cond354_out),
    .reset(cond354_reset),
    .write_en(cond354_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire354 (
    .in(cond_wire354_in),
    .out(cond_wire354_out)
);
std_reg # (
    .WIDTH(1)
) cond355 (
    .clk(cond355_clk),
    .done(cond355_done),
    .in(cond355_in),
    .out(cond355_out),
    .reset(cond355_reset),
    .write_en(cond355_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire355 (
    .in(cond_wire355_in),
    .out(cond_wire355_out)
);
std_reg # (
    .WIDTH(1)
) cond356 (
    .clk(cond356_clk),
    .done(cond356_done),
    .in(cond356_in),
    .out(cond356_out),
    .reset(cond356_reset),
    .write_en(cond356_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire356 (
    .in(cond_wire356_in),
    .out(cond_wire356_out)
);
std_reg # (
    .WIDTH(1)
) cond357 (
    .clk(cond357_clk),
    .done(cond357_done),
    .in(cond357_in),
    .out(cond357_out),
    .reset(cond357_reset),
    .write_en(cond357_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire357 (
    .in(cond_wire357_in),
    .out(cond_wire357_out)
);
std_reg # (
    .WIDTH(1)
) cond358 (
    .clk(cond358_clk),
    .done(cond358_done),
    .in(cond358_in),
    .out(cond358_out),
    .reset(cond358_reset),
    .write_en(cond358_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire358 (
    .in(cond_wire358_in),
    .out(cond_wire358_out)
);
std_reg # (
    .WIDTH(1)
) cond359 (
    .clk(cond359_clk),
    .done(cond359_done),
    .in(cond359_in),
    .out(cond359_out),
    .reset(cond359_reset),
    .write_en(cond359_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire359 (
    .in(cond_wire359_in),
    .out(cond_wire359_out)
);
std_reg # (
    .WIDTH(1)
) cond360 (
    .clk(cond360_clk),
    .done(cond360_done),
    .in(cond360_in),
    .out(cond360_out),
    .reset(cond360_reset),
    .write_en(cond360_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire360 (
    .in(cond_wire360_in),
    .out(cond_wire360_out)
);
std_reg # (
    .WIDTH(1)
) cond361 (
    .clk(cond361_clk),
    .done(cond361_done),
    .in(cond361_in),
    .out(cond361_out),
    .reset(cond361_reset),
    .write_en(cond361_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire361 (
    .in(cond_wire361_in),
    .out(cond_wire361_out)
);
std_reg # (
    .WIDTH(1)
) cond362 (
    .clk(cond362_clk),
    .done(cond362_done),
    .in(cond362_in),
    .out(cond362_out),
    .reset(cond362_reset),
    .write_en(cond362_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire362 (
    .in(cond_wire362_in),
    .out(cond_wire362_out)
);
std_reg # (
    .WIDTH(1)
) cond363 (
    .clk(cond363_clk),
    .done(cond363_done),
    .in(cond363_in),
    .out(cond363_out),
    .reset(cond363_reset),
    .write_en(cond363_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire363 (
    .in(cond_wire363_in),
    .out(cond_wire363_out)
);
std_reg # (
    .WIDTH(1)
) cond364 (
    .clk(cond364_clk),
    .done(cond364_done),
    .in(cond364_in),
    .out(cond364_out),
    .reset(cond364_reset),
    .write_en(cond364_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire364 (
    .in(cond_wire364_in),
    .out(cond_wire364_out)
);
std_reg # (
    .WIDTH(1)
) cond365 (
    .clk(cond365_clk),
    .done(cond365_done),
    .in(cond365_in),
    .out(cond365_out),
    .reset(cond365_reset),
    .write_en(cond365_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire365 (
    .in(cond_wire365_in),
    .out(cond_wire365_out)
);
std_reg # (
    .WIDTH(1)
) cond366 (
    .clk(cond366_clk),
    .done(cond366_done),
    .in(cond366_in),
    .out(cond366_out),
    .reset(cond366_reset),
    .write_en(cond366_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire366 (
    .in(cond_wire366_in),
    .out(cond_wire366_out)
);
std_reg # (
    .WIDTH(1)
) cond367 (
    .clk(cond367_clk),
    .done(cond367_done),
    .in(cond367_in),
    .out(cond367_out),
    .reset(cond367_reset),
    .write_en(cond367_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire367 (
    .in(cond_wire367_in),
    .out(cond_wire367_out)
);
std_reg # (
    .WIDTH(1)
) cond368 (
    .clk(cond368_clk),
    .done(cond368_done),
    .in(cond368_in),
    .out(cond368_out),
    .reset(cond368_reset),
    .write_en(cond368_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire368 (
    .in(cond_wire368_in),
    .out(cond_wire368_out)
);
std_reg # (
    .WIDTH(1)
) cond369 (
    .clk(cond369_clk),
    .done(cond369_done),
    .in(cond369_in),
    .out(cond369_out),
    .reset(cond369_reset),
    .write_en(cond369_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire369 (
    .in(cond_wire369_in),
    .out(cond_wire369_out)
);
std_reg # (
    .WIDTH(1)
) cond370 (
    .clk(cond370_clk),
    .done(cond370_done),
    .in(cond370_in),
    .out(cond370_out),
    .reset(cond370_reset),
    .write_en(cond370_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire370 (
    .in(cond_wire370_in),
    .out(cond_wire370_out)
);
std_reg # (
    .WIDTH(1)
) cond371 (
    .clk(cond371_clk),
    .done(cond371_done),
    .in(cond371_in),
    .out(cond371_out),
    .reset(cond371_reset),
    .write_en(cond371_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire371 (
    .in(cond_wire371_in),
    .out(cond_wire371_out)
);
std_reg # (
    .WIDTH(1)
) cond372 (
    .clk(cond372_clk),
    .done(cond372_done),
    .in(cond372_in),
    .out(cond372_out),
    .reset(cond372_reset),
    .write_en(cond372_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire372 (
    .in(cond_wire372_in),
    .out(cond_wire372_out)
);
std_reg # (
    .WIDTH(1)
) cond373 (
    .clk(cond373_clk),
    .done(cond373_done),
    .in(cond373_in),
    .out(cond373_out),
    .reset(cond373_reset),
    .write_en(cond373_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire373 (
    .in(cond_wire373_in),
    .out(cond_wire373_out)
);
std_reg # (
    .WIDTH(1)
) cond374 (
    .clk(cond374_clk),
    .done(cond374_done),
    .in(cond374_in),
    .out(cond374_out),
    .reset(cond374_reset),
    .write_en(cond374_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire374 (
    .in(cond_wire374_in),
    .out(cond_wire374_out)
);
std_reg # (
    .WIDTH(1)
) cond375 (
    .clk(cond375_clk),
    .done(cond375_done),
    .in(cond375_in),
    .out(cond375_out),
    .reset(cond375_reset),
    .write_en(cond375_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire375 (
    .in(cond_wire375_in),
    .out(cond_wire375_out)
);
std_reg # (
    .WIDTH(1)
) cond376 (
    .clk(cond376_clk),
    .done(cond376_done),
    .in(cond376_in),
    .out(cond376_out),
    .reset(cond376_reset),
    .write_en(cond376_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire376 (
    .in(cond_wire376_in),
    .out(cond_wire376_out)
);
std_reg # (
    .WIDTH(1)
) cond377 (
    .clk(cond377_clk),
    .done(cond377_done),
    .in(cond377_in),
    .out(cond377_out),
    .reset(cond377_reset),
    .write_en(cond377_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire377 (
    .in(cond_wire377_in),
    .out(cond_wire377_out)
);
std_reg # (
    .WIDTH(1)
) cond378 (
    .clk(cond378_clk),
    .done(cond378_done),
    .in(cond378_in),
    .out(cond378_out),
    .reset(cond378_reset),
    .write_en(cond378_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire378 (
    .in(cond_wire378_in),
    .out(cond_wire378_out)
);
std_reg # (
    .WIDTH(1)
) cond379 (
    .clk(cond379_clk),
    .done(cond379_done),
    .in(cond379_in),
    .out(cond379_out),
    .reset(cond379_reset),
    .write_en(cond379_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire379 (
    .in(cond_wire379_in),
    .out(cond_wire379_out)
);
std_reg # (
    .WIDTH(1)
) cond380 (
    .clk(cond380_clk),
    .done(cond380_done),
    .in(cond380_in),
    .out(cond380_out),
    .reset(cond380_reset),
    .write_en(cond380_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire380 (
    .in(cond_wire380_in),
    .out(cond_wire380_out)
);
std_reg # (
    .WIDTH(1)
) cond381 (
    .clk(cond381_clk),
    .done(cond381_done),
    .in(cond381_in),
    .out(cond381_out),
    .reset(cond381_reset),
    .write_en(cond381_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire381 (
    .in(cond_wire381_in),
    .out(cond_wire381_out)
);
std_reg # (
    .WIDTH(1)
) cond382 (
    .clk(cond382_clk),
    .done(cond382_done),
    .in(cond382_in),
    .out(cond382_out),
    .reset(cond382_reset),
    .write_en(cond382_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire382 (
    .in(cond_wire382_in),
    .out(cond_wire382_out)
);
std_reg # (
    .WIDTH(1)
) cond383 (
    .clk(cond383_clk),
    .done(cond383_done),
    .in(cond383_in),
    .out(cond383_out),
    .reset(cond383_reset),
    .write_en(cond383_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire383 (
    .in(cond_wire383_in),
    .out(cond_wire383_out)
);
std_reg # (
    .WIDTH(1)
) cond384 (
    .clk(cond384_clk),
    .done(cond384_done),
    .in(cond384_in),
    .out(cond384_out),
    .reset(cond384_reset),
    .write_en(cond384_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire384 (
    .in(cond_wire384_in),
    .out(cond_wire384_out)
);
std_reg # (
    .WIDTH(1)
) cond385 (
    .clk(cond385_clk),
    .done(cond385_done),
    .in(cond385_in),
    .out(cond385_out),
    .reset(cond385_reset),
    .write_en(cond385_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire385 (
    .in(cond_wire385_in),
    .out(cond_wire385_out)
);
std_reg # (
    .WIDTH(1)
) cond386 (
    .clk(cond386_clk),
    .done(cond386_done),
    .in(cond386_in),
    .out(cond386_out),
    .reset(cond386_reset),
    .write_en(cond386_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire386 (
    .in(cond_wire386_in),
    .out(cond_wire386_out)
);
std_reg # (
    .WIDTH(1)
) cond387 (
    .clk(cond387_clk),
    .done(cond387_done),
    .in(cond387_in),
    .out(cond387_out),
    .reset(cond387_reset),
    .write_en(cond387_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire387 (
    .in(cond_wire387_in),
    .out(cond_wire387_out)
);
std_reg # (
    .WIDTH(1)
) cond388 (
    .clk(cond388_clk),
    .done(cond388_done),
    .in(cond388_in),
    .out(cond388_out),
    .reset(cond388_reset),
    .write_en(cond388_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire388 (
    .in(cond_wire388_in),
    .out(cond_wire388_out)
);
std_reg # (
    .WIDTH(1)
) cond389 (
    .clk(cond389_clk),
    .done(cond389_done),
    .in(cond389_in),
    .out(cond389_out),
    .reset(cond389_reset),
    .write_en(cond389_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire389 (
    .in(cond_wire389_in),
    .out(cond_wire389_out)
);
std_reg # (
    .WIDTH(1)
) cond390 (
    .clk(cond390_clk),
    .done(cond390_done),
    .in(cond390_in),
    .out(cond390_out),
    .reset(cond390_reset),
    .write_en(cond390_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire390 (
    .in(cond_wire390_in),
    .out(cond_wire390_out)
);
std_reg # (
    .WIDTH(1)
) cond391 (
    .clk(cond391_clk),
    .done(cond391_done),
    .in(cond391_in),
    .out(cond391_out),
    .reset(cond391_reset),
    .write_en(cond391_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire391 (
    .in(cond_wire391_in),
    .out(cond_wire391_out)
);
std_reg # (
    .WIDTH(1)
) cond392 (
    .clk(cond392_clk),
    .done(cond392_done),
    .in(cond392_in),
    .out(cond392_out),
    .reset(cond392_reset),
    .write_en(cond392_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire392 (
    .in(cond_wire392_in),
    .out(cond_wire392_out)
);
std_reg # (
    .WIDTH(1)
) cond393 (
    .clk(cond393_clk),
    .done(cond393_done),
    .in(cond393_in),
    .out(cond393_out),
    .reset(cond393_reset),
    .write_en(cond393_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire393 (
    .in(cond_wire393_in),
    .out(cond_wire393_out)
);
std_reg # (
    .WIDTH(1)
) cond394 (
    .clk(cond394_clk),
    .done(cond394_done),
    .in(cond394_in),
    .out(cond394_out),
    .reset(cond394_reset),
    .write_en(cond394_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire394 (
    .in(cond_wire394_in),
    .out(cond_wire394_out)
);
std_reg # (
    .WIDTH(1)
) cond395 (
    .clk(cond395_clk),
    .done(cond395_done),
    .in(cond395_in),
    .out(cond395_out),
    .reset(cond395_reset),
    .write_en(cond395_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire395 (
    .in(cond_wire395_in),
    .out(cond_wire395_out)
);
std_reg # (
    .WIDTH(1)
) cond396 (
    .clk(cond396_clk),
    .done(cond396_done),
    .in(cond396_in),
    .out(cond396_out),
    .reset(cond396_reset),
    .write_en(cond396_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire396 (
    .in(cond_wire396_in),
    .out(cond_wire396_out)
);
std_reg # (
    .WIDTH(1)
) cond397 (
    .clk(cond397_clk),
    .done(cond397_done),
    .in(cond397_in),
    .out(cond397_out),
    .reset(cond397_reset),
    .write_en(cond397_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire397 (
    .in(cond_wire397_in),
    .out(cond_wire397_out)
);
std_reg # (
    .WIDTH(1)
) cond398 (
    .clk(cond398_clk),
    .done(cond398_done),
    .in(cond398_in),
    .out(cond398_out),
    .reset(cond398_reset),
    .write_en(cond398_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire398 (
    .in(cond_wire398_in),
    .out(cond_wire398_out)
);
std_reg # (
    .WIDTH(1)
) cond399 (
    .clk(cond399_clk),
    .done(cond399_done),
    .in(cond399_in),
    .out(cond399_out),
    .reset(cond399_reset),
    .write_en(cond399_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire399 (
    .in(cond_wire399_in),
    .out(cond_wire399_out)
);
std_reg # (
    .WIDTH(1)
) cond400 (
    .clk(cond400_clk),
    .done(cond400_done),
    .in(cond400_in),
    .out(cond400_out),
    .reset(cond400_reset),
    .write_en(cond400_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire400 (
    .in(cond_wire400_in),
    .out(cond_wire400_out)
);
std_reg # (
    .WIDTH(1)
) cond401 (
    .clk(cond401_clk),
    .done(cond401_done),
    .in(cond401_in),
    .out(cond401_out),
    .reset(cond401_reset),
    .write_en(cond401_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire401 (
    .in(cond_wire401_in),
    .out(cond_wire401_out)
);
std_reg # (
    .WIDTH(1)
) cond402 (
    .clk(cond402_clk),
    .done(cond402_done),
    .in(cond402_in),
    .out(cond402_out),
    .reset(cond402_reset),
    .write_en(cond402_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire402 (
    .in(cond_wire402_in),
    .out(cond_wire402_out)
);
std_reg # (
    .WIDTH(1)
) cond403 (
    .clk(cond403_clk),
    .done(cond403_done),
    .in(cond403_in),
    .out(cond403_out),
    .reset(cond403_reset),
    .write_en(cond403_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire403 (
    .in(cond_wire403_in),
    .out(cond_wire403_out)
);
std_reg # (
    .WIDTH(1)
) cond404 (
    .clk(cond404_clk),
    .done(cond404_done),
    .in(cond404_in),
    .out(cond404_out),
    .reset(cond404_reset),
    .write_en(cond404_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire404 (
    .in(cond_wire404_in),
    .out(cond_wire404_out)
);
std_reg # (
    .WIDTH(1)
) cond405 (
    .clk(cond405_clk),
    .done(cond405_done),
    .in(cond405_in),
    .out(cond405_out),
    .reset(cond405_reset),
    .write_en(cond405_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire405 (
    .in(cond_wire405_in),
    .out(cond_wire405_out)
);
std_reg # (
    .WIDTH(1)
) cond406 (
    .clk(cond406_clk),
    .done(cond406_done),
    .in(cond406_in),
    .out(cond406_out),
    .reset(cond406_reset),
    .write_en(cond406_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire406 (
    .in(cond_wire406_in),
    .out(cond_wire406_out)
);
std_reg # (
    .WIDTH(1)
) cond407 (
    .clk(cond407_clk),
    .done(cond407_done),
    .in(cond407_in),
    .out(cond407_out),
    .reset(cond407_reset),
    .write_en(cond407_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire407 (
    .in(cond_wire407_in),
    .out(cond_wire407_out)
);
std_reg # (
    .WIDTH(1)
) cond408 (
    .clk(cond408_clk),
    .done(cond408_done),
    .in(cond408_in),
    .out(cond408_out),
    .reset(cond408_reset),
    .write_en(cond408_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire408 (
    .in(cond_wire408_in),
    .out(cond_wire408_out)
);
std_reg # (
    .WIDTH(1)
) cond409 (
    .clk(cond409_clk),
    .done(cond409_done),
    .in(cond409_in),
    .out(cond409_out),
    .reset(cond409_reset),
    .write_en(cond409_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire409 (
    .in(cond_wire409_in),
    .out(cond_wire409_out)
);
std_reg # (
    .WIDTH(1)
) cond410 (
    .clk(cond410_clk),
    .done(cond410_done),
    .in(cond410_in),
    .out(cond410_out),
    .reset(cond410_reset),
    .write_en(cond410_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire410 (
    .in(cond_wire410_in),
    .out(cond_wire410_out)
);
std_reg # (
    .WIDTH(1)
) cond411 (
    .clk(cond411_clk),
    .done(cond411_done),
    .in(cond411_in),
    .out(cond411_out),
    .reset(cond411_reset),
    .write_en(cond411_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire411 (
    .in(cond_wire411_in),
    .out(cond_wire411_out)
);
std_reg # (
    .WIDTH(1)
) cond412 (
    .clk(cond412_clk),
    .done(cond412_done),
    .in(cond412_in),
    .out(cond412_out),
    .reset(cond412_reset),
    .write_en(cond412_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire412 (
    .in(cond_wire412_in),
    .out(cond_wire412_out)
);
std_reg # (
    .WIDTH(1)
) cond413 (
    .clk(cond413_clk),
    .done(cond413_done),
    .in(cond413_in),
    .out(cond413_out),
    .reset(cond413_reset),
    .write_en(cond413_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire413 (
    .in(cond_wire413_in),
    .out(cond_wire413_out)
);
std_reg # (
    .WIDTH(1)
) cond414 (
    .clk(cond414_clk),
    .done(cond414_done),
    .in(cond414_in),
    .out(cond414_out),
    .reset(cond414_reset),
    .write_en(cond414_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire414 (
    .in(cond_wire414_in),
    .out(cond_wire414_out)
);
std_reg # (
    .WIDTH(1)
) cond415 (
    .clk(cond415_clk),
    .done(cond415_done),
    .in(cond415_in),
    .out(cond415_out),
    .reset(cond415_reset),
    .write_en(cond415_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire415 (
    .in(cond_wire415_in),
    .out(cond_wire415_out)
);
std_reg # (
    .WIDTH(1)
) cond416 (
    .clk(cond416_clk),
    .done(cond416_done),
    .in(cond416_in),
    .out(cond416_out),
    .reset(cond416_reset),
    .write_en(cond416_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire416 (
    .in(cond_wire416_in),
    .out(cond_wire416_out)
);
std_reg # (
    .WIDTH(1)
) cond417 (
    .clk(cond417_clk),
    .done(cond417_done),
    .in(cond417_in),
    .out(cond417_out),
    .reset(cond417_reset),
    .write_en(cond417_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire417 (
    .in(cond_wire417_in),
    .out(cond_wire417_out)
);
std_reg # (
    .WIDTH(1)
) cond418 (
    .clk(cond418_clk),
    .done(cond418_done),
    .in(cond418_in),
    .out(cond418_out),
    .reset(cond418_reset),
    .write_en(cond418_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire418 (
    .in(cond_wire418_in),
    .out(cond_wire418_out)
);
std_reg # (
    .WIDTH(1)
) cond419 (
    .clk(cond419_clk),
    .done(cond419_done),
    .in(cond419_in),
    .out(cond419_out),
    .reset(cond419_reset),
    .write_en(cond419_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire419 (
    .in(cond_wire419_in),
    .out(cond_wire419_out)
);
std_reg # (
    .WIDTH(1)
) cond420 (
    .clk(cond420_clk),
    .done(cond420_done),
    .in(cond420_in),
    .out(cond420_out),
    .reset(cond420_reset),
    .write_en(cond420_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire420 (
    .in(cond_wire420_in),
    .out(cond_wire420_out)
);
std_reg # (
    .WIDTH(1)
) cond421 (
    .clk(cond421_clk),
    .done(cond421_done),
    .in(cond421_in),
    .out(cond421_out),
    .reset(cond421_reset),
    .write_en(cond421_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire421 (
    .in(cond_wire421_in),
    .out(cond_wire421_out)
);
std_reg # (
    .WIDTH(1)
) cond422 (
    .clk(cond422_clk),
    .done(cond422_done),
    .in(cond422_in),
    .out(cond422_out),
    .reset(cond422_reset),
    .write_en(cond422_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire422 (
    .in(cond_wire422_in),
    .out(cond_wire422_out)
);
std_reg # (
    .WIDTH(1)
) cond423 (
    .clk(cond423_clk),
    .done(cond423_done),
    .in(cond423_in),
    .out(cond423_out),
    .reset(cond423_reset),
    .write_en(cond423_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire423 (
    .in(cond_wire423_in),
    .out(cond_wire423_out)
);
std_reg # (
    .WIDTH(1)
) cond424 (
    .clk(cond424_clk),
    .done(cond424_done),
    .in(cond424_in),
    .out(cond424_out),
    .reset(cond424_reset),
    .write_en(cond424_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire424 (
    .in(cond_wire424_in),
    .out(cond_wire424_out)
);
std_reg # (
    .WIDTH(1)
) cond425 (
    .clk(cond425_clk),
    .done(cond425_done),
    .in(cond425_in),
    .out(cond425_out),
    .reset(cond425_reset),
    .write_en(cond425_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire425 (
    .in(cond_wire425_in),
    .out(cond_wire425_out)
);
std_reg # (
    .WIDTH(1)
) cond426 (
    .clk(cond426_clk),
    .done(cond426_done),
    .in(cond426_in),
    .out(cond426_out),
    .reset(cond426_reset),
    .write_en(cond426_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire426 (
    .in(cond_wire426_in),
    .out(cond_wire426_out)
);
std_reg # (
    .WIDTH(1)
) cond427 (
    .clk(cond427_clk),
    .done(cond427_done),
    .in(cond427_in),
    .out(cond427_out),
    .reset(cond427_reset),
    .write_en(cond427_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire427 (
    .in(cond_wire427_in),
    .out(cond_wire427_out)
);
std_reg # (
    .WIDTH(1)
) cond428 (
    .clk(cond428_clk),
    .done(cond428_done),
    .in(cond428_in),
    .out(cond428_out),
    .reset(cond428_reset),
    .write_en(cond428_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire428 (
    .in(cond_wire428_in),
    .out(cond_wire428_out)
);
std_reg # (
    .WIDTH(1)
) cond429 (
    .clk(cond429_clk),
    .done(cond429_done),
    .in(cond429_in),
    .out(cond429_out),
    .reset(cond429_reset),
    .write_en(cond429_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire429 (
    .in(cond_wire429_in),
    .out(cond_wire429_out)
);
std_reg # (
    .WIDTH(1)
) cond430 (
    .clk(cond430_clk),
    .done(cond430_done),
    .in(cond430_in),
    .out(cond430_out),
    .reset(cond430_reset),
    .write_en(cond430_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire430 (
    .in(cond_wire430_in),
    .out(cond_wire430_out)
);
std_reg # (
    .WIDTH(1)
) cond431 (
    .clk(cond431_clk),
    .done(cond431_done),
    .in(cond431_in),
    .out(cond431_out),
    .reset(cond431_reset),
    .write_en(cond431_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire431 (
    .in(cond_wire431_in),
    .out(cond_wire431_out)
);
std_reg # (
    .WIDTH(1)
) cond432 (
    .clk(cond432_clk),
    .done(cond432_done),
    .in(cond432_in),
    .out(cond432_out),
    .reset(cond432_reset),
    .write_en(cond432_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire432 (
    .in(cond_wire432_in),
    .out(cond_wire432_out)
);
std_reg # (
    .WIDTH(1)
) cond433 (
    .clk(cond433_clk),
    .done(cond433_done),
    .in(cond433_in),
    .out(cond433_out),
    .reset(cond433_reset),
    .write_en(cond433_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire433 (
    .in(cond_wire433_in),
    .out(cond_wire433_out)
);
std_reg # (
    .WIDTH(1)
) cond434 (
    .clk(cond434_clk),
    .done(cond434_done),
    .in(cond434_in),
    .out(cond434_out),
    .reset(cond434_reset),
    .write_en(cond434_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire434 (
    .in(cond_wire434_in),
    .out(cond_wire434_out)
);
std_reg # (
    .WIDTH(1)
) cond435 (
    .clk(cond435_clk),
    .done(cond435_done),
    .in(cond435_in),
    .out(cond435_out),
    .reset(cond435_reset),
    .write_en(cond435_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire435 (
    .in(cond_wire435_in),
    .out(cond_wire435_out)
);
std_reg # (
    .WIDTH(1)
) cond436 (
    .clk(cond436_clk),
    .done(cond436_done),
    .in(cond436_in),
    .out(cond436_out),
    .reset(cond436_reset),
    .write_en(cond436_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire436 (
    .in(cond_wire436_in),
    .out(cond_wire436_out)
);
std_reg # (
    .WIDTH(1)
) cond437 (
    .clk(cond437_clk),
    .done(cond437_done),
    .in(cond437_in),
    .out(cond437_out),
    .reset(cond437_reset),
    .write_en(cond437_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire437 (
    .in(cond_wire437_in),
    .out(cond_wire437_out)
);
std_reg # (
    .WIDTH(1)
) cond438 (
    .clk(cond438_clk),
    .done(cond438_done),
    .in(cond438_in),
    .out(cond438_out),
    .reset(cond438_reset),
    .write_en(cond438_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire438 (
    .in(cond_wire438_in),
    .out(cond_wire438_out)
);
std_reg # (
    .WIDTH(1)
) cond439 (
    .clk(cond439_clk),
    .done(cond439_done),
    .in(cond439_in),
    .out(cond439_out),
    .reset(cond439_reset),
    .write_en(cond439_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire439 (
    .in(cond_wire439_in),
    .out(cond_wire439_out)
);
std_reg # (
    .WIDTH(1)
) cond440 (
    .clk(cond440_clk),
    .done(cond440_done),
    .in(cond440_in),
    .out(cond440_out),
    .reset(cond440_reset),
    .write_en(cond440_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire440 (
    .in(cond_wire440_in),
    .out(cond_wire440_out)
);
std_reg # (
    .WIDTH(1)
) cond441 (
    .clk(cond441_clk),
    .done(cond441_done),
    .in(cond441_in),
    .out(cond441_out),
    .reset(cond441_reset),
    .write_en(cond441_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire441 (
    .in(cond_wire441_in),
    .out(cond_wire441_out)
);
std_reg # (
    .WIDTH(1)
) cond442 (
    .clk(cond442_clk),
    .done(cond442_done),
    .in(cond442_in),
    .out(cond442_out),
    .reset(cond442_reset),
    .write_en(cond442_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire442 (
    .in(cond_wire442_in),
    .out(cond_wire442_out)
);
std_reg # (
    .WIDTH(1)
) cond443 (
    .clk(cond443_clk),
    .done(cond443_done),
    .in(cond443_in),
    .out(cond443_out),
    .reset(cond443_reset),
    .write_en(cond443_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire443 (
    .in(cond_wire443_in),
    .out(cond_wire443_out)
);
std_reg # (
    .WIDTH(1)
) cond444 (
    .clk(cond444_clk),
    .done(cond444_done),
    .in(cond444_in),
    .out(cond444_out),
    .reset(cond444_reset),
    .write_en(cond444_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire444 (
    .in(cond_wire444_in),
    .out(cond_wire444_out)
);
std_reg # (
    .WIDTH(1)
) cond445 (
    .clk(cond445_clk),
    .done(cond445_done),
    .in(cond445_in),
    .out(cond445_out),
    .reset(cond445_reset),
    .write_en(cond445_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire445 (
    .in(cond_wire445_in),
    .out(cond_wire445_out)
);
std_reg # (
    .WIDTH(1)
) cond446 (
    .clk(cond446_clk),
    .done(cond446_done),
    .in(cond446_in),
    .out(cond446_out),
    .reset(cond446_reset),
    .write_en(cond446_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire446 (
    .in(cond_wire446_in),
    .out(cond_wire446_out)
);
std_reg # (
    .WIDTH(1)
) cond447 (
    .clk(cond447_clk),
    .done(cond447_done),
    .in(cond447_in),
    .out(cond447_out),
    .reset(cond447_reset),
    .write_en(cond447_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire447 (
    .in(cond_wire447_in),
    .out(cond_wire447_out)
);
std_reg # (
    .WIDTH(1)
) cond448 (
    .clk(cond448_clk),
    .done(cond448_done),
    .in(cond448_in),
    .out(cond448_out),
    .reset(cond448_reset),
    .write_en(cond448_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire448 (
    .in(cond_wire448_in),
    .out(cond_wire448_out)
);
std_reg # (
    .WIDTH(1)
) cond449 (
    .clk(cond449_clk),
    .done(cond449_done),
    .in(cond449_in),
    .out(cond449_out),
    .reset(cond449_reset),
    .write_en(cond449_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire449 (
    .in(cond_wire449_in),
    .out(cond_wire449_out)
);
std_reg # (
    .WIDTH(1)
) cond450 (
    .clk(cond450_clk),
    .done(cond450_done),
    .in(cond450_in),
    .out(cond450_out),
    .reset(cond450_reset),
    .write_en(cond450_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire450 (
    .in(cond_wire450_in),
    .out(cond_wire450_out)
);
std_reg # (
    .WIDTH(1)
) cond451 (
    .clk(cond451_clk),
    .done(cond451_done),
    .in(cond451_in),
    .out(cond451_out),
    .reset(cond451_reset),
    .write_en(cond451_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire451 (
    .in(cond_wire451_in),
    .out(cond_wire451_out)
);
std_reg # (
    .WIDTH(1)
) cond452 (
    .clk(cond452_clk),
    .done(cond452_done),
    .in(cond452_in),
    .out(cond452_out),
    .reset(cond452_reset),
    .write_en(cond452_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire452 (
    .in(cond_wire452_in),
    .out(cond_wire452_out)
);
std_reg # (
    .WIDTH(1)
) cond453 (
    .clk(cond453_clk),
    .done(cond453_done),
    .in(cond453_in),
    .out(cond453_out),
    .reset(cond453_reset),
    .write_en(cond453_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire453 (
    .in(cond_wire453_in),
    .out(cond_wire453_out)
);
std_reg # (
    .WIDTH(1)
) cond454 (
    .clk(cond454_clk),
    .done(cond454_done),
    .in(cond454_in),
    .out(cond454_out),
    .reset(cond454_reset),
    .write_en(cond454_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire454 (
    .in(cond_wire454_in),
    .out(cond_wire454_out)
);
std_reg # (
    .WIDTH(1)
) cond455 (
    .clk(cond455_clk),
    .done(cond455_done),
    .in(cond455_in),
    .out(cond455_out),
    .reset(cond455_reset),
    .write_en(cond455_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire455 (
    .in(cond_wire455_in),
    .out(cond_wire455_out)
);
std_reg # (
    .WIDTH(1)
) cond456 (
    .clk(cond456_clk),
    .done(cond456_done),
    .in(cond456_in),
    .out(cond456_out),
    .reset(cond456_reset),
    .write_en(cond456_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire456 (
    .in(cond_wire456_in),
    .out(cond_wire456_out)
);
std_reg # (
    .WIDTH(1)
) cond457 (
    .clk(cond457_clk),
    .done(cond457_done),
    .in(cond457_in),
    .out(cond457_out),
    .reset(cond457_reset),
    .write_en(cond457_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire457 (
    .in(cond_wire457_in),
    .out(cond_wire457_out)
);
std_reg # (
    .WIDTH(1)
) cond458 (
    .clk(cond458_clk),
    .done(cond458_done),
    .in(cond458_in),
    .out(cond458_out),
    .reset(cond458_reset),
    .write_en(cond458_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire458 (
    .in(cond_wire458_in),
    .out(cond_wire458_out)
);
std_reg # (
    .WIDTH(1)
) cond459 (
    .clk(cond459_clk),
    .done(cond459_done),
    .in(cond459_in),
    .out(cond459_out),
    .reset(cond459_reset),
    .write_en(cond459_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire459 (
    .in(cond_wire459_in),
    .out(cond_wire459_out)
);
std_reg # (
    .WIDTH(1)
) cond460 (
    .clk(cond460_clk),
    .done(cond460_done),
    .in(cond460_in),
    .out(cond460_out),
    .reset(cond460_reset),
    .write_en(cond460_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire460 (
    .in(cond_wire460_in),
    .out(cond_wire460_out)
);
std_reg # (
    .WIDTH(1)
) cond461 (
    .clk(cond461_clk),
    .done(cond461_done),
    .in(cond461_in),
    .out(cond461_out),
    .reset(cond461_reset),
    .write_en(cond461_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire461 (
    .in(cond_wire461_in),
    .out(cond_wire461_out)
);
std_reg # (
    .WIDTH(1)
) cond462 (
    .clk(cond462_clk),
    .done(cond462_done),
    .in(cond462_in),
    .out(cond462_out),
    .reset(cond462_reset),
    .write_en(cond462_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire462 (
    .in(cond_wire462_in),
    .out(cond_wire462_out)
);
std_reg # (
    .WIDTH(1)
) cond463 (
    .clk(cond463_clk),
    .done(cond463_done),
    .in(cond463_in),
    .out(cond463_out),
    .reset(cond463_reset),
    .write_en(cond463_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire463 (
    .in(cond_wire463_in),
    .out(cond_wire463_out)
);
std_reg # (
    .WIDTH(1)
) cond464 (
    .clk(cond464_clk),
    .done(cond464_done),
    .in(cond464_in),
    .out(cond464_out),
    .reset(cond464_reset),
    .write_en(cond464_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire464 (
    .in(cond_wire464_in),
    .out(cond_wire464_out)
);
std_reg # (
    .WIDTH(1)
) cond465 (
    .clk(cond465_clk),
    .done(cond465_done),
    .in(cond465_in),
    .out(cond465_out),
    .reset(cond465_reset),
    .write_en(cond465_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire465 (
    .in(cond_wire465_in),
    .out(cond_wire465_out)
);
std_reg # (
    .WIDTH(1)
) cond466 (
    .clk(cond466_clk),
    .done(cond466_done),
    .in(cond466_in),
    .out(cond466_out),
    .reset(cond466_reset),
    .write_en(cond466_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire466 (
    .in(cond_wire466_in),
    .out(cond_wire466_out)
);
std_reg # (
    .WIDTH(1)
) cond467 (
    .clk(cond467_clk),
    .done(cond467_done),
    .in(cond467_in),
    .out(cond467_out),
    .reset(cond467_reset),
    .write_en(cond467_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire467 (
    .in(cond_wire467_in),
    .out(cond_wire467_out)
);
std_reg # (
    .WIDTH(1)
) cond468 (
    .clk(cond468_clk),
    .done(cond468_done),
    .in(cond468_in),
    .out(cond468_out),
    .reset(cond468_reset),
    .write_en(cond468_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire468 (
    .in(cond_wire468_in),
    .out(cond_wire468_out)
);
std_reg # (
    .WIDTH(1)
) cond469 (
    .clk(cond469_clk),
    .done(cond469_done),
    .in(cond469_in),
    .out(cond469_out),
    .reset(cond469_reset),
    .write_en(cond469_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire469 (
    .in(cond_wire469_in),
    .out(cond_wire469_out)
);
std_reg # (
    .WIDTH(1)
) cond470 (
    .clk(cond470_clk),
    .done(cond470_done),
    .in(cond470_in),
    .out(cond470_out),
    .reset(cond470_reset),
    .write_en(cond470_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire470 (
    .in(cond_wire470_in),
    .out(cond_wire470_out)
);
std_reg # (
    .WIDTH(1)
) cond471 (
    .clk(cond471_clk),
    .done(cond471_done),
    .in(cond471_in),
    .out(cond471_out),
    .reset(cond471_reset),
    .write_en(cond471_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire471 (
    .in(cond_wire471_in),
    .out(cond_wire471_out)
);
std_reg # (
    .WIDTH(1)
) cond472 (
    .clk(cond472_clk),
    .done(cond472_done),
    .in(cond472_in),
    .out(cond472_out),
    .reset(cond472_reset),
    .write_en(cond472_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire472 (
    .in(cond_wire472_in),
    .out(cond_wire472_out)
);
std_reg # (
    .WIDTH(1)
) cond473 (
    .clk(cond473_clk),
    .done(cond473_done),
    .in(cond473_in),
    .out(cond473_out),
    .reset(cond473_reset),
    .write_en(cond473_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire473 (
    .in(cond_wire473_in),
    .out(cond_wire473_out)
);
std_reg # (
    .WIDTH(1)
) cond474 (
    .clk(cond474_clk),
    .done(cond474_done),
    .in(cond474_in),
    .out(cond474_out),
    .reset(cond474_reset),
    .write_en(cond474_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire474 (
    .in(cond_wire474_in),
    .out(cond_wire474_out)
);
std_reg # (
    .WIDTH(1)
) cond475 (
    .clk(cond475_clk),
    .done(cond475_done),
    .in(cond475_in),
    .out(cond475_out),
    .reset(cond475_reset),
    .write_en(cond475_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire475 (
    .in(cond_wire475_in),
    .out(cond_wire475_out)
);
std_reg # (
    .WIDTH(1)
) cond476 (
    .clk(cond476_clk),
    .done(cond476_done),
    .in(cond476_in),
    .out(cond476_out),
    .reset(cond476_reset),
    .write_en(cond476_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire476 (
    .in(cond_wire476_in),
    .out(cond_wire476_out)
);
std_reg # (
    .WIDTH(1)
) cond477 (
    .clk(cond477_clk),
    .done(cond477_done),
    .in(cond477_in),
    .out(cond477_out),
    .reset(cond477_reset),
    .write_en(cond477_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire477 (
    .in(cond_wire477_in),
    .out(cond_wire477_out)
);
std_reg # (
    .WIDTH(1)
) cond478 (
    .clk(cond478_clk),
    .done(cond478_done),
    .in(cond478_in),
    .out(cond478_out),
    .reset(cond478_reset),
    .write_en(cond478_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire478 (
    .in(cond_wire478_in),
    .out(cond_wire478_out)
);
std_reg # (
    .WIDTH(1)
) cond479 (
    .clk(cond479_clk),
    .done(cond479_done),
    .in(cond479_in),
    .out(cond479_out),
    .reset(cond479_reset),
    .write_en(cond479_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire479 (
    .in(cond_wire479_in),
    .out(cond_wire479_out)
);
std_reg # (
    .WIDTH(1)
) cond480 (
    .clk(cond480_clk),
    .done(cond480_done),
    .in(cond480_in),
    .out(cond480_out),
    .reset(cond480_reset),
    .write_en(cond480_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire480 (
    .in(cond_wire480_in),
    .out(cond_wire480_out)
);
std_reg # (
    .WIDTH(1)
) cond481 (
    .clk(cond481_clk),
    .done(cond481_done),
    .in(cond481_in),
    .out(cond481_out),
    .reset(cond481_reset),
    .write_en(cond481_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire481 (
    .in(cond_wire481_in),
    .out(cond_wire481_out)
);
std_reg # (
    .WIDTH(1)
) cond482 (
    .clk(cond482_clk),
    .done(cond482_done),
    .in(cond482_in),
    .out(cond482_out),
    .reset(cond482_reset),
    .write_en(cond482_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire482 (
    .in(cond_wire482_in),
    .out(cond_wire482_out)
);
std_reg # (
    .WIDTH(1)
) cond483 (
    .clk(cond483_clk),
    .done(cond483_done),
    .in(cond483_in),
    .out(cond483_out),
    .reset(cond483_reset),
    .write_en(cond483_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire483 (
    .in(cond_wire483_in),
    .out(cond_wire483_out)
);
std_reg # (
    .WIDTH(1)
) cond484 (
    .clk(cond484_clk),
    .done(cond484_done),
    .in(cond484_in),
    .out(cond484_out),
    .reset(cond484_reset),
    .write_en(cond484_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire484 (
    .in(cond_wire484_in),
    .out(cond_wire484_out)
);
std_reg # (
    .WIDTH(1)
) cond485 (
    .clk(cond485_clk),
    .done(cond485_done),
    .in(cond485_in),
    .out(cond485_out),
    .reset(cond485_reset),
    .write_en(cond485_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire485 (
    .in(cond_wire485_in),
    .out(cond_wire485_out)
);
std_reg # (
    .WIDTH(1)
) cond486 (
    .clk(cond486_clk),
    .done(cond486_done),
    .in(cond486_in),
    .out(cond486_out),
    .reset(cond486_reset),
    .write_en(cond486_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire486 (
    .in(cond_wire486_in),
    .out(cond_wire486_out)
);
std_reg # (
    .WIDTH(1)
) cond487 (
    .clk(cond487_clk),
    .done(cond487_done),
    .in(cond487_in),
    .out(cond487_out),
    .reset(cond487_reset),
    .write_en(cond487_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire487 (
    .in(cond_wire487_in),
    .out(cond_wire487_out)
);
std_reg # (
    .WIDTH(1)
) cond488 (
    .clk(cond488_clk),
    .done(cond488_done),
    .in(cond488_in),
    .out(cond488_out),
    .reset(cond488_reset),
    .write_en(cond488_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire488 (
    .in(cond_wire488_in),
    .out(cond_wire488_out)
);
std_reg # (
    .WIDTH(1)
) cond489 (
    .clk(cond489_clk),
    .done(cond489_done),
    .in(cond489_in),
    .out(cond489_out),
    .reset(cond489_reset),
    .write_en(cond489_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire489 (
    .in(cond_wire489_in),
    .out(cond_wire489_out)
);
std_reg # (
    .WIDTH(1)
) cond490 (
    .clk(cond490_clk),
    .done(cond490_done),
    .in(cond490_in),
    .out(cond490_out),
    .reset(cond490_reset),
    .write_en(cond490_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire490 (
    .in(cond_wire490_in),
    .out(cond_wire490_out)
);
std_reg # (
    .WIDTH(1)
) cond491 (
    .clk(cond491_clk),
    .done(cond491_done),
    .in(cond491_in),
    .out(cond491_out),
    .reset(cond491_reset),
    .write_en(cond491_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire491 (
    .in(cond_wire491_in),
    .out(cond_wire491_out)
);
std_reg # (
    .WIDTH(1)
) cond492 (
    .clk(cond492_clk),
    .done(cond492_done),
    .in(cond492_in),
    .out(cond492_out),
    .reset(cond492_reset),
    .write_en(cond492_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire492 (
    .in(cond_wire492_in),
    .out(cond_wire492_out)
);
std_reg # (
    .WIDTH(1)
) cond493 (
    .clk(cond493_clk),
    .done(cond493_done),
    .in(cond493_in),
    .out(cond493_out),
    .reset(cond493_reset),
    .write_en(cond493_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire493 (
    .in(cond_wire493_in),
    .out(cond_wire493_out)
);
std_reg # (
    .WIDTH(1)
) cond494 (
    .clk(cond494_clk),
    .done(cond494_done),
    .in(cond494_in),
    .out(cond494_out),
    .reset(cond494_reset),
    .write_en(cond494_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire494 (
    .in(cond_wire494_in),
    .out(cond_wire494_out)
);
std_reg # (
    .WIDTH(1)
) cond495 (
    .clk(cond495_clk),
    .done(cond495_done),
    .in(cond495_in),
    .out(cond495_out),
    .reset(cond495_reset),
    .write_en(cond495_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire495 (
    .in(cond_wire495_in),
    .out(cond_wire495_out)
);
std_reg # (
    .WIDTH(1)
) cond496 (
    .clk(cond496_clk),
    .done(cond496_done),
    .in(cond496_in),
    .out(cond496_out),
    .reset(cond496_reset),
    .write_en(cond496_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire496 (
    .in(cond_wire496_in),
    .out(cond_wire496_out)
);
std_reg # (
    .WIDTH(1)
) cond497 (
    .clk(cond497_clk),
    .done(cond497_done),
    .in(cond497_in),
    .out(cond497_out),
    .reset(cond497_reset),
    .write_en(cond497_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire497 (
    .in(cond_wire497_in),
    .out(cond_wire497_out)
);
std_reg # (
    .WIDTH(1)
) cond498 (
    .clk(cond498_clk),
    .done(cond498_done),
    .in(cond498_in),
    .out(cond498_out),
    .reset(cond498_reset),
    .write_en(cond498_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire498 (
    .in(cond_wire498_in),
    .out(cond_wire498_out)
);
std_reg # (
    .WIDTH(1)
) cond499 (
    .clk(cond499_clk),
    .done(cond499_done),
    .in(cond499_in),
    .out(cond499_out),
    .reset(cond499_reset),
    .write_en(cond499_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire499 (
    .in(cond_wire499_in),
    .out(cond_wire499_out)
);
std_reg # (
    .WIDTH(1)
) cond500 (
    .clk(cond500_clk),
    .done(cond500_done),
    .in(cond500_in),
    .out(cond500_out),
    .reset(cond500_reset),
    .write_en(cond500_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire500 (
    .in(cond_wire500_in),
    .out(cond_wire500_out)
);
std_reg # (
    .WIDTH(1)
) cond501 (
    .clk(cond501_clk),
    .done(cond501_done),
    .in(cond501_in),
    .out(cond501_out),
    .reset(cond501_reset),
    .write_en(cond501_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire501 (
    .in(cond_wire501_in),
    .out(cond_wire501_out)
);
std_reg # (
    .WIDTH(1)
) cond502 (
    .clk(cond502_clk),
    .done(cond502_done),
    .in(cond502_in),
    .out(cond502_out),
    .reset(cond502_reset),
    .write_en(cond502_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire502 (
    .in(cond_wire502_in),
    .out(cond_wire502_out)
);
std_reg # (
    .WIDTH(1)
) cond503 (
    .clk(cond503_clk),
    .done(cond503_done),
    .in(cond503_in),
    .out(cond503_out),
    .reset(cond503_reset),
    .write_en(cond503_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire503 (
    .in(cond_wire503_in),
    .out(cond_wire503_out)
);
std_reg # (
    .WIDTH(1)
) cond504 (
    .clk(cond504_clk),
    .done(cond504_done),
    .in(cond504_in),
    .out(cond504_out),
    .reset(cond504_reset),
    .write_en(cond504_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire504 (
    .in(cond_wire504_in),
    .out(cond_wire504_out)
);
std_reg # (
    .WIDTH(1)
) cond505 (
    .clk(cond505_clk),
    .done(cond505_done),
    .in(cond505_in),
    .out(cond505_out),
    .reset(cond505_reset),
    .write_en(cond505_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire505 (
    .in(cond_wire505_in),
    .out(cond_wire505_out)
);
std_reg # (
    .WIDTH(1)
) cond506 (
    .clk(cond506_clk),
    .done(cond506_done),
    .in(cond506_in),
    .out(cond506_out),
    .reset(cond506_reset),
    .write_en(cond506_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire506 (
    .in(cond_wire506_in),
    .out(cond_wire506_out)
);
std_reg # (
    .WIDTH(1)
) cond507 (
    .clk(cond507_clk),
    .done(cond507_done),
    .in(cond507_in),
    .out(cond507_out),
    .reset(cond507_reset),
    .write_en(cond507_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire507 (
    .in(cond_wire507_in),
    .out(cond_wire507_out)
);
std_reg # (
    .WIDTH(1)
) cond508 (
    .clk(cond508_clk),
    .done(cond508_done),
    .in(cond508_in),
    .out(cond508_out),
    .reset(cond508_reset),
    .write_en(cond508_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire508 (
    .in(cond_wire508_in),
    .out(cond_wire508_out)
);
std_reg # (
    .WIDTH(1)
) cond509 (
    .clk(cond509_clk),
    .done(cond509_done),
    .in(cond509_in),
    .out(cond509_out),
    .reset(cond509_reset),
    .write_en(cond509_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire509 (
    .in(cond_wire509_in),
    .out(cond_wire509_out)
);
std_reg # (
    .WIDTH(1)
) cond510 (
    .clk(cond510_clk),
    .done(cond510_done),
    .in(cond510_in),
    .out(cond510_out),
    .reset(cond510_reset),
    .write_en(cond510_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire510 (
    .in(cond_wire510_in),
    .out(cond_wire510_out)
);
std_reg # (
    .WIDTH(1)
) cond511 (
    .clk(cond511_clk),
    .done(cond511_done),
    .in(cond511_in),
    .out(cond511_out),
    .reset(cond511_reset),
    .write_en(cond511_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire511 (
    .in(cond_wire511_in),
    .out(cond_wire511_out)
);
std_reg # (
    .WIDTH(1)
) cond512 (
    .clk(cond512_clk),
    .done(cond512_done),
    .in(cond512_in),
    .out(cond512_out),
    .reset(cond512_reset),
    .write_en(cond512_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire512 (
    .in(cond_wire512_in),
    .out(cond_wire512_out)
);
std_reg # (
    .WIDTH(1)
) cond513 (
    .clk(cond513_clk),
    .done(cond513_done),
    .in(cond513_in),
    .out(cond513_out),
    .reset(cond513_reset),
    .write_en(cond513_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire513 (
    .in(cond_wire513_in),
    .out(cond_wire513_out)
);
std_reg # (
    .WIDTH(1)
) cond514 (
    .clk(cond514_clk),
    .done(cond514_done),
    .in(cond514_in),
    .out(cond514_out),
    .reset(cond514_reset),
    .write_en(cond514_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire514 (
    .in(cond_wire514_in),
    .out(cond_wire514_out)
);
std_reg # (
    .WIDTH(1)
) cond515 (
    .clk(cond515_clk),
    .done(cond515_done),
    .in(cond515_in),
    .out(cond515_out),
    .reset(cond515_reset),
    .write_en(cond515_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire515 (
    .in(cond_wire515_in),
    .out(cond_wire515_out)
);
std_reg # (
    .WIDTH(1)
) cond516 (
    .clk(cond516_clk),
    .done(cond516_done),
    .in(cond516_in),
    .out(cond516_out),
    .reset(cond516_reset),
    .write_en(cond516_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire516 (
    .in(cond_wire516_in),
    .out(cond_wire516_out)
);
std_reg # (
    .WIDTH(1)
) cond517 (
    .clk(cond517_clk),
    .done(cond517_done),
    .in(cond517_in),
    .out(cond517_out),
    .reset(cond517_reset),
    .write_en(cond517_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire517 (
    .in(cond_wire517_in),
    .out(cond_wire517_out)
);
std_reg # (
    .WIDTH(1)
) cond518 (
    .clk(cond518_clk),
    .done(cond518_done),
    .in(cond518_in),
    .out(cond518_out),
    .reset(cond518_reset),
    .write_en(cond518_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire518 (
    .in(cond_wire518_in),
    .out(cond_wire518_out)
);
std_reg # (
    .WIDTH(1)
) cond519 (
    .clk(cond519_clk),
    .done(cond519_done),
    .in(cond519_in),
    .out(cond519_out),
    .reset(cond519_reset),
    .write_en(cond519_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire519 (
    .in(cond_wire519_in),
    .out(cond_wire519_out)
);
std_reg # (
    .WIDTH(1)
) cond520 (
    .clk(cond520_clk),
    .done(cond520_done),
    .in(cond520_in),
    .out(cond520_out),
    .reset(cond520_reset),
    .write_en(cond520_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire520 (
    .in(cond_wire520_in),
    .out(cond_wire520_out)
);
std_reg # (
    .WIDTH(1)
) cond521 (
    .clk(cond521_clk),
    .done(cond521_done),
    .in(cond521_in),
    .out(cond521_out),
    .reset(cond521_reset),
    .write_en(cond521_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire521 (
    .in(cond_wire521_in),
    .out(cond_wire521_out)
);
std_reg # (
    .WIDTH(1)
) cond522 (
    .clk(cond522_clk),
    .done(cond522_done),
    .in(cond522_in),
    .out(cond522_out),
    .reset(cond522_reset),
    .write_en(cond522_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire522 (
    .in(cond_wire522_in),
    .out(cond_wire522_out)
);
std_reg # (
    .WIDTH(1)
) cond523 (
    .clk(cond523_clk),
    .done(cond523_done),
    .in(cond523_in),
    .out(cond523_out),
    .reset(cond523_reset),
    .write_en(cond523_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire523 (
    .in(cond_wire523_in),
    .out(cond_wire523_out)
);
std_reg # (
    .WIDTH(1)
) cond524 (
    .clk(cond524_clk),
    .done(cond524_done),
    .in(cond524_in),
    .out(cond524_out),
    .reset(cond524_reset),
    .write_en(cond524_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire524 (
    .in(cond_wire524_in),
    .out(cond_wire524_out)
);
std_reg # (
    .WIDTH(1)
) cond525 (
    .clk(cond525_clk),
    .done(cond525_done),
    .in(cond525_in),
    .out(cond525_out),
    .reset(cond525_reset),
    .write_en(cond525_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire525 (
    .in(cond_wire525_in),
    .out(cond_wire525_out)
);
std_reg # (
    .WIDTH(1)
) cond526 (
    .clk(cond526_clk),
    .done(cond526_done),
    .in(cond526_in),
    .out(cond526_out),
    .reset(cond526_reset),
    .write_en(cond526_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire526 (
    .in(cond_wire526_in),
    .out(cond_wire526_out)
);
std_reg # (
    .WIDTH(1)
) cond527 (
    .clk(cond527_clk),
    .done(cond527_done),
    .in(cond527_in),
    .out(cond527_out),
    .reset(cond527_reset),
    .write_en(cond527_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire527 (
    .in(cond_wire527_in),
    .out(cond_wire527_out)
);
std_reg # (
    .WIDTH(1)
) cond528 (
    .clk(cond528_clk),
    .done(cond528_done),
    .in(cond528_in),
    .out(cond528_out),
    .reset(cond528_reset),
    .write_en(cond528_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire528 (
    .in(cond_wire528_in),
    .out(cond_wire528_out)
);
std_reg # (
    .WIDTH(1)
) cond529 (
    .clk(cond529_clk),
    .done(cond529_done),
    .in(cond529_in),
    .out(cond529_out),
    .reset(cond529_reset),
    .write_en(cond529_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire529 (
    .in(cond_wire529_in),
    .out(cond_wire529_out)
);
std_reg # (
    .WIDTH(1)
) cond530 (
    .clk(cond530_clk),
    .done(cond530_done),
    .in(cond530_in),
    .out(cond530_out),
    .reset(cond530_reset),
    .write_en(cond530_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire530 (
    .in(cond_wire530_in),
    .out(cond_wire530_out)
);
std_reg # (
    .WIDTH(1)
) cond531 (
    .clk(cond531_clk),
    .done(cond531_done),
    .in(cond531_in),
    .out(cond531_out),
    .reset(cond531_reset),
    .write_en(cond531_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire531 (
    .in(cond_wire531_in),
    .out(cond_wire531_out)
);
std_reg # (
    .WIDTH(1)
) cond532 (
    .clk(cond532_clk),
    .done(cond532_done),
    .in(cond532_in),
    .out(cond532_out),
    .reset(cond532_reset),
    .write_en(cond532_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire532 (
    .in(cond_wire532_in),
    .out(cond_wire532_out)
);
std_reg # (
    .WIDTH(1)
) cond533 (
    .clk(cond533_clk),
    .done(cond533_done),
    .in(cond533_in),
    .out(cond533_out),
    .reset(cond533_reset),
    .write_en(cond533_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire533 (
    .in(cond_wire533_in),
    .out(cond_wire533_out)
);
std_reg # (
    .WIDTH(1)
) cond534 (
    .clk(cond534_clk),
    .done(cond534_done),
    .in(cond534_in),
    .out(cond534_out),
    .reset(cond534_reset),
    .write_en(cond534_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire534 (
    .in(cond_wire534_in),
    .out(cond_wire534_out)
);
std_reg # (
    .WIDTH(1)
) cond535 (
    .clk(cond535_clk),
    .done(cond535_done),
    .in(cond535_in),
    .out(cond535_out),
    .reset(cond535_reset),
    .write_en(cond535_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire535 (
    .in(cond_wire535_in),
    .out(cond_wire535_out)
);
std_reg # (
    .WIDTH(1)
) cond536 (
    .clk(cond536_clk),
    .done(cond536_done),
    .in(cond536_in),
    .out(cond536_out),
    .reset(cond536_reset),
    .write_en(cond536_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire536 (
    .in(cond_wire536_in),
    .out(cond_wire536_out)
);
std_reg # (
    .WIDTH(1)
) cond537 (
    .clk(cond537_clk),
    .done(cond537_done),
    .in(cond537_in),
    .out(cond537_out),
    .reset(cond537_reset),
    .write_en(cond537_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire537 (
    .in(cond_wire537_in),
    .out(cond_wire537_out)
);
std_reg # (
    .WIDTH(1)
) cond538 (
    .clk(cond538_clk),
    .done(cond538_done),
    .in(cond538_in),
    .out(cond538_out),
    .reset(cond538_reset),
    .write_en(cond538_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire538 (
    .in(cond_wire538_in),
    .out(cond_wire538_out)
);
std_reg # (
    .WIDTH(1)
) cond539 (
    .clk(cond539_clk),
    .done(cond539_done),
    .in(cond539_in),
    .out(cond539_out),
    .reset(cond539_reset),
    .write_en(cond539_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire539 (
    .in(cond_wire539_in),
    .out(cond_wire539_out)
);
std_reg # (
    .WIDTH(1)
) cond540 (
    .clk(cond540_clk),
    .done(cond540_done),
    .in(cond540_in),
    .out(cond540_out),
    .reset(cond540_reset),
    .write_en(cond540_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire540 (
    .in(cond_wire540_in),
    .out(cond_wire540_out)
);
std_reg # (
    .WIDTH(1)
) cond541 (
    .clk(cond541_clk),
    .done(cond541_done),
    .in(cond541_in),
    .out(cond541_out),
    .reset(cond541_reset),
    .write_en(cond541_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire541 (
    .in(cond_wire541_in),
    .out(cond_wire541_out)
);
std_reg # (
    .WIDTH(1)
) cond542 (
    .clk(cond542_clk),
    .done(cond542_done),
    .in(cond542_in),
    .out(cond542_out),
    .reset(cond542_reset),
    .write_en(cond542_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire542 (
    .in(cond_wire542_in),
    .out(cond_wire542_out)
);
std_reg # (
    .WIDTH(1)
) cond543 (
    .clk(cond543_clk),
    .done(cond543_done),
    .in(cond543_in),
    .out(cond543_out),
    .reset(cond543_reset),
    .write_en(cond543_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire543 (
    .in(cond_wire543_in),
    .out(cond_wire543_out)
);
std_reg # (
    .WIDTH(1)
) cond544 (
    .clk(cond544_clk),
    .done(cond544_done),
    .in(cond544_in),
    .out(cond544_out),
    .reset(cond544_reset),
    .write_en(cond544_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire544 (
    .in(cond_wire544_in),
    .out(cond_wire544_out)
);
std_reg # (
    .WIDTH(1)
) cond545 (
    .clk(cond545_clk),
    .done(cond545_done),
    .in(cond545_in),
    .out(cond545_out),
    .reset(cond545_reset),
    .write_en(cond545_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire545 (
    .in(cond_wire545_in),
    .out(cond_wire545_out)
);
std_reg # (
    .WIDTH(1)
) cond546 (
    .clk(cond546_clk),
    .done(cond546_done),
    .in(cond546_in),
    .out(cond546_out),
    .reset(cond546_reset),
    .write_en(cond546_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire546 (
    .in(cond_wire546_in),
    .out(cond_wire546_out)
);
std_reg # (
    .WIDTH(1)
) cond547 (
    .clk(cond547_clk),
    .done(cond547_done),
    .in(cond547_in),
    .out(cond547_out),
    .reset(cond547_reset),
    .write_en(cond547_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire547 (
    .in(cond_wire547_in),
    .out(cond_wire547_out)
);
std_reg # (
    .WIDTH(1)
) cond548 (
    .clk(cond548_clk),
    .done(cond548_done),
    .in(cond548_in),
    .out(cond548_out),
    .reset(cond548_reset),
    .write_en(cond548_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire548 (
    .in(cond_wire548_in),
    .out(cond_wire548_out)
);
std_reg # (
    .WIDTH(1)
) cond549 (
    .clk(cond549_clk),
    .done(cond549_done),
    .in(cond549_in),
    .out(cond549_out),
    .reset(cond549_reset),
    .write_en(cond549_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire549 (
    .in(cond_wire549_in),
    .out(cond_wire549_out)
);
std_reg # (
    .WIDTH(1)
) cond550 (
    .clk(cond550_clk),
    .done(cond550_done),
    .in(cond550_in),
    .out(cond550_out),
    .reset(cond550_reset),
    .write_en(cond550_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire550 (
    .in(cond_wire550_in),
    .out(cond_wire550_out)
);
std_reg # (
    .WIDTH(1)
) cond551 (
    .clk(cond551_clk),
    .done(cond551_done),
    .in(cond551_in),
    .out(cond551_out),
    .reset(cond551_reset),
    .write_en(cond551_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire551 (
    .in(cond_wire551_in),
    .out(cond_wire551_out)
);
std_reg # (
    .WIDTH(1)
) cond552 (
    .clk(cond552_clk),
    .done(cond552_done),
    .in(cond552_in),
    .out(cond552_out),
    .reset(cond552_reset),
    .write_en(cond552_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire552 (
    .in(cond_wire552_in),
    .out(cond_wire552_out)
);
std_reg # (
    .WIDTH(1)
) cond553 (
    .clk(cond553_clk),
    .done(cond553_done),
    .in(cond553_in),
    .out(cond553_out),
    .reset(cond553_reset),
    .write_en(cond553_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire553 (
    .in(cond_wire553_in),
    .out(cond_wire553_out)
);
std_reg # (
    .WIDTH(1)
) cond554 (
    .clk(cond554_clk),
    .done(cond554_done),
    .in(cond554_in),
    .out(cond554_out),
    .reset(cond554_reset),
    .write_en(cond554_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire554 (
    .in(cond_wire554_in),
    .out(cond_wire554_out)
);
std_reg # (
    .WIDTH(1)
) cond555 (
    .clk(cond555_clk),
    .done(cond555_done),
    .in(cond555_in),
    .out(cond555_out),
    .reset(cond555_reset),
    .write_en(cond555_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire555 (
    .in(cond_wire555_in),
    .out(cond_wire555_out)
);
std_reg # (
    .WIDTH(1)
) cond556 (
    .clk(cond556_clk),
    .done(cond556_done),
    .in(cond556_in),
    .out(cond556_out),
    .reset(cond556_reset),
    .write_en(cond556_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire556 (
    .in(cond_wire556_in),
    .out(cond_wire556_out)
);
std_reg # (
    .WIDTH(1)
) cond557 (
    .clk(cond557_clk),
    .done(cond557_done),
    .in(cond557_in),
    .out(cond557_out),
    .reset(cond557_reset),
    .write_en(cond557_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire557 (
    .in(cond_wire557_in),
    .out(cond_wire557_out)
);
std_reg # (
    .WIDTH(1)
) cond558 (
    .clk(cond558_clk),
    .done(cond558_done),
    .in(cond558_in),
    .out(cond558_out),
    .reset(cond558_reset),
    .write_en(cond558_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire558 (
    .in(cond_wire558_in),
    .out(cond_wire558_out)
);
std_reg # (
    .WIDTH(1)
) cond559 (
    .clk(cond559_clk),
    .done(cond559_done),
    .in(cond559_in),
    .out(cond559_out),
    .reset(cond559_reset),
    .write_en(cond559_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire559 (
    .in(cond_wire559_in),
    .out(cond_wire559_out)
);
std_reg # (
    .WIDTH(1)
) cond560 (
    .clk(cond560_clk),
    .done(cond560_done),
    .in(cond560_in),
    .out(cond560_out),
    .reset(cond560_reset),
    .write_en(cond560_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire560 (
    .in(cond_wire560_in),
    .out(cond_wire560_out)
);
std_reg # (
    .WIDTH(1)
) cond561 (
    .clk(cond561_clk),
    .done(cond561_done),
    .in(cond561_in),
    .out(cond561_out),
    .reset(cond561_reset),
    .write_en(cond561_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire561 (
    .in(cond_wire561_in),
    .out(cond_wire561_out)
);
std_reg # (
    .WIDTH(1)
) cond562 (
    .clk(cond562_clk),
    .done(cond562_done),
    .in(cond562_in),
    .out(cond562_out),
    .reset(cond562_reset),
    .write_en(cond562_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire562 (
    .in(cond_wire562_in),
    .out(cond_wire562_out)
);
std_reg # (
    .WIDTH(1)
) cond563 (
    .clk(cond563_clk),
    .done(cond563_done),
    .in(cond563_in),
    .out(cond563_out),
    .reset(cond563_reset),
    .write_en(cond563_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire563 (
    .in(cond_wire563_in),
    .out(cond_wire563_out)
);
std_reg # (
    .WIDTH(1)
) cond564 (
    .clk(cond564_clk),
    .done(cond564_done),
    .in(cond564_in),
    .out(cond564_out),
    .reset(cond564_reset),
    .write_en(cond564_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire564 (
    .in(cond_wire564_in),
    .out(cond_wire564_out)
);
std_reg # (
    .WIDTH(1)
) cond565 (
    .clk(cond565_clk),
    .done(cond565_done),
    .in(cond565_in),
    .out(cond565_out),
    .reset(cond565_reset),
    .write_en(cond565_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire565 (
    .in(cond_wire565_in),
    .out(cond_wire565_out)
);
std_reg # (
    .WIDTH(1)
) cond566 (
    .clk(cond566_clk),
    .done(cond566_done),
    .in(cond566_in),
    .out(cond566_out),
    .reset(cond566_reset),
    .write_en(cond566_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire566 (
    .in(cond_wire566_in),
    .out(cond_wire566_out)
);
std_reg # (
    .WIDTH(1)
) cond567 (
    .clk(cond567_clk),
    .done(cond567_done),
    .in(cond567_in),
    .out(cond567_out),
    .reset(cond567_reset),
    .write_en(cond567_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire567 (
    .in(cond_wire567_in),
    .out(cond_wire567_out)
);
std_reg # (
    .WIDTH(1)
) cond568 (
    .clk(cond568_clk),
    .done(cond568_done),
    .in(cond568_in),
    .out(cond568_out),
    .reset(cond568_reset),
    .write_en(cond568_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire568 (
    .in(cond_wire568_in),
    .out(cond_wire568_out)
);
std_reg # (
    .WIDTH(1)
) cond569 (
    .clk(cond569_clk),
    .done(cond569_done),
    .in(cond569_in),
    .out(cond569_out),
    .reset(cond569_reset),
    .write_en(cond569_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire569 (
    .in(cond_wire569_in),
    .out(cond_wire569_out)
);
std_reg # (
    .WIDTH(1)
) cond570 (
    .clk(cond570_clk),
    .done(cond570_done),
    .in(cond570_in),
    .out(cond570_out),
    .reset(cond570_reset),
    .write_en(cond570_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire570 (
    .in(cond_wire570_in),
    .out(cond_wire570_out)
);
std_reg # (
    .WIDTH(1)
) cond571 (
    .clk(cond571_clk),
    .done(cond571_done),
    .in(cond571_in),
    .out(cond571_out),
    .reset(cond571_reset),
    .write_en(cond571_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire571 (
    .in(cond_wire571_in),
    .out(cond_wire571_out)
);
std_reg # (
    .WIDTH(1)
) cond572 (
    .clk(cond572_clk),
    .done(cond572_done),
    .in(cond572_in),
    .out(cond572_out),
    .reset(cond572_reset),
    .write_en(cond572_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire572 (
    .in(cond_wire572_in),
    .out(cond_wire572_out)
);
std_reg # (
    .WIDTH(1)
) cond573 (
    .clk(cond573_clk),
    .done(cond573_done),
    .in(cond573_in),
    .out(cond573_out),
    .reset(cond573_reset),
    .write_en(cond573_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire573 (
    .in(cond_wire573_in),
    .out(cond_wire573_out)
);
std_reg # (
    .WIDTH(1)
) cond574 (
    .clk(cond574_clk),
    .done(cond574_done),
    .in(cond574_in),
    .out(cond574_out),
    .reset(cond574_reset),
    .write_en(cond574_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire574 (
    .in(cond_wire574_in),
    .out(cond_wire574_out)
);
std_reg # (
    .WIDTH(1)
) cond575 (
    .clk(cond575_clk),
    .done(cond575_done),
    .in(cond575_in),
    .out(cond575_out),
    .reset(cond575_reset),
    .write_en(cond575_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire575 (
    .in(cond_wire575_in),
    .out(cond_wire575_out)
);
std_reg # (
    .WIDTH(1)
) cond576 (
    .clk(cond576_clk),
    .done(cond576_done),
    .in(cond576_in),
    .out(cond576_out),
    .reset(cond576_reset),
    .write_en(cond576_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire576 (
    .in(cond_wire576_in),
    .out(cond_wire576_out)
);
std_reg # (
    .WIDTH(1)
) cond577 (
    .clk(cond577_clk),
    .done(cond577_done),
    .in(cond577_in),
    .out(cond577_out),
    .reset(cond577_reset),
    .write_en(cond577_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire577 (
    .in(cond_wire577_in),
    .out(cond_wire577_out)
);
std_reg # (
    .WIDTH(1)
) cond578 (
    .clk(cond578_clk),
    .done(cond578_done),
    .in(cond578_in),
    .out(cond578_out),
    .reset(cond578_reset),
    .write_en(cond578_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire578 (
    .in(cond_wire578_in),
    .out(cond_wire578_out)
);
std_reg # (
    .WIDTH(1)
) cond579 (
    .clk(cond579_clk),
    .done(cond579_done),
    .in(cond579_in),
    .out(cond579_out),
    .reset(cond579_reset),
    .write_en(cond579_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire579 (
    .in(cond_wire579_in),
    .out(cond_wire579_out)
);
std_reg # (
    .WIDTH(1)
) cond580 (
    .clk(cond580_clk),
    .done(cond580_done),
    .in(cond580_in),
    .out(cond580_out),
    .reset(cond580_reset),
    .write_en(cond580_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire580 (
    .in(cond_wire580_in),
    .out(cond_wire580_out)
);
std_reg # (
    .WIDTH(1)
) cond581 (
    .clk(cond581_clk),
    .done(cond581_done),
    .in(cond581_in),
    .out(cond581_out),
    .reset(cond581_reset),
    .write_en(cond581_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire581 (
    .in(cond_wire581_in),
    .out(cond_wire581_out)
);
std_reg # (
    .WIDTH(1)
) cond582 (
    .clk(cond582_clk),
    .done(cond582_done),
    .in(cond582_in),
    .out(cond582_out),
    .reset(cond582_reset),
    .write_en(cond582_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire582 (
    .in(cond_wire582_in),
    .out(cond_wire582_out)
);
std_reg # (
    .WIDTH(1)
) cond583 (
    .clk(cond583_clk),
    .done(cond583_done),
    .in(cond583_in),
    .out(cond583_out),
    .reset(cond583_reset),
    .write_en(cond583_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire583 (
    .in(cond_wire583_in),
    .out(cond_wire583_out)
);
std_reg # (
    .WIDTH(1)
) cond584 (
    .clk(cond584_clk),
    .done(cond584_done),
    .in(cond584_in),
    .out(cond584_out),
    .reset(cond584_reset),
    .write_en(cond584_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire584 (
    .in(cond_wire584_in),
    .out(cond_wire584_out)
);
std_reg # (
    .WIDTH(1)
) cond585 (
    .clk(cond585_clk),
    .done(cond585_done),
    .in(cond585_in),
    .out(cond585_out),
    .reset(cond585_reset),
    .write_en(cond585_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire585 (
    .in(cond_wire585_in),
    .out(cond_wire585_out)
);
std_reg # (
    .WIDTH(1)
) cond586 (
    .clk(cond586_clk),
    .done(cond586_done),
    .in(cond586_in),
    .out(cond586_out),
    .reset(cond586_reset),
    .write_en(cond586_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire586 (
    .in(cond_wire586_in),
    .out(cond_wire586_out)
);
std_reg # (
    .WIDTH(1)
) cond587 (
    .clk(cond587_clk),
    .done(cond587_done),
    .in(cond587_in),
    .out(cond587_out),
    .reset(cond587_reset),
    .write_en(cond587_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire587 (
    .in(cond_wire587_in),
    .out(cond_wire587_out)
);
std_reg # (
    .WIDTH(1)
) cond588 (
    .clk(cond588_clk),
    .done(cond588_done),
    .in(cond588_in),
    .out(cond588_out),
    .reset(cond588_reset),
    .write_en(cond588_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire588 (
    .in(cond_wire588_in),
    .out(cond_wire588_out)
);
std_reg # (
    .WIDTH(1)
) cond589 (
    .clk(cond589_clk),
    .done(cond589_done),
    .in(cond589_in),
    .out(cond589_out),
    .reset(cond589_reset),
    .write_en(cond589_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire589 (
    .in(cond_wire589_in),
    .out(cond_wire589_out)
);
std_reg # (
    .WIDTH(1)
) cond590 (
    .clk(cond590_clk),
    .done(cond590_done),
    .in(cond590_in),
    .out(cond590_out),
    .reset(cond590_reset),
    .write_en(cond590_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire590 (
    .in(cond_wire590_in),
    .out(cond_wire590_out)
);
std_reg # (
    .WIDTH(1)
) cond591 (
    .clk(cond591_clk),
    .done(cond591_done),
    .in(cond591_in),
    .out(cond591_out),
    .reset(cond591_reset),
    .write_en(cond591_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire591 (
    .in(cond_wire591_in),
    .out(cond_wire591_out)
);
std_reg # (
    .WIDTH(1)
) cond592 (
    .clk(cond592_clk),
    .done(cond592_done),
    .in(cond592_in),
    .out(cond592_out),
    .reset(cond592_reset),
    .write_en(cond592_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire592 (
    .in(cond_wire592_in),
    .out(cond_wire592_out)
);
std_reg # (
    .WIDTH(1)
) cond593 (
    .clk(cond593_clk),
    .done(cond593_done),
    .in(cond593_in),
    .out(cond593_out),
    .reset(cond593_reset),
    .write_en(cond593_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire593 (
    .in(cond_wire593_in),
    .out(cond_wire593_out)
);
std_reg # (
    .WIDTH(1)
) cond594 (
    .clk(cond594_clk),
    .done(cond594_done),
    .in(cond594_in),
    .out(cond594_out),
    .reset(cond594_reset),
    .write_en(cond594_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire594 (
    .in(cond_wire594_in),
    .out(cond_wire594_out)
);
std_reg # (
    .WIDTH(1)
) cond595 (
    .clk(cond595_clk),
    .done(cond595_done),
    .in(cond595_in),
    .out(cond595_out),
    .reset(cond595_reset),
    .write_en(cond595_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire595 (
    .in(cond_wire595_in),
    .out(cond_wire595_out)
);
std_reg # (
    .WIDTH(1)
) cond596 (
    .clk(cond596_clk),
    .done(cond596_done),
    .in(cond596_in),
    .out(cond596_out),
    .reset(cond596_reset),
    .write_en(cond596_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire596 (
    .in(cond_wire596_in),
    .out(cond_wire596_out)
);
std_reg # (
    .WIDTH(1)
) cond597 (
    .clk(cond597_clk),
    .done(cond597_done),
    .in(cond597_in),
    .out(cond597_out),
    .reset(cond597_reset),
    .write_en(cond597_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire597 (
    .in(cond_wire597_in),
    .out(cond_wire597_out)
);
std_reg # (
    .WIDTH(1)
) cond598 (
    .clk(cond598_clk),
    .done(cond598_done),
    .in(cond598_in),
    .out(cond598_out),
    .reset(cond598_reset),
    .write_en(cond598_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire598 (
    .in(cond_wire598_in),
    .out(cond_wire598_out)
);
std_reg # (
    .WIDTH(1)
) cond599 (
    .clk(cond599_clk),
    .done(cond599_done),
    .in(cond599_in),
    .out(cond599_out),
    .reset(cond599_reset),
    .write_en(cond599_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire599 (
    .in(cond_wire599_in),
    .out(cond_wire599_out)
);
std_reg # (
    .WIDTH(1)
) cond600 (
    .clk(cond600_clk),
    .done(cond600_done),
    .in(cond600_in),
    .out(cond600_out),
    .reset(cond600_reset),
    .write_en(cond600_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire600 (
    .in(cond_wire600_in),
    .out(cond_wire600_out)
);
std_reg # (
    .WIDTH(1)
) cond601 (
    .clk(cond601_clk),
    .done(cond601_done),
    .in(cond601_in),
    .out(cond601_out),
    .reset(cond601_reset),
    .write_en(cond601_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire601 (
    .in(cond_wire601_in),
    .out(cond_wire601_out)
);
std_reg # (
    .WIDTH(1)
) cond602 (
    .clk(cond602_clk),
    .done(cond602_done),
    .in(cond602_in),
    .out(cond602_out),
    .reset(cond602_reset),
    .write_en(cond602_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire602 (
    .in(cond_wire602_in),
    .out(cond_wire602_out)
);
std_reg # (
    .WIDTH(1)
) cond603 (
    .clk(cond603_clk),
    .done(cond603_done),
    .in(cond603_in),
    .out(cond603_out),
    .reset(cond603_reset),
    .write_en(cond603_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire603 (
    .in(cond_wire603_in),
    .out(cond_wire603_out)
);
std_reg # (
    .WIDTH(1)
) cond604 (
    .clk(cond604_clk),
    .done(cond604_done),
    .in(cond604_in),
    .out(cond604_out),
    .reset(cond604_reset),
    .write_en(cond604_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire604 (
    .in(cond_wire604_in),
    .out(cond_wire604_out)
);
std_reg # (
    .WIDTH(1)
) cond605 (
    .clk(cond605_clk),
    .done(cond605_done),
    .in(cond605_in),
    .out(cond605_out),
    .reset(cond605_reset),
    .write_en(cond605_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire605 (
    .in(cond_wire605_in),
    .out(cond_wire605_out)
);
std_reg # (
    .WIDTH(1)
) cond606 (
    .clk(cond606_clk),
    .done(cond606_done),
    .in(cond606_in),
    .out(cond606_out),
    .reset(cond606_reset),
    .write_en(cond606_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire606 (
    .in(cond_wire606_in),
    .out(cond_wire606_out)
);
std_reg # (
    .WIDTH(1)
) cond607 (
    .clk(cond607_clk),
    .done(cond607_done),
    .in(cond607_in),
    .out(cond607_out),
    .reset(cond607_reset),
    .write_en(cond607_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire607 (
    .in(cond_wire607_in),
    .out(cond_wire607_out)
);
std_reg # (
    .WIDTH(1)
) cond608 (
    .clk(cond608_clk),
    .done(cond608_done),
    .in(cond608_in),
    .out(cond608_out),
    .reset(cond608_reset),
    .write_en(cond608_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire608 (
    .in(cond_wire608_in),
    .out(cond_wire608_out)
);
std_reg # (
    .WIDTH(1)
) cond609 (
    .clk(cond609_clk),
    .done(cond609_done),
    .in(cond609_in),
    .out(cond609_out),
    .reset(cond609_reset),
    .write_en(cond609_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire609 (
    .in(cond_wire609_in),
    .out(cond_wire609_out)
);
std_reg # (
    .WIDTH(1)
) cond610 (
    .clk(cond610_clk),
    .done(cond610_done),
    .in(cond610_in),
    .out(cond610_out),
    .reset(cond610_reset),
    .write_en(cond610_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire610 (
    .in(cond_wire610_in),
    .out(cond_wire610_out)
);
std_reg # (
    .WIDTH(1)
) cond611 (
    .clk(cond611_clk),
    .done(cond611_done),
    .in(cond611_in),
    .out(cond611_out),
    .reset(cond611_reset),
    .write_en(cond611_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire611 (
    .in(cond_wire611_in),
    .out(cond_wire611_out)
);
std_reg # (
    .WIDTH(1)
) cond612 (
    .clk(cond612_clk),
    .done(cond612_done),
    .in(cond612_in),
    .out(cond612_out),
    .reset(cond612_reset),
    .write_en(cond612_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire612 (
    .in(cond_wire612_in),
    .out(cond_wire612_out)
);
std_reg # (
    .WIDTH(1)
) cond613 (
    .clk(cond613_clk),
    .done(cond613_done),
    .in(cond613_in),
    .out(cond613_out),
    .reset(cond613_reset),
    .write_en(cond613_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire613 (
    .in(cond_wire613_in),
    .out(cond_wire613_out)
);
std_reg # (
    .WIDTH(1)
) cond614 (
    .clk(cond614_clk),
    .done(cond614_done),
    .in(cond614_in),
    .out(cond614_out),
    .reset(cond614_reset),
    .write_en(cond614_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire614 (
    .in(cond_wire614_in),
    .out(cond_wire614_out)
);
std_reg # (
    .WIDTH(1)
) cond615 (
    .clk(cond615_clk),
    .done(cond615_done),
    .in(cond615_in),
    .out(cond615_out),
    .reset(cond615_reset),
    .write_en(cond615_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire615 (
    .in(cond_wire615_in),
    .out(cond_wire615_out)
);
std_reg # (
    .WIDTH(1)
) cond616 (
    .clk(cond616_clk),
    .done(cond616_done),
    .in(cond616_in),
    .out(cond616_out),
    .reset(cond616_reset),
    .write_en(cond616_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire616 (
    .in(cond_wire616_in),
    .out(cond_wire616_out)
);
std_reg # (
    .WIDTH(1)
) cond617 (
    .clk(cond617_clk),
    .done(cond617_done),
    .in(cond617_in),
    .out(cond617_out),
    .reset(cond617_reset),
    .write_en(cond617_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire617 (
    .in(cond_wire617_in),
    .out(cond_wire617_out)
);
std_reg # (
    .WIDTH(1)
) cond618 (
    .clk(cond618_clk),
    .done(cond618_done),
    .in(cond618_in),
    .out(cond618_out),
    .reset(cond618_reset),
    .write_en(cond618_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire618 (
    .in(cond_wire618_in),
    .out(cond_wire618_out)
);
std_reg # (
    .WIDTH(1)
) cond619 (
    .clk(cond619_clk),
    .done(cond619_done),
    .in(cond619_in),
    .out(cond619_out),
    .reset(cond619_reset),
    .write_en(cond619_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire619 (
    .in(cond_wire619_in),
    .out(cond_wire619_out)
);
std_reg # (
    .WIDTH(1)
) cond620 (
    .clk(cond620_clk),
    .done(cond620_done),
    .in(cond620_in),
    .out(cond620_out),
    .reset(cond620_reset),
    .write_en(cond620_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire620 (
    .in(cond_wire620_in),
    .out(cond_wire620_out)
);
std_reg # (
    .WIDTH(1)
) cond621 (
    .clk(cond621_clk),
    .done(cond621_done),
    .in(cond621_in),
    .out(cond621_out),
    .reset(cond621_reset),
    .write_en(cond621_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire621 (
    .in(cond_wire621_in),
    .out(cond_wire621_out)
);
std_reg # (
    .WIDTH(1)
) cond622 (
    .clk(cond622_clk),
    .done(cond622_done),
    .in(cond622_in),
    .out(cond622_out),
    .reset(cond622_reset),
    .write_en(cond622_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire622 (
    .in(cond_wire622_in),
    .out(cond_wire622_out)
);
std_reg # (
    .WIDTH(1)
) cond623 (
    .clk(cond623_clk),
    .done(cond623_done),
    .in(cond623_in),
    .out(cond623_out),
    .reset(cond623_reset),
    .write_en(cond623_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire623 (
    .in(cond_wire623_in),
    .out(cond_wire623_out)
);
std_reg # (
    .WIDTH(1)
) cond624 (
    .clk(cond624_clk),
    .done(cond624_done),
    .in(cond624_in),
    .out(cond624_out),
    .reset(cond624_reset),
    .write_en(cond624_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire624 (
    .in(cond_wire624_in),
    .out(cond_wire624_out)
);
std_reg # (
    .WIDTH(1)
) cond625 (
    .clk(cond625_clk),
    .done(cond625_done),
    .in(cond625_in),
    .out(cond625_out),
    .reset(cond625_reset),
    .write_en(cond625_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire625 (
    .in(cond_wire625_in),
    .out(cond_wire625_out)
);
std_reg # (
    .WIDTH(1)
) cond626 (
    .clk(cond626_clk),
    .done(cond626_done),
    .in(cond626_in),
    .out(cond626_out),
    .reset(cond626_reset),
    .write_en(cond626_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire626 (
    .in(cond_wire626_in),
    .out(cond_wire626_out)
);
std_reg # (
    .WIDTH(1)
) cond627 (
    .clk(cond627_clk),
    .done(cond627_done),
    .in(cond627_in),
    .out(cond627_out),
    .reset(cond627_reset),
    .write_en(cond627_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire627 (
    .in(cond_wire627_in),
    .out(cond_wire627_out)
);
std_reg # (
    .WIDTH(1)
) cond628 (
    .clk(cond628_clk),
    .done(cond628_done),
    .in(cond628_in),
    .out(cond628_out),
    .reset(cond628_reset),
    .write_en(cond628_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire628 (
    .in(cond_wire628_in),
    .out(cond_wire628_out)
);
std_reg # (
    .WIDTH(1)
) cond629 (
    .clk(cond629_clk),
    .done(cond629_done),
    .in(cond629_in),
    .out(cond629_out),
    .reset(cond629_reset),
    .write_en(cond629_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire629 (
    .in(cond_wire629_in),
    .out(cond_wire629_out)
);
std_reg # (
    .WIDTH(1)
) cond630 (
    .clk(cond630_clk),
    .done(cond630_done),
    .in(cond630_in),
    .out(cond630_out),
    .reset(cond630_reset),
    .write_en(cond630_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire630 (
    .in(cond_wire630_in),
    .out(cond_wire630_out)
);
std_reg # (
    .WIDTH(1)
) cond631 (
    .clk(cond631_clk),
    .done(cond631_done),
    .in(cond631_in),
    .out(cond631_out),
    .reset(cond631_reset),
    .write_en(cond631_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire631 (
    .in(cond_wire631_in),
    .out(cond_wire631_out)
);
std_reg # (
    .WIDTH(1)
) cond632 (
    .clk(cond632_clk),
    .done(cond632_done),
    .in(cond632_in),
    .out(cond632_out),
    .reset(cond632_reset),
    .write_en(cond632_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire632 (
    .in(cond_wire632_in),
    .out(cond_wire632_out)
);
std_reg # (
    .WIDTH(1)
) cond633 (
    .clk(cond633_clk),
    .done(cond633_done),
    .in(cond633_in),
    .out(cond633_out),
    .reset(cond633_reset),
    .write_en(cond633_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire633 (
    .in(cond_wire633_in),
    .out(cond_wire633_out)
);
std_reg # (
    .WIDTH(1)
) cond634 (
    .clk(cond634_clk),
    .done(cond634_done),
    .in(cond634_in),
    .out(cond634_out),
    .reset(cond634_reset),
    .write_en(cond634_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire634 (
    .in(cond_wire634_in),
    .out(cond_wire634_out)
);
std_reg # (
    .WIDTH(1)
) cond635 (
    .clk(cond635_clk),
    .done(cond635_done),
    .in(cond635_in),
    .out(cond635_out),
    .reset(cond635_reset),
    .write_en(cond635_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire635 (
    .in(cond_wire635_in),
    .out(cond_wire635_out)
);
std_reg # (
    .WIDTH(1)
) cond636 (
    .clk(cond636_clk),
    .done(cond636_done),
    .in(cond636_in),
    .out(cond636_out),
    .reset(cond636_reset),
    .write_en(cond636_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire636 (
    .in(cond_wire636_in),
    .out(cond_wire636_out)
);
std_reg # (
    .WIDTH(1)
) cond637 (
    .clk(cond637_clk),
    .done(cond637_done),
    .in(cond637_in),
    .out(cond637_out),
    .reset(cond637_reset),
    .write_en(cond637_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire637 (
    .in(cond_wire637_in),
    .out(cond_wire637_out)
);
std_reg # (
    .WIDTH(1)
) cond638 (
    .clk(cond638_clk),
    .done(cond638_done),
    .in(cond638_in),
    .out(cond638_out),
    .reset(cond638_reset),
    .write_en(cond638_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire638 (
    .in(cond_wire638_in),
    .out(cond_wire638_out)
);
std_reg # (
    .WIDTH(1)
) cond639 (
    .clk(cond639_clk),
    .done(cond639_done),
    .in(cond639_in),
    .out(cond639_out),
    .reset(cond639_reset),
    .write_en(cond639_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire639 (
    .in(cond_wire639_in),
    .out(cond_wire639_out)
);
std_reg # (
    .WIDTH(1)
) cond640 (
    .clk(cond640_clk),
    .done(cond640_done),
    .in(cond640_in),
    .out(cond640_out),
    .reset(cond640_reset),
    .write_en(cond640_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire640 (
    .in(cond_wire640_in),
    .out(cond_wire640_out)
);
std_reg # (
    .WIDTH(1)
) cond641 (
    .clk(cond641_clk),
    .done(cond641_done),
    .in(cond641_in),
    .out(cond641_out),
    .reset(cond641_reset),
    .write_en(cond641_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire641 (
    .in(cond_wire641_in),
    .out(cond_wire641_out)
);
std_reg # (
    .WIDTH(1)
) cond642 (
    .clk(cond642_clk),
    .done(cond642_done),
    .in(cond642_in),
    .out(cond642_out),
    .reset(cond642_reset),
    .write_en(cond642_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire642 (
    .in(cond_wire642_in),
    .out(cond_wire642_out)
);
std_reg # (
    .WIDTH(1)
) cond643 (
    .clk(cond643_clk),
    .done(cond643_done),
    .in(cond643_in),
    .out(cond643_out),
    .reset(cond643_reset),
    .write_en(cond643_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire643 (
    .in(cond_wire643_in),
    .out(cond_wire643_out)
);
std_reg # (
    .WIDTH(1)
) cond644 (
    .clk(cond644_clk),
    .done(cond644_done),
    .in(cond644_in),
    .out(cond644_out),
    .reset(cond644_reset),
    .write_en(cond644_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire644 (
    .in(cond_wire644_in),
    .out(cond_wire644_out)
);
std_reg # (
    .WIDTH(1)
) cond645 (
    .clk(cond645_clk),
    .done(cond645_done),
    .in(cond645_in),
    .out(cond645_out),
    .reset(cond645_reset),
    .write_en(cond645_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire645 (
    .in(cond_wire645_in),
    .out(cond_wire645_out)
);
std_reg # (
    .WIDTH(1)
) cond646 (
    .clk(cond646_clk),
    .done(cond646_done),
    .in(cond646_in),
    .out(cond646_out),
    .reset(cond646_reset),
    .write_en(cond646_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire646 (
    .in(cond_wire646_in),
    .out(cond_wire646_out)
);
std_reg # (
    .WIDTH(1)
) cond647 (
    .clk(cond647_clk),
    .done(cond647_done),
    .in(cond647_in),
    .out(cond647_out),
    .reset(cond647_reset),
    .write_en(cond647_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire647 (
    .in(cond_wire647_in),
    .out(cond_wire647_out)
);
std_reg # (
    .WIDTH(1)
) cond648 (
    .clk(cond648_clk),
    .done(cond648_done),
    .in(cond648_in),
    .out(cond648_out),
    .reset(cond648_reset),
    .write_en(cond648_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire648 (
    .in(cond_wire648_in),
    .out(cond_wire648_out)
);
std_reg # (
    .WIDTH(1)
) cond649 (
    .clk(cond649_clk),
    .done(cond649_done),
    .in(cond649_in),
    .out(cond649_out),
    .reset(cond649_reset),
    .write_en(cond649_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire649 (
    .in(cond_wire649_in),
    .out(cond_wire649_out)
);
std_reg # (
    .WIDTH(1)
) cond650 (
    .clk(cond650_clk),
    .done(cond650_done),
    .in(cond650_in),
    .out(cond650_out),
    .reset(cond650_reset),
    .write_en(cond650_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire650 (
    .in(cond_wire650_in),
    .out(cond_wire650_out)
);
std_reg # (
    .WIDTH(1)
) cond651 (
    .clk(cond651_clk),
    .done(cond651_done),
    .in(cond651_in),
    .out(cond651_out),
    .reset(cond651_reset),
    .write_en(cond651_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire651 (
    .in(cond_wire651_in),
    .out(cond_wire651_out)
);
std_reg # (
    .WIDTH(1)
) cond652 (
    .clk(cond652_clk),
    .done(cond652_done),
    .in(cond652_in),
    .out(cond652_out),
    .reset(cond652_reset),
    .write_en(cond652_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire652 (
    .in(cond_wire652_in),
    .out(cond_wire652_out)
);
std_reg # (
    .WIDTH(1)
) cond653 (
    .clk(cond653_clk),
    .done(cond653_done),
    .in(cond653_in),
    .out(cond653_out),
    .reset(cond653_reset),
    .write_en(cond653_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire653 (
    .in(cond_wire653_in),
    .out(cond_wire653_out)
);
std_reg # (
    .WIDTH(1)
) cond654 (
    .clk(cond654_clk),
    .done(cond654_done),
    .in(cond654_in),
    .out(cond654_out),
    .reset(cond654_reset),
    .write_en(cond654_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire654 (
    .in(cond_wire654_in),
    .out(cond_wire654_out)
);
std_reg # (
    .WIDTH(1)
) cond655 (
    .clk(cond655_clk),
    .done(cond655_done),
    .in(cond655_in),
    .out(cond655_out),
    .reset(cond655_reset),
    .write_en(cond655_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire655 (
    .in(cond_wire655_in),
    .out(cond_wire655_out)
);
std_reg # (
    .WIDTH(1)
) cond656 (
    .clk(cond656_clk),
    .done(cond656_done),
    .in(cond656_in),
    .out(cond656_out),
    .reset(cond656_reset),
    .write_en(cond656_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire656 (
    .in(cond_wire656_in),
    .out(cond_wire656_out)
);
std_reg # (
    .WIDTH(1)
) cond657 (
    .clk(cond657_clk),
    .done(cond657_done),
    .in(cond657_in),
    .out(cond657_out),
    .reset(cond657_reset),
    .write_en(cond657_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire657 (
    .in(cond_wire657_in),
    .out(cond_wire657_out)
);
std_reg # (
    .WIDTH(1)
) cond658 (
    .clk(cond658_clk),
    .done(cond658_done),
    .in(cond658_in),
    .out(cond658_out),
    .reset(cond658_reset),
    .write_en(cond658_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire658 (
    .in(cond_wire658_in),
    .out(cond_wire658_out)
);
std_reg # (
    .WIDTH(1)
) cond659 (
    .clk(cond659_clk),
    .done(cond659_done),
    .in(cond659_in),
    .out(cond659_out),
    .reset(cond659_reset),
    .write_en(cond659_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire659 (
    .in(cond_wire659_in),
    .out(cond_wire659_out)
);
std_reg # (
    .WIDTH(1)
) cond660 (
    .clk(cond660_clk),
    .done(cond660_done),
    .in(cond660_in),
    .out(cond660_out),
    .reset(cond660_reset),
    .write_en(cond660_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire660 (
    .in(cond_wire660_in),
    .out(cond_wire660_out)
);
std_reg # (
    .WIDTH(1)
) cond661 (
    .clk(cond661_clk),
    .done(cond661_done),
    .in(cond661_in),
    .out(cond661_out),
    .reset(cond661_reset),
    .write_en(cond661_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire661 (
    .in(cond_wire661_in),
    .out(cond_wire661_out)
);
std_reg # (
    .WIDTH(1)
) cond662 (
    .clk(cond662_clk),
    .done(cond662_done),
    .in(cond662_in),
    .out(cond662_out),
    .reset(cond662_reset),
    .write_en(cond662_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire662 (
    .in(cond_wire662_in),
    .out(cond_wire662_out)
);
std_reg # (
    .WIDTH(1)
) cond663 (
    .clk(cond663_clk),
    .done(cond663_done),
    .in(cond663_in),
    .out(cond663_out),
    .reset(cond663_reset),
    .write_en(cond663_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire663 (
    .in(cond_wire663_in),
    .out(cond_wire663_out)
);
std_reg # (
    .WIDTH(1)
) cond664 (
    .clk(cond664_clk),
    .done(cond664_done),
    .in(cond664_in),
    .out(cond664_out),
    .reset(cond664_reset),
    .write_en(cond664_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire664 (
    .in(cond_wire664_in),
    .out(cond_wire664_out)
);
std_reg # (
    .WIDTH(1)
) cond665 (
    .clk(cond665_clk),
    .done(cond665_done),
    .in(cond665_in),
    .out(cond665_out),
    .reset(cond665_reset),
    .write_en(cond665_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire665 (
    .in(cond_wire665_in),
    .out(cond_wire665_out)
);
std_reg # (
    .WIDTH(1)
) cond666 (
    .clk(cond666_clk),
    .done(cond666_done),
    .in(cond666_in),
    .out(cond666_out),
    .reset(cond666_reset),
    .write_en(cond666_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire666 (
    .in(cond_wire666_in),
    .out(cond_wire666_out)
);
std_reg # (
    .WIDTH(1)
) cond667 (
    .clk(cond667_clk),
    .done(cond667_done),
    .in(cond667_in),
    .out(cond667_out),
    .reset(cond667_reset),
    .write_en(cond667_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire667 (
    .in(cond_wire667_in),
    .out(cond_wire667_out)
);
std_reg # (
    .WIDTH(1)
) cond668 (
    .clk(cond668_clk),
    .done(cond668_done),
    .in(cond668_in),
    .out(cond668_out),
    .reset(cond668_reset),
    .write_en(cond668_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire668 (
    .in(cond_wire668_in),
    .out(cond_wire668_out)
);
std_reg # (
    .WIDTH(1)
) cond669 (
    .clk(cond669_clk),
    .done(cond669_done),
    .in(cond669_in),
    .out(cond669_out),
    .reset(cond669_reset),
    .write_en(cond669_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire669 (
    .in(cond_wire669_in),
    .out(cond_wire669_out)
);
std_reg # (
    .WIDTH(1)
) cond670 (
    .clk(cond670_clk),
    .done(cond670_done),
    .in(cond670_in),
    .out(cond670_out),
    .reset(cond670_reset),
    .write_en(cond670_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire670 (
    .in(cond_wire670_in),
    .out(cond_wire670_out)
);
std_reg # (
    .WIDTH(1)
) cond671 (
    .clk(cond671_clk),
    .done(cond671_done),
    .in(cond671_in),
    .out(cond671_out),
    .reset(cond671_reset),
    .write_en(cond671_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire671 (
    .in(cond_wire671_in),
    .out(cond_wire671_out)
);
std_reg # (
    .WIDTH(1)
) cond672 (
    .clk(cond672_clk),
    .done(cond672_done),
    .in(cond672_in),
    .out(cond672_out),
    .reset(cond672_reset),
    .write_en(cond672_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire672 (
    .in(cond_wire672_in),
    .out(cond_wire672_out)
);
std_reg # (
    .WIDTH(1)
) cond673 (
    .clk(cond673_clk),
    .done(cond673_done),
    .in(cond673_in),
    .out(cond673_out),
    .reset(cond673_reset),
    .write_en(cond673_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire673 (
    .in(cond_wire673_in),
    .out(cond_wire673_out)
);
std_reg # (
    .WIDTH(1)
) cond674 (
    .clk(cond674_clk),
    .done(cond674_done),
    .in(cond674_in),
    .out(cond674_out),
    .reset(cond674_reset),
    .write_en(cond674_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire674 (
    .in(cond_wire674_in),
    .out(cond_wire674_out)
);
std_reg # (
    .WIDTH(1)
) cond675 (
    .clk(cond675_clk),
    .done(cond675_done),
    .in(cond675_in),
    .out(cond675_out),
    .reset(cond675_reset),
    .write_en(cond675_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire675 (
    .in(cond_wire675_in),
    .out(cond_wire675_out)
);
std_reg # (
    .WIDTH(1)
) cond676 (
    .clk(cond676_clk),
    .done(cond676_done),
    .in(cond676_in),
    .out(cond676_out),
    .reset(cond676_reset),
    .write_en(cond676_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire676 (
    .in(cond_wire676_in),
    .out(cond_wire676_out)
);
std_reg # (
    .WIDTH(1)
) cond677 (
    .clk(cond677_clk),
    .done(cond677_done),
    .in(cond677_in),
    .out(cond677_out),
    .reset(cond677_reset),
    .write_en(cond677_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire677 (
    .in(cond_wire677_in),
    .out(cond_wire677_out)
);
std_reg # (
    .WIDTH(1)
) cond678 (
    .clk(cond678_clk),
    .done(cond678_done),
    .in(cond678_in),
    .out(cond678_out),
    .reset(cond678_reset),
    .write_en(cond678_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire678 (
    .in(cond_wire678_in),
    .out(cond_wire678_out)
);
std_reg # (
    .WIDTH(1)
) cond679 (
    .clk(cond679_clk),
    .done(cond679_done),
    .in(cond679_in),
    .out(cond679_out),
    .reset(cond679_reset),
    .write_en(cond679_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire679 (
    .in(cond_wire679_in),
    .out(cond_wire679_out)
);
std_reg # (
    .WIDTH(1)
) cond680 (
    .clk(cond680_clk),
    .done(cond680_done),
    .in(cond680_in),
    .out(cond680_out),
    .reset(cond680_reset),
    .write_en(cond680_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire680 (
    .in(cond_wire680_in),
    .out(cond_wire680_out)
);
std_reg # (
    .WIDTH(1)
) cond681 (
    .clk(cond681_clk),
    .done(cond681_done),
    .in(cond681_in),
    .out(cond681_out),
    .reset(cond681_reset),
    .write_en(cond681_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire681 (
    .in(cond_wire681_in),
    .out(cond_wire681_out)
);
std_reg # (
    .WIDTH(1)
) cond682 (
    .clk(cond682_clk),
    .done(cond682_done),
    .in(cond682_in),
    .out(cond682_out),
    .reset(cond682_reset),
    .write_en(cond682_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire682 (
    .in(cond_wire682_in),
    .out(cond_wire682_out)
);
std_reg # (
    .WIDTH(1)
) cond683 (
    .clk(cond683_clk),
    .done(cond683_done),
    .in(cond683_in),
    .out(cond683_out),
    .reset(cond683_reset),
    .write_en(cond683_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire683 (
    .in(cond_wire683_in),
    .out(cond_wire683_out)
);
std_reg # (
    .WIDTH(1)
) cond684 (
    .clk(cond684_clk),
    .done(cond684_done),
    .in(cond684_in),
    .out(cond684_out),
    .reset(cond684_reset),
    .write_en(cond684_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire684 (
    .in(cond_wire684_in),
    .out(cond_wire684_out)
);
std_reg # (
    .WIDTH(1)
) cond685 (
    .clk(cond685_clk),
    .done(cond685_done),
    .in(cond685_in),
    .out(cond685_out),
    .reset(cond685_reset),
    .write_en(cond685_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire685 (
    .in(cond_wire685_in),
    .out(cond_wire685_out)
);
std_reg # (
    .WIDTH(1)
) cond686 (
    .clk(cond686_clk),
    .done(cond686_done),
    .in(cond686_in),
    .out(cond686_out),
    .reset(cond686_reset),
    .write_en(cond686_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire686 (
    .in(cond_wire686_in),
    .out(cond_wire686_out)
);
std_reg # (
    .WIDTH(1)
) cond687 (
    .clk(cond687_clk),
    .done(cond687_done),
    .in(cond687_in),
    .out(cond687_out),
    .reset(cond687_reset),
    .write_en(cond687_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire687 (
    .in(cond_wire687_in),
    .out(cond_wire687_out)
);
std_reg # (
    .WIDTH(1)
) cond688 (
    .clk(cond688_clk),
    .done(cond688_done),
    .in(cond688_in),
    .out(cond688_out),
    .reset(cond688_reset),
    .write_en(cond688_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire688 (
    .in(cond_wire688_in),
    .out(cond_wire688_out)
);
std_reg # (
    .WIDTH(1)
) cond689 (
    .clk(cond689_clk),
    .done(cond689_done),
    .in(cond689_in),
    .out(cond689_out),
    .reset(cond689_reset),
    .write_en(cond689_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire689 (
    .in(cond_wire689_in),
    .out(cond_wire689_out)
);
std_reg # (
    .WIDTH(1)
) cond690 (
    .clk(cond690_clk),
    .done(cond690_done),
    .in(cond690_in),
    .out(cond690_out),
    .reset(cond690_reset),
    .write_en(cond690_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire690 (
    .in(cond_wire690_in),
    .out(cond_wire690_out)
);
std_reg # (
    .WIDTH(1)
) cond691 (
    .clk(cond691_clk),
    .done(cond691_done),
    .in(cond691_in),
    .out(cond691_out),
    .reset(cond691_reset),
    .write_en(cond691_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire691 (
    .in(cond_wire691_in),
    .out(cond_wire691_out)
);
std_reg # (
    .WIDTH(1)
) cond692 (
    .clk(cond692_clk),
    .done(cond692_done),
    .in(cond692_in),
    .out(cond692_out),
    .reset(cond692_reset),
    .write_en(cond692_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire692 (
    .in(cond_wire692_in),
    .out(cond_wire692_out)
);
std_reg # (
    .WIDTH(1)
) cond693 (
    .clk(cond693_clk),
    .done(cond693_done),
    .in(cond693_in),
    .out(cond693_out),
    .reset(cond693_reset),
    .write_en(cond693_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire693 (
    .in(cond_wire693_in),
    .out(cond_wire693_out)
);
std_reg # (
    .WIDTH(1)
) cond694 (
    .clk(cond694_clk),
    .done(cond694_done),
    .in(cond694_in),
    .out(cond694_out),
    .reset(cond694_reset),
    .write_en(cond694_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire694 (
    .in(cond_wire694_in),
    .out(cond_wire694_out)
);
std_reg # (
    .WIDTH(1)
) cond695 (
    .clk(cond695_clk),
    .done(cond695_done),
    .in(cond695_in),
    .out(cond695_out),
    .reset(cond695_reset),
    .write_en(cond695_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire695 (
    .in(cond_wire695_in),
    .out(cond_wire695_out)
);
std_reg # (
    .WIDTH(1)
) cond696 (
    .clk(cond696_clk),
    .done(cond696_done),
    .in(cond696_in),
    .out(cond696_out),
    .reset(cond696_reset),
    .write_en(cond696_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire696 (
    .in(cond_wire696_in),
    .out(cond_wire696_out)
);
std_reg # (
    .WIDTH(1)
) cond697 (
    .clk(cond697_clk),
    .done(cond697_done),
    .in(cond697_in),
    .out(cond697_out),
    .reset(cond697_reset),
    .write_en(cond697_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire697 (
    .in(cond_wire697_in),
    .out(cond_wire697_out)
);
std_reg # (
    .WIDTH(1)
) cond698 (
    .clk(cond698_clk),
    .done(cond698_done),
    .in(cond698_in),
    .out(cond698_out),
    .reset(cond698_reset),
    .write_en(cond698_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire698 (
    .in(cond_wire698_in),
    .out(cond_wire698_out)
);
std_reg # (
    .WIDTH(1)
) cond699 (
    .clk(cond699_clk),
    .done(cond699_done),
    .in(cond699_in),
    .out(cond699_out),
    .reset(cond699_reset),
    .write_en(cond699_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire699 (
    .in(cond_wire699_in),
    .out(cond_wire699_out)
);
std_reg # (
    .WIDTH(1)
) cond700 (
    .clk(cond700_clk),
    .done(cond700_done),
    .in(cond700_in),
    .out(cond700_out),
    .reset(cond700_reset),
    .write_en(cond700_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire700 (
    .in(cond_wire700_in),
    .out(cond_wire700_out)
);
std_reg # (
    .WIDTH(1)
) cond701 (
    .clk(cond701_clk),
    .done(cond701_done),
    .in(cond701_in),
    .out(cond701_out),
    .reset(cond701_reset),
    .write_en(cond701_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire701 (
    .in(cond_wire701_in),
    .out(cond_wire701_out)
);
std_reg # (
    .WIDTH(1)
) cond702 (
    .clk(cond702_clk),
    .done(cond702_done),
    .in(cond702_in),
    .out(cond702_out),
    .reset(cond702_reset),
    .write_en(cond702_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire702 (
    .in(cond_wire702_in),
    .out(cond_wire702_out)
);
std_reg # (
    .WIDTH(1)
) cond703 (
    .clk(cond703_clk),
    .done(cond703_done),
    .in(cond703_in),
    .out(cond703_out),
    .reset(cond703_reset),
    .write_en(cond703_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire703 (
    .in(cond_wire703_in),
    .out(cond_wire703_out)
);
std_reg # (
    .WIDTH(1)
) cond704 (
    .clk(cond704_clk),
    .done(cond704_done),
    .in(cond704_in),
    .out(cond704_out),
    .reset(cond704_reset),
    .write_en(cond704_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire704 (
    .in(cond_wire704_in),
    .out(cond_wire704_out)
);
std_reg # (
    .WIDTH(1)
) cond705 (
    .clk(cond705_clk),
    .done(cond705_done),
    .in(cond705_in),
    .out(cond705_out),
    .reset(cond705_reset),
    .write_en(cond705_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire705 (
    .in(cond_wire705_in),
    .out(cond_wire705_out)
);
std_reg # (
    .WIDTH(1)
) cond706 (
    .clk(cond706_clk),
    .done(cond706_done),
    .in(cond706_in),
    .out(cond706_out),
    .reset(cond706_reset),
    .write_en(cond706_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire706 (
    .in(cond_wire706_in),
    .out(cond_wire706_out)
);
std_reg # (
    .WIDTH(1)
) cond707 (
    .clk(cond707_clk),
    .done(cond707_done),
    .in(cond707_in),
    .out(cond707_out),
    .reset(cond707_reset),
    .write_en(cond707_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire707 (
    .in(cond_wire707_in),
    .out(cond_wire707_out)
);
std_reg # (
    .WIDTH(1)
) cond708 (
    .clk(cond708_clk),
    .done(cond708_done),
    .in(cond708_in),
    .out(cond708_out),
    .reset(cond708_reset),
    .write_en(cond708_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire708 (
    .in(cond_wire708_in),
    .out(cond_wire708_out)
);
std_reg # (
    .WIDTH(1)
) cond709 (
    .clk(cond709_clk),
    .done(cond709_done),
    .in(cond709_in),
    .out(cond709_out),
    .reset(cond709_reset),
    .write_en(cond709_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire709 (
    .in(cond_wire709_in),
    .out(cond_wire709_out)
);
std_reg # (
    .WIDTH(1)
) cond710 (
    .clk(cond710_clk),
    .done(cond710_done),
    .in(cond710_in),
    .out(cond710_out),
    .reset(cond710_reset),
    .write_en(cond710_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire710 (
    .in(cond_wire710_in),
    .out(cond_wire710_out)
);
std_reg # (
    .WIDTH(1)
) cond711 (
    .clk(cond711_clk),
    .done(cond711_done),
    .in(cond711_in),
    .out(cond711_out),
    .reset(cond711_reset),
    .write_en(cond711_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire711 (
    .in(cond_wire711_in),
    .out(cond_wire711_out)
);
std_reg # (
    .WIDTH(1)
) cond712 (
    .clk(cond712_clk),
    .done(cond712_done),
    .in(cond712_in),
    .out(cond712_out),
    .reset(cond712_reset),
    .write_en(cond712_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire712 (
    .in(cond_wire712_in),
    .out(cond_wire712_out)
);
std_reg # (
    .WIDTH(1)
) cond713 (
    .clk(cond713_clk),
    .done(cond713_done),
    .in(cond713_in),
    .out(cond713_out),
    .reset(cond713_reset),
    .write_en(cond713_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire713 (
    .in(cond_wire713_in),
    .out(cond_wire713_out)
);
std_reg # (
    .WIDTH(1)
) cond714 (
    .clk(cond714_clk),
    .done(cond714_done),
    .in(cond714_in),
    .out(cond714_out),
    .reset(cond714_reset),
    .write_en(cond714_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire714 (
    .in(cond_wire714_in),
    .out(cond_wire714_out)
);
std_reg # (
    .WIDTH(1)
) cond715 (
    .clk(cond715_clk),
    .done(cond715_done),
    .in(cond715_in),
    .out(cond715_out),
    .reset(cond715_reset),
    .write_en(cond715_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire715 (
    .in(cond_wire715_in),
    .out(cond_wire715_out)
);
std_reg # (
    .WIDTH(1)
) cond716 (
    .clk(cond716_clk),
    .done(cond716_done),
    .in(cond716_in),
    .out(cond716_out),
    .reset(cond716_reset),
    .write_en(cond716_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire716 (
    .in(cond_wire716_in),
    .out(cond_wire716_out)
);
std_reg # (
    .WIDTH(1)
) cond717 (
    .clk(cond717_clk),
    .done(cond717_done),
    .in(cond717_in),
    .out(cond717_out),
    .reset(cond717_reset),
    .write_en(cond717_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire717 (
    .in(cond_wire717_in),
    .out(cond_wire717_out)
);
std_reg # (
    .WIDTH(1)
) cond718 (
    .clk(cond718_clk),
    .done(cond718_done),
    .in(cond718_in),
    .out(cond718_out),
    .reset(cond718_reset),
    .write_en(cond718_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire718 (
    .in(cond_wire718_in),
    .out(cond_wire718_out)
);
std_reg # (
    .WIDTH(1)
) cond719 (
    .clk(cond719_clk),
    .done(cond719_done),
    .in(cond719_in),
    .out(cond719_out),
    .reset(cond719_reset),
    .write_en(cond719_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire719 (
    .in(cond_wire719_in),
    .out(cond_wire719_out)
);
std_reg # (
    .WIDTH(1)
) cond720 (
    .clk(cond720_clk),
    .done(cond720_done),
    .in(cond720_in),
    .out(cond720_out),
    .reset(cond720_reset),
    .write_en(cond720_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire720 (
    .in(cond_wire720_in),
    .out(cond_wire720_out)
);
std_reg # (
    .WIDTH(1)
) cond721 (
    .clk(cond721_clk),
    .done(cond721_done),
    .in(cond721_in),
    .out(cond721_out),
    .reset(cond721_reset),
    .write_en(cond721_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire721 (
    .in(cond_wire721_in),
    .out(cond_wire721_out)
);
std_reg # (
    .WIDTH(1)
) cond722 (
    .clk(cond722_clk),
    .done(cond722_done),
    .in(cond722_in),
    .out(cond722_out),
    .reset(cond722_reset),
    .write_en(cond722_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire722 (
    .in(cond_wire722_in),
    .out(cond_wire722_out)
);
std_reg # (
    .WIDTH(1)
) cond723 (
    .clk(cond723_clk),
    .done(cond723_done),
    .in(cond723_in),
    .out(cond723_out),
    .reset(cond723_reset),
    .write_en(cond723_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire723 (
    .in(cond_wire723_in),
    .out(cond_wire723_out)
);
std_reg # (
    .WIDTH(1)
) cond724 (
    .clk(cond724_clk),
    .done(cond724_done),
    .in(cond724_in),
    .out(cond724_out),
    .reset(cond724_reset),
    .write_en(cond724_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire724 (
    .in(cond_wire724_in),
    .out(cond_wire724_out)
);
std_reg # (
    .WIDTH(1)
) cond725 (
    .clk(cond725_clk),
    .done(cond725_done),
    .in(cond725_in),
    .out(cond725_out),
    .reset(cond725_reset),
    .write_en(cond725_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire725 (
    .in(cond_wire725_in),
    .out(cond_wire725_out)
);
std_reg # (
    .WIDTH(1)
) cond726 (
    .clk(cond726_clk),
    .done(cond726_done),
    .in(cond726_in),
    .out(cond726_out),
    .reset(cond726_reset),
    .write_en(cond726_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire726 (
    .in(cond_wire726_in),
    .out(cond_wire726_out)
);
std_reg # (
    .WIDTH(1)
) cond727 (
    .clk(cond727_clk),
    .done(cond727_done),
    .in(cond727_in),
    .out(cond727_out),
    .reset(cond727_reset),
    .write_en(cond727_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire727 (
    .in(cond_wire727_in),
    .out(cond_wire727_out)
);
std_reg # (
    .WIDTH(1)
) cond728 (
    .clk(cond728_clk),
    .done(cond728_done),
    .in(cond728_in),
    .out(cond728_out),
    .reset(cond728_reset),
    .write_en(cond728_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire728 (
    .in(cond_wire728_in),
    .out(cond_wire728_out)
);
std_reg # (
    .WIDTH(1)
) cond729 (
    .clk(cond729_clk),
    .done(cond729_done),
    .in(cond729_in),
    .out(cond729_out),
    .reset(cond729_reset),
    .write_en(cond729_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire729 (
    .in(cond_wire729_in),
    .out(cond_wire729_out)
);
std_reg # (
    .WIDTH(1)
) cond730 (
    .clk(cond730_clk),
    .done(cond730_done),
    .in(cond730_in),
    .out(cond730_out),
    .reset(cond730_reset),
    .write_en(cond730_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire730 (
    .in(cond_wire730_in),
    .out(cond_wire730_out)
);
std_reg # (
    .WIDTH(1)
) cond731 (
    .clk(cond731_clk),
    .done(cond731_done),
    .in(cond731_in),
    .out(cond731_out),
    .reset(cond731_reset),
    .write_en(cond731_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire731 (
    .in(cond_wire731_in),
    .out(cond_wire731_out)
);
std_reg # (
    .WIDTH(1)
) cond732 (
    .clk(cond732_clk),
    .done(cond732_done),
    .in(cond732_in),
    .out(cond732_out),
    .reset(cond732_reset),
    .write_en(cond732_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire732 (
    .in(cond_wire732_in),
    .out(cond_wire732_out)
);
std_reg # (
    .WIDTH(1)
) cond733 (
    .clk(cond733_clk),
    .done(cond733_done),
    .in(cond733_in),
    .out(cond733_out),
    .reset(cond733_reset),
    .write_en(cond733_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire733 (
    .in(cond_wire733_in),
    .out(cond_wire733_out)
);
std_reg # (
    .WIDTH(1)
) cond734 (
    .clk(cond734_clk),
    .done(cond734_done),
    .in(cond734_in),
    .out(cond734_out),
    .reset(cond734_reset),
    .write_en(cond734_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire734 (
    .in(cond_wire734_in),
    .out(cond_wire734_out)
);
std_reg # (
    .WIDTH(1)
) cond735 (
    .clk(cond735_clk),
    .done(cond735_done),
    .in(cond735_in),
    .out(cond735_out),
    .reset(cond735_reset),
    .write_en(cond735_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire735 (
    .in(cond_wire735_in),
    .out(cond_wire735_out)
);
std_reg # (
    .WIDTH(1)
) cond736 (
    .clk(cond736_clk),
    .done(cond736_done),
    .in(cond736_in),
    .out(cond736_out),
    .reset(cond736_reset),
    .write_en(cond736_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire736 (
    .in(cond_wire736_in),
    .out(cond_wire736_out)
);
std_reg # (
    .WIDTH(1)
) cond737 (
    .clk(cond737_clk),
    .done(cond737_done),
    .in(cond737_in),
    .out(cond737_out),
    .reset(cond737_reset),
    .write_en(cond737_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire737 (
    .in(cond_wire737_in),
    .out(cond_wire737_out)
);
std_reg # (
    .WIDTH(1)
) cond738 (
    .clk(cond738_clk),
    .done(cond738_done),
    .in(cond738_in),
    .out(cond738_out),
    .reset(cond738_reset),
    .write_en(cond738_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire738 (
    .in(cond_wire738_in),
    .out(cond_wire738_out)
);
std_reg # (
    .WIDTH(1)
) cond739 (
    .clk(cond739_clk),
    .done(cond739_done),
    .in(cond739_in),
    .out(cond739_out),
    .reset(cond739_reset),
    .write_en(cond739_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire739 (
    .in(cond_wire739_in),
    .out(cond_wire739_out)
);
std_reg # (
    .WIDTH(1)
) cond740 (
    .clk(cond740_clk),
    .done(cond740_done),
    .in(cond740_in),
    .out(cond740_out),
    .reset(cond740_reset),
    .write_en(cond740_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire740 (
    .in(cond_wire740_in),
    .out(cond_wire740_out)
);
std_reg # (
    .WIDTH(1)
) cond741 (
    .clk(cond741_clk),
    .done(cond741_done),
    .in(cond741_in),
    .out(cond741_out),
    .reset(cond741_reset),
    .write_en(cond741_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire741 (
    .in(cond_wire741_in),
    .out(cond_wire741_out)
);
std_reg # (
    .WIDTH(1)
) cond742 (
    .clk(cond742_clk),
    .done(cond742_done),
    .in(cond742_in),
    .out(cond742_out),
    .reset(cond742_reset),
    .write_en(cond742_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire742 (
    .in(cond_wire742_in),
    .out(cond_wire742_out)
);
std_reg # (
    .WIDTH(1)
) cond743 (
    .clk(cond743_clk),
    .done(cond743_done),
    .in(cond743_in),
    .out(cond743_out),
    .reset(cond743_reset),
    .write_en(cond743_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire743 (
    .in(cond_wire743_in),
    .out(cond_wire743_out)
);
std_reg # (
    .WIDTH(1)
) cond744 (
    .clk(cond744_clk),
    .done(cond744_done),
    .in(cond744_in),
    .out(cond744_out),
    .reset(cond744_reset),
    .write_en(cond744_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire744 (
    .in(cond_wire744_in),
    .out(cond_wire744_out)
);
std_reg # (
    .WIDTH(1)
) cond745 (
    .clk(cond745_clk),
    .done(cond745_done),
    .in(cond745_in),
    .out(cond745_out),
    .reset(cond745_reset),
    .write_en(cond745_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire745 (
    .in(cond_wire745_in),
    .out(cond_wire745_out)
);
std_reg # (
    .WIDTH(1)
) cond746 (
    .clk(cond746_clk),
    .done(cond746_done),
    .in(cond746_in),
    .out(cond746_out),
    .reset(cond746_reset),
    .write_en(cond746_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire746 (
    .in(cond_wire746_in),
    .out(cond_wire746_out)
);
std_reg # (
    .WIDTH(1)
) cond747 (
    .clk(cond747_clk),
    .done(cond747_done),
    .in(cond747_in),
    .out(cond747_out),
    .reset(cond747_reset),
    .write_en(cond747_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire747 (
    .in(cond_wire747_in),
    .out(cond_wire747_out)
);
std_reg # (
    .WIDTH(1)
) cond748 (
    .clk(cond748_clk),
    .done(cond748_done),
    .in(cond748_in),
    .out(cond748_out),
    .reset(cond748_reset),
    .write_en(cond748_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire748 (
    .in(cond_wire748_in),
    .out(cond_wire748_out)
);
std_reg # (
    .WIDTH(1)
) cond749 (
    .clk(cond749_clk),
    .done(cond749_done),
    .in(cond749_in),
    .out(cond749_out),
    .reset(cond749_reset),
    .write_en(cond749_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire749 (
    .in(cond_wire749_in),
    .out(cond_wire749_out)
);
std_reg # (
    .WIDTH(1)
) cond750 (
    .clk(cond750_clk),
    .done(cond750_done),
    .in(cond750_in),
    .out(cond750_out),
    .reset(cond750_reset),
    .write_en(cond750_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire750 (
    .in(cond_wire750_in),
    .out(cond_wire750_out)
);
std_reg # (
    .WIDTH(1)
) cond751 (
    .clk(cond751_clk),
    .done(cond751_done),
    .in(cond751_in),
    .out(cond751_out),
    .reset(cond751_reset),
    .write_en(cond751_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire751 (
    .in(cond_wire751_in),
    .out(cond_wire751_out)
);
std_reg # (
    .WIDTH(1)
) cond752 (
    .clk(cond752_clk),
    .done(cond752_done),
    .in(cond752_in),
    .out(cond752_out),
    .reset(cond752_reset),
    .write_en(cond752_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire752 (
    .in(cond_wire752_in),
    .out(cond_wire752_out)
);
std_reg # (
    .WIDTH(1)
) cond753 (
    .clk(cond753_clk),
    .done(cond753_done),
    .in(cond753_in),
    .out(cond753_out),
    .reset(cond753_reset),
    .write_en(cond753_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire753 (
    .in(cond_wire753_in),
    .out(cond_wire753_out)
);
std_reg # (
    .WIDTH(1)
) cond754 (
    .clk(cond754_clk),
    .done(cond754_done),
    .in(cond754_in),
    .out(cond754_out),
    .reset(cond754_reset),
    .write_en(cond754_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire754 (
    .in(cond_wire754_in),
    .out(cond_wire754_out)
);
std_reg # (
    .WIDTH(1)
) cond755 (
    .clk(cond755_clk),
    .done(cond755_done),
    .in(cond755_in),
    .out(cond755_out),
    .reset(cond755_reset),
    .write_en(cond755_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire755 (
    .in(cond_wire755_in),
    .out(cond_wire755_out)
);
std_reg # (
    .WIDTH(1)
) cond756 (
    .clk(cond756_clk),
    .done(cond756_done),
    .in(cond756_in),
    .out(cond756_out),
    .reset(cond756_reset),
    .write_en(cond756_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire756 (
    .in(cond_wire756_in),
    .out(cond_wire756_out)
);
std_reg # (
    .WIDTH(1)
) cond757 (
    .clk(cond757_clk),
    .done(cond757_done),
    .in(cond757_in),
    .out(cond757_out),
    .reset(cond757_reset),
    .write_en(cond757_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire757 (
    .in(cond_wire757_in),
    .out(cond_wire757_out)
);
std_reg # (
    .WIDTH(1)
) cond758 (
    .clk(cond758_clk),
    .done(cond758_done),
    .in(cond758_in),
    .out(cond758_out),
    .reset(cond758_reset),
    .write_en(cond758_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire758 (
    .in(cond_wire758_in),
    .out(cond_wire758_out)
);
std_reg # (
    .WIDTH(1)
) cond759 (
    .clk(cond759_clk),
    .done(cond759_done),
    .in(cond759_in),
    .out(cond759_out),
    .reset(cond759_reset),
    .write_en(cond759_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire759 (
    .in(cond_wire759_in),
    .out(cond_wire759_out)
);
std_reg # (
    .WIDTH(1)
) cond760 (
    .clk(cond760_clk),
    .done(cond760_done),
    .in(cond760_in),
    .out(cond760_out),
    .reset(cond760_reset),
    .write_en(cond760_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire760 (
    .in(cond_wire760_in),
    .out(cond_wire760_out)
);
std_reg # (
    .WIDTH(1)
) cond761 (
    .clk(cond761_clk),
    .done(cond761_done),
    .in(cond761_in),
    .out(cond761_out),
    .reset(cond761_reset),
    .write_en(cond761_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire761 (
    .in(cond_wire761_in),
    .out(cond_wire761_out)
);
std_reg # (
    .WIDTH(1)
) cond762 (
    .clk(cond762_clk),
    .done(cond762_done),
    .in(cond762_in),
    .out(cond762_out),
    .reset(cond762_reset),
    .write_en(cond762_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire762 (
    .in(cond_wire762_in),
    .out(cond_wire762_out)
);
std_reg # (
    .WIDTH(1)
) cond763 (
    .clk(cond763_clk),
    .done(cond763_done),
    .in(cond763_in),
    .out(cond763_out),
    .reset(cond763_reset),
    .write_en(cond763_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire763 (
    .in(cond_wire763_in),
    .out(cond_wire763_out)
);
std_reg # (
    .WIDTH(1)
) cond764 (
    .clk(cond764_clk),
    .done(cond764_done),
    .in(cond764_in),
    .out(cond764_out),
    .reset(cond764_reset),
    .write_en(cond764_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire764 (
    .in(cond_wire764_in),
    .out(cond_wire764_out)
);
std_reg # (
    .WIDTH(1)
) cond765 (
    .clk(cond765_clk),
    .done(cond765_done),
    .in(cond765_in),
    .out(cond765_out),
    .reset(cond765_reset),
    .write_en(cond765_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire765 (
    .in(cond_wire765_in),
    .out(cond_wire765_out)
);
std_reg # (
    .WIDTH(1)
) cond766 (
    .clk(cond766_clk),
    .done(cond766_done),
    .in(cond766_in),
    .out(cond766_out),
    .reset(cond766_reset),
    .write_en(cond766_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire766 (
    .in(cond_wire766_in),
    .out(cond_wire766_out)
);
std_reg # (
    .WIDTH(1)
) cond767 (
    .clk(cond767_clk),
    .done(cond767_done),
    .in(cond767_in),
    .out(cond767_out),
    .reset(cond767_reset),
    .write_en(cond767_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire767 (
    .in(cond_wire767_in),
    .out(cond_wire767_out)
);
std_reg # (
    .WIDTH(1)
) cond768 (
    .clk(cond768_clk),
    .done(cond768_done),
    .in(cond768_in),
    .out(cond768_out),
    .reset(cond768_reset),
    .write_en(cond768_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire768 (
    .in(cond_wire768_in),
    .out(cond_wire768_out)
);
std_reg # (
    .WIDTH(1)
) cond769 (
    .clk(cond769_clk),
    .done(cond769_done),
    .in(cond769_in),
    .out(cond769_out),
    .reset(cond769_reset),
    .write_en(cond769_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire769 (
    .in(cond_wire769_in),
    .out(cond_wire769_out)
);
std_reg # (
    .WIDTH(1)
) cond770 (
    .clk(cond770_clk),
    .done(cond770_done),
    .in(cond770_in),
    .out(cond770_out),
    .reset(cond770_reset),
    .write_en(cond770_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire770 (
    .in(cond_wire770_in),
    .out(cond_wire770_out)
);
std_reg # (
    .WIDTH(1)
) cond771 (
    .clk(cond771_clk),
    .done(cond771_done),
    .in(cond771_in),
    .out(cond771_out),
    .reset(cond771_reset),
    .write_en(cond771_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire771 (
    .in(cond_wire771_in),
    .out(cond_wire771_out)
);
std_reg # (
    .WIDTH(1)
) cond772 (
    .clk(cond772_clk),
    .done(cond772_done),
    .in(cond772_in),
    .out(cond772_out),
    .reset(cond772_reset),
    .write_en(cond772_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire772 (
    .in(cond_wire772_in),
    .out(cond_wire772_out)
);
std_reg # (
    .WIDTH(1)
) cond773 (
    .clk(cond773_clk),
    .done(cond773_done),
    .in(cond773_in),
    .out(cond773_out),
    .reset(cond773_reset),
    .write_en(cond773_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire773 (
    .in(cond_wire773_in),
    .out(cond_wire773_out)
);
std_reg # (
    .WIDTH(1)
) cond774 (
    .clk(cond774_clk),
    .done(cond774_done),
    .in(cond774_in),
    .out(cond774_out),
    .reset(cond774_reset),
    .write_en(cond774_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire774 (
    .in(cond_wire774_in),
    .out(cond_wire774_out)
);
std_reg # (
    .WIDTH(1)
) cond775 (
    .clk(cond775_clk),
    .done(cond775_done),
    .in(cond775_in),
    .out(cond775_out),
    .reset(cond775_reset),
    .write_en(cond775_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire775 (
    .in(cond_wire775_in),
    .out(cond_wire775_out)
);
std_reg # (
    .WIDTH(1)
) cond776 (
    .clk(cond776_clk),
    .done(cond776_done),
    .in(cond776_in),
    .out(cond776_out),
    .reset(cond776_reset),
    .write_en(cond776_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire776 (
    .in(cond_wire776_in),
    .out(cond_wire776_out)
);
std_reg # (
    .WIDTH(1)
) cond777 (
    .clk(cond777_clk),
    .done(cond777_done),
    .in(cond777_in),
    .out(cond777_out),
    .reset(cond777_reset),
    .write_en(cond777_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire777 (
    .in(cond_wire777_in),
    .out(cond_wire777_out)
);
std_reg # (
    .WIDTH(1)
) cond778 (
    .clk(cond778_clk),
    .done(cond778_done),
    .in(cond778_in),
    .out(cond778_out),
    .reset(cond778_reset),
    .write_en(cond778_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire778 (
    .in(cond_wire778_in),
    .out(cond_wire778_out)
);
std_reg # (
    .WIDTH(1)
) cond779 (
    .clk(cond779_clk),
    .done(cond779_done),
    .in(cond779_in),
    .out(cond779_out),
    .reset(cond779_reset),
    .write_en(cond779_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire779 (
    .in(cond_wire779_in),
    .out(cond_wire779_out)
);
std_reg # (
    .WIDTH(1)
) cond780 (
    .clk(cond780_clk),
    .done(cond780_done),
    .in(cond780_in),
    .out(cond780_out),
    .reset(cond780_reset),
    .write_en(cond780_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire780 (
    .in(cond_wire780_in),
    .out(cond_wire780_out)
);
std_reg # (
    .WIDTH(1)
) cond781 (
    .clk(cond781_clk),
    .done(cond781_done),
    .in(cond781_in),
    .out(cond781_out),
    .reset(cond781_reset),
    .write_en(cond781_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire781 (
    .in(cond_wire781_in),
    .out(cond_wire781_out)
);
std_reg # (
    .WIDTH(1)
) cond782 (
    .clk(cond782_clk),
    .done(cond782_done),
    .in(cond782_in),
    .out(cond782_out),
    .reset(cond782_reset),
    .write_en(cond782_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire782 (
    .in(cond_wire782_in),
    .out(cond_wire782_out)
);
std_reg # (
    .WIDTH(1)
) cond783 (
    .clk(cond783_clk),
    .done(cond783_done),
    .in(cond783_in),
    .out(cond783_out),
    .reset(cond783_reset),
    .write_en(cond783_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire783 (
    .in(cond_wire783_in),
    .out(cond_wire783_out)
);
std_reg # (
    .WIDTH(1)
) cond784 (
    .clk(cond784_clk),
    .done(cond784_done),
    .in(cond784_in),
    .out(cond784_out),
    .reset(cond784_reset),
    .write_en(cond784_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire784 (
    .in(cond_wire784_in),
    .out(cond_wire784_out)
);
std_reg # (
    .WIDTH(1)
) cond785 (
    .clk(cond785_clk),
    .done(cond785_done),
    .in(cond785_in),
    .out(cond785_out),
    .reset(cond785_reset),
    .write_en(cond785_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire785 (
    .in(cond_wire785_in),
    .out(cond_wire785_out)
);
std_reg # (
    .WIDTH(1)
) cond786 (
    .clk(cond786_clk),
    .done(cond786_done),
    .in(cond786_in),
    .out(cond786_out),
    .reset(cond786_reset),
    .write_en(cond786_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire786 (
    .in(cond_wire786_in),
    .out(cond_wire786_out)
);
std_reg # (
    .WIDTH(1)
) cond787 (
    .clk(cond787_clk),
    .done(cond787_done),
    .in(cond787_in),
    .out(cond787_out),
    .reset(cond787_reset),
    .write_en(cond787_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire787 (
    .in(cond_wire787_in),
    .out(cond_wire787_out)
);
std_reg # (
    .WIDTH(1)
) cond788 (
    .clk(cond788_clk),
    .done(cond788_done),
    .in(cond788_in),
    .out(cond788_out),
    .reset(cond788_reset),
    .write_en(cond788_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire788 (
    .in(cond_wire788_in),
    .out(cond_wire788_out)
);
std_reg # (
    .WIDTH(1)
) cond789 (
    .clk(cond789_clk),
    .done(cond789_done),
    .in(cond789_in),
    .out(cond789_out),
    .reset(cond789_reset),
    .write_en(cond789_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire789 (
    .in(cond_wire789_in),
    .out(cond_wire789_out)
);
std_reg # (
    .WIDTH(1)
) cond790 (
    .clk(cond790_clk),
    .done(cond790_done),
    .in(cond790_in),
    .out(cond790_out),
    .reset(cond790_reset),
    .write_en(cond790_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire790 (
    .in(cond_wire790_in),
    .out(cond_wire790_out)
);
std_reg # (
    .WIDTH(1)
) cond791 (
    .clk(cond791_clk),
    .done(cond791_done),
    .in(cond791_in),
    .out(cond791_out),
    .reset(cond791_reset),
    .write_en(cond791_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire791 (
    .in(cond_wire791_in),
    .out(cond_wire791_out)
);
std_reg # (
    .WIDTH(1)
) cond792 (
    .clk(cond792_clk),
    .done(cond792_done),
    .in(cond792_in),
    .out(cond792_out),
    .reset(cond792_reset),
    .write_en(cond792_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire792 (
    .in(cond_wire792_in),
    .out(cond_wire792_out)
);
std_reg # (
    .WIDTH(1)
) cond793 (
    .clk(cond793_clk),
    .done(cond793_done),
    .in(cond793_in),
    .out(cond793_out),
    .reset(cond793_reset),
    .write_en(cond793_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire793 (
    .in(cond_wire793_in),
    .out(cond_wire793_out)
);
std_reg # (
    .WIDTH(1)
) cond794 (
    .clk(cond794_clk),
    .done(cond794_done),
    .in(cond794_in),
    .out(cond794_out),
    .reset(cond794_reset),
    .write_en(cond794_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire794 (
    .in(cond_wire794_in),
    .out(cond_wire794_out)
);
std_reg # (
    .WIDTH(1)
) cond795 (
    .clk(cond795_clk),
    .done(cond795_done),
    .in(cond795_in),
    .out(cond795_out),
    .reset(cond795_reset),
    .write_en(cond795_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire795 (
    .in(cond_wire795_in),
    .out(cond_wire795_out)
);
std_reg # (
    .WIDTH(1)
) cond796 (
    .clk(cond796_clk),
    .done(cond796_done),
    .in(cond796_in),
    .out(cond796_out),
    .reset(cond796_reset),
    .write_en(cond796_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire796 (
    .in(cond_wire796_in),
    .out(cond_wire796_out)
);
std_reg # (
    .WIDTH(1)
) cond797 (
    .clk(cond797_clk),
    .done(cond797_done),
    .in(cond797_in),
    .out(cond797_out),
    .reset(cond797_reset),
    .write_en(cond797_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire797 (
    .in(cond_wire797_in),
    .out(cond_wire797_out)
);
std_reg # (
    .WIDTH(1)
) cond798 (
    .clk(cond798_clk),
    .done(cond798_done),
    .in(cond798_in),
    .out(cond798_out),
    .reset(cond798_reset),
    .write_en(cond798_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire798 (
    .in(cond_wire798_in),
    .out(cond_wire798_out)
);
std_reg # (
    .WIDTH(1)
) cond799 (
    .clk(cond799_clk),
    .done(cond799_done),
    .in(cond799_in),
    .out(cond799_out),
    .reset(cond799_reset),
    .write_en(cond799_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire799 (
    .in(cond_wire799_in),
    .out(cond_wire799_out)
);
std_reg # (
    .WIDTH(1)
) cond800 (
    .clk(cond800_clk),
    .done(cond800_done),
    .in(cond800_in),
    .out(cond800_out),
    .reset(cond800_reset),
    .write_en(cond800_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire800 (
    .in(cond_wire800_in),
    .out(cond_wire800_out)
);
std_reg # (
    .WIDTH(1)
) cond801 (
    .clk(cond801_clk),
    .done(cond801_done),
    .in(cond801_in),
    .out(cond801_out),
    .reset(cond801_reset),
    .write_en(cond801_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire801 (
    .in(cond_wire801_in),
    .out(cond_wire801_out)
);
std_reg # (
    .WIDTH(1)
) cond802 (
    .clk(cond802_clk),
    .done(cond802_done),
    .in(cond802_in),
    .out(cond802_out),
    .reset(cond802_reset),
    .write_en(cond802_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire802 (
    .in(cond_wire802_in),
    .out(cond_wire802_out)
);
std_reg # (
    .WIDTH(1)
) cond803 (
    .clk(cond803_clk),
    .done(cond803_done),
    .in(cond803_in),
    .out(cond803_out),
    .reset(cond803_reset),
    .write_en(cond803_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire803 (
    .in(cond_wire803_in),
    .out(cond_wire803_out)
);
std_reg # (
    .WIDTH(1)
) cond804 (
    .clk(cond804_clk),
    .done(cond804_done),
    .in(cond804_in),
    .out(cond804_out),
    .reset(cond804_reset),
    .write_en(cond804_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire804 (
    .in(cond_wire804_in),
    .out(cond_wire804_out)
);
std_reg # (
    .WIDTH(1)
) cond805 (
    .clk(cond805_clk),
    .done(cond805_done),
    .in(cond805_in),
    .out(cond805_out),
    .reset(cond805_reset),
    .write_en(cond805_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire805 (
    .in(cond_wire805_in),
    .out(cond_wire805_out)
);
std_reg # (
    .WIDTH(1)
) cond806 (
    .clk(cond806_clk),
    .done(cond806_done),
    .in(cond806_in),
    .out(cond806_out),
    .reset(cond806_reset),
    .write_en(cond806_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire806 (
    .in(cond_wire806_in),
    .out(cond_wire806_out)
);
std_reg # (
    .WIDTH(1)
) cond807 (
    .clk(cond807_clk),
    .done(cond807_done),
    .in(cond807_in),
    .out(cond807_out),
    .reset(cond807_reset),
    .write_en(cond807_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire807 (
    .in(cond_wire807_in),
    .out(cond_wire807_out)
);
std_reg # (
    .WIDTH(1)
) cond808 (
    .clk(cond808_clk),
    .done(cond808_done),
    .in(cond808_in),
    .out(cond808_out),
    .reset(cond808_reset),
    .write_en(cond808_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire808 (
    .in(cond_wire808_in),
    .out(cond_wire808_out)
);
std_reg # (
    .WIDTH(1)
) cond809 (
    .clk(cond809_clk),
    .done(cond809_done),
    .in(cond809_in),
    .out(cond809_out),
    .reset(cond809_reset),
    .write_en(cond809_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire809 (
    .in(cond_wire809_in),
    .out(cond_wire809_out)
);
std_reg # (
    .WIDTH(1)
) cond810 (
    .clk(cond810_clk),
    .done(cond810_done),
    .in(cond810_in),
    .out(cond810_out),
    .reset(cond810_reset),
    .write_en(cond810_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire810 (
    .in(cond_wire810_in),
    .out(cond_wire810_out)
);
std_reg # (
    .WIDTH(1)
) cond811 (
    .clk(cond811_clk),
    .done(cond811_done),
    .in(cond811_in),
    .out(cond811_out),
    .reset(cond811_reset),
    .write_en(cond811_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire811 (
    .in(cond_wire811_in),
    .out(cond_wire811_out)
);
std_reg # (
    .WIDTH(1)
) cond812 (
    .clk(cond812_clk),
    .done(cond812_done),
    .in(cond812_in),
    .out(cond812_out),
    .reset(cond812_reset),
    .write_en(cond812_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire812 (
    .in(cond_wire812_in),
    .out(cond_wire812_out)
);
std_reg # (
    .WIDTH(1)
) cond813 (
    .clk(cond813_clk),
    .done(cond813_done),
    .in(cond813_in),
    .out(cond813_out),
    .reset(cond813_reset),
    .write_en(cond813_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire813 (
    .in(cond_wire813_in),
    .out(cond_wire813_out)
);
std_reg # (
    .WIDTH(1)
) cond814 (
    .clk(cond814_clk),
    .done(cond814_done),
    .in(cond814_in),
    .out(cond814_out),
    .reset(cond814_reset),
    .write_en(cond814_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire814 (
    .in(cond_wire814_in),
    .out(cond_wire814_out)
);
std_reg # (
    .WIDTH(1)
) cond815 (
    .clk(cond815_clk),
    .done(cond815_done),
    .in(cond815_in),
    .out(cond815_out),
    .reset(cond815_reset),
    .write_en(cond815_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire815 (
    .in(cond_wire815_in),
    .out(cond_wire815_out)
);
std_reg # (
    .WIDTH(1)
) cond816 (
    .clk(cond816_clk),
    .done(cond816_done),
    .in(cond816_in),
    .out(cond816_out),
    .reset(cond816_reset),
    .write_en(cond816_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire816 (
    .in(cond_wire816_in),
    .out(cond_wire816_out)
);
std_reg # (
    .WIDTH(1)
) cond817 (
    .clk(cond817_clk),
    .done(cond817_done),
    .in(cond817_in),
    .out(cond817_out),
    .reset(cond817_reset),
    .write_en(cond817_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire817 (
    .in(cond_wire817_in),
    .out(cond_wire817_out)
);
std_reg # (
    .WIDTH(1)
) cond818 (
    .clk(cond818_clk),
    .done(cond818_done),
    .in(cond818_in),
    .out(cond818_out),
    .reset(cond818_reset),
    .write_en(cond818_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire818 (
    .in(cond_wire818_in),
    .out(cond_wire818_out)
);
std_reg # (
    .WIDTH(1)
) cond819 (
    .clk(cond819_clk),
    .done(cond819_done),
    .in(cond819_in),
    .out(cond819_out),
    .reset(cond819_reset),
    .write_en(cond819_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire819 (
    .in(cond_wire819_in),
    .out(cond_wire819_out)
);
std_reg # (
    .WIDTH(1)
) cond820 (
    .clk(cond820_clk),
    .done(cond820_done),
    .in(cond820_in),
    .out(cond820_out),
    .reset(cond820_reset),
    .write_en(cond820_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire820 (
    .in(cond_wire820_in),
    .out(cond_wire820_out)
);
std_reg # (
    .WIDTH(1)
) cond821 (
    .clk(cond821_clk),
    .done(cond821_done),
    .in(cond821_in),
    .out(cond821_out),
    .reset(cond821_reset),
    .write_en(cond821_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire821 (
    .in(cond_wire821_in),
    .out(cond_wire821_out)
);
std_reg # (
    .WIDTH(1)
) cond822 (
    .clk(cond822_clk),
    .done(cond822_done),
    .in(cond822_in),
    .out(cond822_out),
    .reset(cond822_reset),
    .write_en(cond822_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire822 (
    .in(cond_wire822_in),
    .out(cond_wire822_out)
);
std_reg # (
    .WIDTH(1)
) cond823 (
    .clk(cond823_clk),
    .done(cond823_done),
    .in(cond823_in),
    .out(cond823_out),
    .reset(cond823_reset),
    .write_en(cond823_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire823 (
    .in(cond_wire823_in),
    .out(cond_wire823_out)
);
std_reg # (
    .WIDTH(1)
) cond824 (
    .clk(cond824_clk),
    .done(cond824_done),
    .in(cond824_in),
    .out(cond824_out),
    .reset(cond824_reset),
    .write_en(cond824_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire824 (
    .in(cond_wire824_in),
    .out(cond_wire824_out)
);
std_reg # (
    .WIDTH(1)
) cond825 (
    .clk(cond825_clk),
    .done(cond825_done),
    .in(cond825_in),
    .out(cond825_out),
    .reset(cond825_reset),
    .write_en(cond825_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire825 (
    .in(cond_wire825_in),
    .out(cond_wire825_out)
);
std_reg # (
    .WIDTH(1)
) cond826 (
    .clk(cond826_clk),
    .done(cond826_done),
    .in(cond826_in),
    .out(cond826_out),
    .reset(cond826_reset),
    .write_en(cond826_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire826 (
    .in(cond_wire826_in),
    .out(cond_wire826_out)
);
std_reg # (
    .WIDTH(1)
) cond827 (
    .clk(cond827_clk),
    .done(cond827_done),
    .in(cond827_in),
    .out(cond827_out),
    .reset(cond827_reset),
    .write_en(cond827_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire827 (
    .in(cond_wire827_in),
    .out(cond_wire827_out)
);
std_reg # (
    .WIDTH(1)
) cond828 (
    .clk(cond828_clk),
    .done(cond828_done),
    .in(cond828_in),
    .out(cond828_out),
    .reset(cond828_reset),
    .write_en(cond828_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire828 (
    .in(cond_wire828_in),
    .out(cond_wire828_out)
);
std_reg # (
    .WIDTH(1)
) cond829 (
    .clk(cond829_clk),
    .done(cond829_done),
    .in(cond829_in),
    .out(cond829_out),
    .reset(cond829_reset),
    .write_en(cond829_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire829 (
    .in(cond_wire829_in),
    .out(cond_wire829_out)
);
std_reg # (
    .WIDTH(1)
) cond830 (
    .clk(cond830_clk),
    .done(cond830_done),
    .in(cond830_in),
    .out(cond830_out),
    .reset(cond830_reset),
    .write_en(cond830_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire830 (
    .in(cond_wire830_in),
    .out(cond_wire830_out)
);
std_reg # (
    .WIDTH(1)
) cond831 (
    .clk(cond831_clk),
    .done(cond831_done),
    .in(cond831_in),
    .out(cond831_out),
    .reset(cond831_reset),
    .write_en(cond831_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire831 (
    .in(cond_wire831_in),
    .out(cond_wire831_out)
);
std_reg # (
    .WIDTH(1)
) cond832 (
    .clk(cond832_clk),
    .done(cond832_done),
    .in(cond832_in),
    .out(cond832_out),
    .reset(cond832_reset),
    .write_en(cond832_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire832 (
    .in(cond_wire832_in),
    .out(cond_wire832_out)
);
std_reg # (
    .WIDTH(1)
) cond833 (
    .clk(cond833_clk),
    .done(cond833_done),
    .in(cond833_in),
    .out(cond833_out),
    .reset(cond833_reset),
    .write_en(cond833_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire833 (
    .in(cond_wire833_in),
    .out(cond_wire833_out)
);
std_reg # (
    .WIDTH(1)
) cond834 (
    .clk(cond834_clk),
    .done(cond834_done),
    .in(cond834_in),
    .out(cond834_out),
    .reset(cond834_reset),
    .write_en(cond834_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire834 (
    .in(cond_wire834_in),
    .out(cond_wire834_out)
);
std_reg # (
    .WIDTH(1)
) cond835 (
    .clk(cond835_clk),
    .done(cond835_done),
    .in(cond835_in),
    .out(cond835_out),
    .reset(cond835_reset),
    .write_en(cond835_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire835 (
    .in(cond_wire835_in),
    .out(cond_wire835_out)
);
std_reg # (
    .WIDTH(1)
) cond836 (
    .clk(cond836_clk),
    .done(cond836_done),
    .in(cond836_in),
    .out(cond836_out),
    .reset(cond836_reset),
    .write_en(cond836_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire836 (
    .in(cond_wire836_in),
    .out(cond_wire836_out)
);
std_reg # (
    .WIDTH(1)
) cond837 (
    .clk(cond837_clk),
    .done(cond837_done),
    .in(cond837_in),
    .out(cond837_out),
    .reset(cond837_reset),
    .write_en(cond837_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire837 (
    .in(cond_wire837_in),
    .out(cond_wire837_out)
);
std_reg # (
    .WIDTH(1)
) cond838 (
    .clk(cond838_clk),
    .done(cond838_done),
    .in(cond838_in),
    .out(cond838_out),
    .reset(cond838_reset),
    .write_en(cond838_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire838 (
    .in(cond_wire838_in),
    .out(cond_wire838_out)
);
std_reg # (
    .WIDTH(1)
) cond839 (
    .clk(cond839_clk),
    .done(cond839_done),
    .in(cond839_in),
    .out(cond839_out),
    .reset(cond839_reset),
    .write_en(cond839_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire839 (
    .in(cond_wire839_in),
    .out(cond_wire839_out)
);
std_reg # (
    .WIDTH(1)
) cond840 (
    .clk(cond840_clk),
    .done(cond840_done),
    .in(cond840_in),
    .out(cond840_out),
    .reset(cond840_reset),
    .write_en(cond840_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire840 (
    .in(cond_wire840_in),
    .out(cond_wire840_out)
);
std_reg # (
    .WIDTH(1)
) cond841 (
    .clk(cond841_clk),
    .done(cond841_done),
    .in(cond841_in),
    .out(cond841_out),
    .reset(cond841_reset),
    .write_en(cond841_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire841 (
    .in(cond_wire841_in),
    .out(cond_wire841_out)
);
std_reg # (
    .WIDTH(1)
) cond842 (
    .clk(cond842_clk),
    .done(cond842_done),
    .in(cond842_in),
    .out(cond842_out),
    .reset(cond842_reset),
    .write_en(cond842_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire842 (
    .in(cond_wire842_in),
    .out(cond_wire842_out)
);
std_reg # (
    .WIDTH(1)
) cond843 (
    .clk(cond843_clk),
    .done(cond843_done),
    .in(cond843_in),
    .out(cond843_out),
    .reset(cond843_reset),
    .write_en(cond843_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire843 (
    .in(cond_wire843_in),
    .out(cond_wire843_out)
);
std_reg # (
    .WIDTH(1)
) cond844 (
    .clk(cond844_clk),
    .done(cond844_done),
    .in(cond844_in),
    .out(cond844_out),
    .reset(cond844_reset),
    .write_en(cond844_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire844 (
    .in(cond_wire844_in),
    .out(cond_wire844_out)
);
std_reg # (
    .WIDTH(1)
) cond845 (
    .clk(cond845_clk),
    .done(cond845_done),
    .in(cond845_in),
    .out(cond845_out),
    .reset(cond845_reset),
    .write_en(cond845_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire845 (
    .in(cond_wire845_in),
    .out(cond_wire845_out)
);
std_reg # (
    .WIDTH(1)
) cond846 (
    .clk(cond846_clk),
    .done(cond846_done),
    .in(cond846_in),
    .out(cond846_out),
    .reset(cond846_reset),
    .write_en(cond846_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire846 (
    .in(cond_wire846_in),
    .out(cond_wire846_out)
);
std_reg # (
    .WIDTH(1)
) cond847 (
    .clk(cond847_clk),
    .done(cond847_done),
    .in(cond847_in),
    .out(cond847_out),
    .reset(cond847_reset),
    .write_en(cond847_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire847 (
    .in(cond_wire847_in),
    .out(cond_wire847_out)
);
std_reg # (
    .WIDTH(1)
) cond848 (
    .clk(cond848_clk),
    .done(cond848_done),
    .in(cond848_in),
    .out(cond848_out),
    .reset(cond848_reset),
    .write_en(cond848_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire848 (
    .in(cond_wire848_in),
    .out(cond_wire848_out)
);
std_reg # (
    .WIDTH(1)
) cond849 (
    .clk(cond849_clk),
    .done(cond849_done),
    .in(cond849_in),
    .out(cond849_out),
    .reset(cond849_reset),
    .write_en(cond849_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire849 (
    .in(cond_wire849_in),
    .out(cond_wire849_out)
);
std_reg # (
    .WIDTH(1)
) cond850 (
    .clk(cond850_clk),
    .done(cond850_done),
    .in(cond850_in),
    .out(cond850_out),
    .reset(cond850_reset),
    .write_en(cond850_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire850 (
    .in(cond_wire850_in),
    .out(cond_wire850_out)
);
std_reg # (
    .WIDTH(1)
) cond851 (
    .clk(cond851_clk),
    .done(cond851_done),
    .in(cond851_in),
    .out(cond851_out),
    .reset(cond851_reset),
    .write_en(cond851_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire851 (
    .in(cond_wire851_in),
    .out(cond_wire851_out)
);
std_reg # (
    .WIDTH(1)
) cond852 (
    .clk(cond852_clk),
    .done(cond852_done),
    .in(cond852_in),
    .out(cond852_out),
    .reset(cond852_reset),
    .write_en(cond852_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire852 (
    .in(cond_wire852_in),
    .out(cond_wire852_out)
);
std_reg # (
    .WIDTH(1)
) cond853 (
    .clk(cond853_clk),
    .done(cond853_done),
    .in(cond853_in),
    .out(cond853_out),
    .reset(cond853_reset),
    .write_en(cond853_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire853 (
    .in(cond_wire853_in),
    .out(cond_wire853_out)
);
std_reg # (
    .WIDTH(1)
) cond854 (
    .clk(cond854_clk),
    .done(cond854_done),
    .in(cond854_in),
    .out(cond854_out),
    .reset(cond854_reset),
    .write_en(cond854_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire854 (
    .in(cond_wire854_in),
    .out(cond_wire854_out)
);
std_reg # (
    .WIDTH(1)
) cond855 (
    .clk(cond855_clk),
    .done(cond855_done),
    .in(cond855_in),
    .out(cond855_out),
    .reset(cond855_reset),
    .write_en(cond855_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire855 (
    .in(cond_wire855_in),
    .out(cond_wire855_out)
);
std_reg # (
    .WIDTH(1)
) cond856 (
    .clk(cond856_clk),
    .done(cond856_done),
    .in(cond856_in),
    .out(cond856_out),
    .reset(cond856_reset),
    .write_en(cond856_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire856 (
    .in(cond_wire856_in),
    .out(cond_wire856_out)
);
std_reg # (
    .WIDTH(1)
) cond857 (
    .clk(cond857_clk),
    .done(cond857_done),
    .in(cond857_in),
    .out(cond857_out),
    .reset(cond857_reset),
    .write_en(cond857_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire857 (
    .in(cond_wire857_in),
    .out(cond_wire857_out)
);
std_reg # (
    .WIDTH(1)
) cond858 (
    .clk(cond858_clk),
    .done(cond858_done),
    .in(cond858_in),
    .out(cond858_out),
    .reset(cond858_reset),
    .write_en(cond858_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire858 (
    .in(cond_wire858_in),
    .out(cond_wire858_out)
);
std_reg # (
    .WIDTH(1)
) cond859 (
    .clk(cond859_clk),
    .done(cond859_done),
    .in(cond859_in),
    .out(cond859_out),
    .reset(cond859_reset),
    .write_en(cond859_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire859 (
    .in(cond_wire859_in),
    .out(cond_wire859_out)
);
std_reg # (
    .WIDTH(1)
) cond860 (
    .clk(cond860_clk),
    .done(cond860_done),
    .in(cond860_in),
    .out(cond860_out),
    .reset(cond860_reset),
    .write_en(cond860_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire860 (
    .in(cond_wire860_in),
    .out(cond_wire860_out)
);
std_reg # (
    .WIDTH(1)
) cond861 (
    .clk(cond861_clk),
    .done(cond861_done),
    .in(cond861_in),
    .out(cond861_out),
    .reset(cond861_reset),
    .write_en(cond861_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire861 (
    .in(cond_wire861_in),
    .out(cond_wire861_out)
);
std_reg # (
    .WIDTH(1)
) cond862 (
    .clk(cond862_clk),
    .done(cond862_done),
    .in(cond862_in),
    .out(cond862_out),
    .reset(cond862_reset),
    .write_en(cond862_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire862 (
    .in(cond_wire862_in),
    .out(cond_wire862_out)
);
std_reg # (
    .WIDTH(1)
) cond863 (
    .clk(cond863_clk),
    .done(cond863_done),
    .in(cond863_in),
    .out(cond863_out),
    .reset(cond863_reset),
    .write_en(cond863_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire863 (
    .in(cond_wire863_in),
    .out(cond_wire863_out)
);
std_reg # (
    .WIDTH(1)
) cond864 (
    .clk(cond864_clk),
    .done(cond864_done),
    .in(cond864_in),
    .out(cond864_out),
    .reset(cond864_reset),
    .write_en(cond864_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire864 (
    .in(cond_wire864_in),
    .out(cond_wire864_out)
);
std_reg # (
    .WIDTH(1)
) cond865 (
    .clk(cond865_clk),
    .done(cond865_done),
    .in(cond865_in),
    .out(cond865_out),
    .reset(cond865_reset),
    .write_en(cond865_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire865 (
    .in(cond_wire865_in),
    .out(cond_wire865_out)
);
std_reg # (
    .WIDTH(1)
) cond866 (
    .clk(cond866_clk),
    .done(cond866_done),
    .in(cond866_in),
    .out(cond866_out),
    .reset(cond866_reset),
    .write_en(cond866_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire866 (
    .in(cond_wire866_in),
    .out(cond_wire866_out)
);
std_reg # (
    .WIDTH(1)
) cond867 (
    .clk(cond867_clk),
    .done(cond867_done),
    .in(cond867_in),
    .out(cond867_out),
    .reset(cond867_reset),
    .write_en(cond867_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire867 (
    .in(cond_wire867_in),
    .out(cond_wire867_out)
);
std_reg # (
    .WIDTH(1)
) cond868 (
    .clk(cond868_clk),
    .done(cond868_done),
    .in(cond868_in),
    .out(cond868_out),
    .reset(cond868_reset),
    .write_en(cond868_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire868 (
    .in(cond_wire868_in),
    .out(cond_wire868_out)
);
std_reg # (
    .WIDTH(1)
) cond869 (
    .clk(cond869_clk),
    .done(cond869_done),
    .in(cond869_in),
    .out(cond869_out),
    .reset(cond869_reset),
    .write_en(cond869_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire869 (
    .in(cond_wire869_in),
    .out(cond_wire869_out)
);
std_reg # (
    .WIDTH(1)
) cond870 (
    .clk(cond870_clk),
    .done(cond870_done),
    .in(cond870_in),
    .out(cond870_out),
    .reset(cond870_reset),
    .write_en(cond870_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire870 (
    .in(cond_wire870_in),
    .out(cond_wire870_out)
);
std_reg # (
    .WIDTH(1)
) cond871 (
    .clk(cond871_clk),
    .done(cond871_done),
    .in(cond871_in),
    .out(cond871_out),
    .reset(cond871_reset),
    .write_en(cond871_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire871 (
    .in(cond_wire871_in),
    .out(cond_wire871_out)
);
std_reg # (
    .WIDTH(1)
) cond872 (
    .clk(cond872_clk),
    .done(cond872_done),
    .in(cond872_in),
    .out(cond872_out),
    .reset(cond872_reset),
    .write_en(cond872_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire872 (
    .in(cond_wire872_in),
    .out(cond_wire872_out)
);
std_reg # (
    .WIDTH(1)
) cond873 (
    .clk(cond873_clk),
    .done(cond873_done),
    .in(cond873_in),
    .out(cond873_out),
    .reset(cond873_reset),
    .write_en(cond873_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire873 (
    .in(cond_wire873_in),
    .out(cond_wire873_out)
);
std_reg # (
    .WIDTH(1)
) cond874 (
    .clk(cond874_clk),
    .done(cond874_done),
    .in(cond874_in),
    .out(cond874_out),
    .reset(cond874_reset),
    .write_en(cond874_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire874 (
    .in(cond_wire874_in),
    .out(cond_wire874_out)
);
std_reg # (
    .WIDTH(1)
) cond875 (
    .clk(cond875_clk),
    .done(cond875_done),
    .in(cond875_in),
    .out(cond875_out),
    .reset(cond875_reset),
    .write_en(cond875_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire875 (
    .in(cond_wire875_in),
    .out(cond_wire875_out)
);
std_reg # (
    .WIDTH(1)
) cond876 (
    .clk(cond876_clk),
    .done(cond876_done),
    .in(cond876_in),
    .out(cond876_out),
    .reset(cond876_reset),
    .write_en(cond876_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire876 (
    .in(cond_wire876_in),
    .out(cond_wire876_out)
);
std_reg # (
    .WIDTH(1)
) cond877 (
    .clk(cond877_clk),
    .done(cond877_done),
    .in(cond877_in),
    .out(cond877_out),
    .reset(cond877_reset),
    .write_en(cond877_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire877 (
    .in(cond_wire877_in),
    .out(cond_wire877_out)
);
std_reg # (
    .WIDTH(1)
) cond878 (
    .clk(cond878_clk),
    .done(cond878_done),
    .in(cond878_in),
    .out(cond878_out),
    .reset(cond878_reset),
    .write_en(cond878_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire878 (
    .in(cond_wire878_in),
    .out(cond_wire878_out)
);
std_reg # (
    .WIDTH(1)
) cond879 (
    .clk(cond879_clk),
    .done(cond879_done),
    .in(cond879_in),
    .out(cond879_out),
    .reset(cond879_reset),
    .write_en(cond879_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire879 (
    .in(cond_wire879_in),
    .out(cond_wire879_out)
);
std_reg # (
    .WIDTH(1)
) cond880 (
    .clk(cond880_clk),
    .done(cond880_done),
    .in(cond880_in),
    .out(cond880_out),
    .reset(cond880_reset),
    .write_en(cond880_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire880 (
    .in(cond_wire880_in),
    .out(cond_wire880_out)
);
std_reg # (
    .WIDTH(1)
) cond881 (
    .clk(cond881_clk),
    .done(cond881_done),
    .in(cond881_in),
    .out(cond881_out),
    .reset(cond881_reset),
    .write_en(cond881_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire881 (
    .in(cond_wire881_in),
    .out(cond_wire881_out)
);
std_reg # (
    .WIDTH(1)
) cond882 (
    .clk(cond882_clk),
    .done(cond882_done),
    .in(cond882_in),
    .out(cond882_out),
    .reset(cond882_reset),
    .write_en(cond882_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire882 (
    .in(cond_wire882_in),
    .out(cond_wire882_out)
);
std_reg # (
    .WIDTH(1)
) cond883 (
    .clk(cond883_clk),
    .done(cond883_done),
    .in(cond883_in),
    .out(cond883_out),
    .reset(cond883_reset),
    .write_en(cond883_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire883 (
    .in(cond_wire883_in),
    .out(cond_wire883_out)
);
std_reg # (
    .WIDTH(1)
) cond884 (
    .clk(cond884_clk),
    .done(cond884_done),
    .in(cond884_in),
    .out(cond884_out),
    .reset(cond884_reset),
    .write_en(cond884_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire884 (
    .in(cond_wire884_in),
    .out(cond_wire884_out)
);
std_reg # (
    .WIDTH(1)
) cond885 (
    .clk(cond885_clk),
    .done(cond885_done),
    .in(cond885_in),
    .out(cond885_out),
    .reset(cond885_reset),
    .write_en(cond885_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire885 (
    .in(cond_wire885_in),
    .out(cond_wire885_out)
);
std_reg # (
    .WIDTH(1)
) cond886 (
    .clk(cond886_clk),
    .done(cond886_done),
    .in(cond886_in),
    .out(cond886_out),
    .reset(cond886_reset),
    .write_en(cond886_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire886 (
    .in(cond_wire886_in),
    .out(cond_wire886_out)
);
std_reg # (
    .WIDTH(1)
) cond887 (
    .clk(cond887_clk),
    .done(cond887_done),
    .in(cond887_in),
    .out(cond887_out),
    .reset(cond887_reset),
    .write_en(cond887_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire887 (
    .in(cond_wire887_in),
    .out(cond_wire887_out)
);
std_reg # (
    .WIDTH(1)
) cond888 (
    .clk(cond888_clk),
    .done(cond888_done),
    .in(cond888_in),
    .out(cond888_out),
    .reset(cond888_reset),
    .write_en(cond888_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire888 (
    .in(cond_wire888_in),
    .out(cond_wire888_out)
);
std_reg # (
    .WIDTH(1)
) cond889 (
    .clk(cond889_clk),
    .done(cond889_done),
    .in(cond889_in),
    .out(cond889_out),
    .reset(cond889_reset),
    .write_en(cond889_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire889 (
    .in(cond_wire889_in),
    .out(cond_wire889_out)
);
std_reg # (
    .WIDTH(1)
) cond890 (
    .clk(cond890_clk),
    .done(cond890_done),
    .in(cond890_in),
    .out(cond890_out),
    .reset(cond890_reset),
    .write_en(cond890_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire890 (
    .in(cond_wire890_in),
    .out(cond_wire890_out)
);
std_reg # (
    .WIDTH(1)
) cond891 (
    .clk(cond891_clk),
    .done(cond891_done),
    .in(cond891_in),
    .out(cond891_out),
    .reset(cond891_reset),
    .write_en(cond891_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire891 (
    .in(cond_wire891_in),
    .out(cond_wire891_out)
);
std_reg # (
    .WIDTH(1)
) cond892 (
    .clk(cond892_clk),
    .done(cond892_done),
    .in(cond892_in),
    .out(cond892_out),
    .reset(cond892_reset),
    .write_en(cond892_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire892 (
    .in(cond_wire892_in),
    .out(cond_wire892_out)
);
std_reg # (
    .WIDTH(1)
) cond893 (
    .clk(cond893_clk),
    .done(cond893_done),
    .in(cond893_in),
    .out(cond893_out),
    .reset(cond893_reset),
    .write_en(cond893_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire893 (
    .in(cond_wire893_in),
    .out(cond_wire893_out)
);
std_reg # (
    .WIDTH(1)
) cond894 (
    .clk(cond894_clk),
    .done(cond894_done),
    .in(cond894_in),
    .out(cond894_out),
    .reset(cond894_reset),
    .write_en(cond894_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire894 (
    .in(cond_wire894_in),
    .out(cond_wire894_out)
);
std_reg # (
    .WIDTH(1)
) cond895 (
    .clk(cond895_clk),
    .done(cond895_done),
    .in(cond895_in),
    .out(cond895_out),
    .reset(cond895_reset),
    .write_en(cond895_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire895 (
    .in(cond_wire895_in),
    .out(cond_wire895_out)
);
std_reg # (
    .WIDTH(1)
) cond896 (
    .clk(cond896_clk),
    .done(cond896_done),
    .in(cond896_in),
    .out(cond896_out),
    .reset(cond896_reset),
    .write_en(cond896_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire896 (
    .in(cond_wire896_in),
    .out(cond_wire896_out)
);
std_reg # (
    .WIDTH(1)
) cond897 (
    .clk(cond897_clk),
    .done(cond897_done),
    .in(cond897_in),
    .out(cond897_out),
    .reset(cond897_reset),
    .write_en(cond897_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire897 (
    .in(cond_wire897_in),
    .out(cond_wire897_out)
);
std_reg # (
    .WIDTH(1)
) cond898 (
    .clk(cond898_clk),
    .done(cond898_done),
    .in(cond898_in),
    .out(cond898_out),
    .reset(cond898_reset),
    .write_en(cond898_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire898 (
    .in(cond_wire898_in),
    .out(cond_wire898_out)
);
std_reg # (
    .WIDTH(1)
) cond899 (
    .clk(cond899_clk),
    .done(cond899_done),
    .in(cond899_in),
    .out(cond899_out),
    .reset(cond899_reset),
    .write_en(cond899_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire899 (
    .in(cond_wire899_in),
    .out(cond_wire899_out)
);
std_reg # (
    .WIDTH(1)
) cond900 (
    .clk(cond900_clk),
    .done(cond900_done),
    .in(cond900_in),
    .out(cond900_out),
    .reset(cond900_reset),
    .write_en(cond900_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire900 (
    .in(cond_wire900_in),
    .out(cond_wire900_out)
);
std_reg # (
    .WIDTH(1)
) cond901 (
    .clk(cond901_clk),
    .done(cond901_done),
    .in(cond901_in),
    .out(cond901_out),
    .reset(cond901_reset),
    .write_en(cond901_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire901 (
    .in(cond_wire901_in),
    .out(cond_wire901_out)
);
std_reg # (
    .WIDTH(1)
) cond902 (
    .clk(cond902_clk),
    .done(cond902_done),
    .in(cond902_in),
    .out(cond902_out),
    .reset(cond902_reset),
    .write_en(cond902_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire902 (
    .in(cond_wire902_in),
    .out(cond_wire902_out)
);
std_reg # (
    .WIDTH(1)
) cond903 (
    .clk(cond903_clk),
    .done(cond903_done),
    .in(cond903_in),
    .out(cond903_out),
    .reset(cond903_reset),
    .write_en(cond903_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire903 (
    .in(cond_wire903_in),
    .out(cond_wire903_out)
);
std_reg # (
    .WIDTH(1)
) cond904 (
    .clk(cond904_clk),
    .done(cond904_done),
    .in(cond904_in),
    .out(cond904_out),
    .reset(cond904_reset),
    .write_en(cond904_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire904 (
    .in(cond_wire904_in),
    .out(cond_wire904_out)
);
std_reg # (
    .WIDTH(1)
) cond905 (
    .clk(cond905_clk),
    .done(cond905_done),
    .in(cond905_in),
    .out(cond905_out),
    .reset(cond905_reset),
    .write_en(cond905_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire905 (
    .in(cond_wire905_in),
    .out(cond_wire905_out)
);
std_reg # (
    .WIDTH(1)
) cond906 (
    .clk(cond906_clk),
    .done(cond906_done),
    .in(cond906_in),
    .out(cond906_out),
    .reset(cond906_reset),
    .write_en(cond906_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire906 (
    .in(cond_wire906_in),
    .out(cond_wire906_out)
);
std_reg # (
    .WIDTH(1)
) cond907 (
    .clk(cond907_clk),
    .done(cond907_done),
    .in(cond907_in),
    .out(cond907_out),
    .reset(cond907_reset),
    .write_en(cond907_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire907 (
    .in(cond_wire907_in),
    .out(cond_wire907_out)
);
std_reg # (
    .WIDTH(1)
) cond908 (
    .clk(cond908_clk),
    .done(cond908_done),
    .in(cond908_in),
    .out(cond908_out),
    .reset(cond908_reset),
    .write_en(cond908_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire908 (
    .in(cond_wire908_in),
    .out(cond_wire908_out)
);
std_reg # (
    .WIDTH(1)
) cond909 (
    .clk(cond909_clk),
    .done(cond909_done),
    .in(cond909_in),
    .out(cond909_out),
    .reset(cond909_reset),
    .write_en(cond909_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire909 (
    .in(cond_wire909_in),
    .out(cond_wire909_out)
);
std_reg # (
    .WIDTH(1)
) cond910 (
    .clk(cond910_clk),
    .done(cond910_done),
    .in(cond910_in),
    .out(cond910_out),
    .reset(cond910_reset),
    .write_en(cond910_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire910 (
    .in(cond_wire910_in),
    .out(cond_wire910_out)
);
std_reg # (
    .WIDTH(1)
) cond911 (
    .clk(cond911_clk),
    .done(cond911_done),
    .in(cond911_in),
    .out(cond911_out),
    .reset(cond911_reset),
    .write_en(cond911_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire911 (
    .in(cond_wire911_in),
    .out(cond_wire911_out)
);
std_reg # (
    .WIDTH(1)
) cond912 (
    .clk(cond912_clk),
    .done(cond912_done),
    .in(cond912_in),
    .out(cond912_out),
    .reset(cond912_reset),
    .write_en(cond912_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire912 (
    .in(cond_wire912_in),
    .out(cond_wire912_out)
);
std_reg # (
    .WIDTH(1)
) cond913 (
    .clk(cond913_clk),
    .done(cond913_done),
    .in(cond913_in),
    .out(cond913_out),
    .reset(cond913_reset),
    .write_en(cond913_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire913 (
    .in(cond_wire913_in),
    .out(cond_wire913_out)
);
std_reg # (
    .WIDTH(1)
) cond914 (
    .clk(cond914_clk),
    .done(cond914_done),
    .in(cond914_in),
    .out(cond914_out),
    .reset(cond914_reset),
    .write_en(cond914_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire914 (
    .in(cond_wire914_in),
    .out(cond_wire914_out)
);
std_reg # (
    .WIDTH(1)
) cond915 (
    .clk(cond915_clk),
    .done(cond915_done),
    .in(cond915_in),
    .out(cond915_out),
    .reset(cond915_reset),
    .write_en(cond915_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire915 (
    .in(cond_wire915_in),
    .out(cond_wire915_out)
);
std_reg # (
    .WIDTH(1)
) cond916 (
    .clk(cond916_clk),
    .done(cond916_done),
    .in(cond916_in),
    .out(cond916_out),
    .reset(cond916_reset),
    .write_en(cond916_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire916 (
    .in(cond_wire916_in),
    .out(cond_wire916_out)
);
std_reg # (
    .WIDTH(1)
) cond917 (
    .clk(cond917_clk),
    .done(cond917_done),
    .in(cond917_in),
    .out(cond917_out),
    .reset(cond917_reset),
    .write_en(cond917_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire917 (
    .in(cond_wire917_in),
    .out(cond_wire917_out)
);
std_reg # (
    .WIDTH(1)
) cond918 (
    .clk(cond918_clk),
    .done(cond918_done),
    .in(cond918_in),
    .out(cond918_out),
    .reset(cond918_reset),
    .write_en(cond918_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire918 (
    .in(cond_wire918_in),
    .out(cond_wire918_out)
);
std_reg # (
    .WIDTH(1)
) cond919 (
    .clk(cond919_clk),
    .done(cond919_done),
    .in(cond919_in),
    .out(cond919_out),
    .reset(cond919_reset),
    .write_en(cond919_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire919 (
    .in(cond_wire919_in),
    .out(cond_wire919_out)
);
std_reg # (
    .WIDTH(1)
) cond920 (
    .clk(cond920_clk),
    .done(cond920_done),
    .in(cond920_in),
    .out(cond920_out),
    .reset(cond920_reset),
    .write_en(cond920_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire920 (
    .in(cond_wire920_in),
    .out(cond_wire920_out)
);
std_reg # (
    .WIDTH(1)
) cond921 (
    .clk(cond921_clk),
    .done(cond921_done),
    .in(cond921_in),
    .out(cond921_out),
    .reset(cond921_reset),
    .write_en(cond921_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire921 (
    .in(cond_wire921_in),
    .out(cond_wire921_out)
);
std_reg # (
    .WIDTH(1)
) cond922 (
    .clk(cond922_clk),
    .done(cond922_done),
    .in(cond922_in),
    .out(cond922_out),
    .reset(cond922_reset),
    .write_en(cond922_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire922 (
    .in(cond_wire922_in),
    .out(cond_wire922_out)
);
std_reg # (
    .WIDTH(1)
) cond923 (
    .clk(cond923_clk),
    .done(cond923_done),
    .in(cond923_in),
    .out(cond923_out),
    .reset(cond923_reset),
    .write_en(cond923_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire923 (
    .in(cond_wire923_in),
    .out(cond_wire923_out)
);
std_reg # (
    .WIDTH(1)
) cond924 (
    .clk(cond924_clk),
    .done(cond924_done),
    .in(cond924_in),
    .out(cond924_out),
    .reset(cond924_reset),
    .write_en(cond924_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire924 (
    .in(cond_wire924_in),
    .out(cond_wire924_out)
);
std_reg # (
    .WIDTH(1)
) cond925 (
    .clk(cond925_clk),
    .done(cond925_done),
    .in(cond925_in),
    .out(cond925_out),
    .reset(cond925_reset),
    .write_en(cond925_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire925 (
    .in(cond_wire925_in),
    .out(cond_wire925_out)
);
std_reg # (
    .WIDTH(1)
) cond926 (
    .clk(cond926_clk),
    .done(cond926_done),
    .in(cond926_in),
    .out(cond926_out),
    .reset(cond926_reset),
    .write_en(cond926_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire926 (
    .in(cond_wire926_in),
    .out(cond_wire926_out)
);
std_reg # (
    .WIDTH(1)
) cond927 (
    .clk(cond927_clk),
    .done(cond927_done),
    .in(cond927_in),
    .out(cond927_out),
    .reset(cond927_reset),
    .write_en(cond927_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire927 (
    .in(cond_wire927_in),
    .out(cond_wire927_out)
);
std_reg # (
    .WIDTH(1)
) cond928 (
    .clk(cond928_clk),
    .done(cond928_done),
    .in(cond928_in),
    .out(cond928_out),
    .reset(cond928_reset),
    .write_en(cond928_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire928 (
    .in(cond_wire928_in),
    .out(cond_wire928_out)
);
std_reg # (
    .WIDTH(1)
) cond929 (
    .clk(cond929_clk),
    .done(cond929_done),
    .in(cond929_in),
    .out(cond929_out),
    .reset(cond929_reset),
    .write_en(cond929_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire929 (
    .in(cond_wire929_in),
    .out(cond_wire929_out)
);
std_reg # (
    .WIDTH(1)
) cond930 (
    .clk(cond930_clk),
    .done(cond930_done),
    .in(cond930_in),
    .out(cond930_out),
    .reset(cond930_reset),
    .write_en(cond930_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire930 (
    .in(cond_wire930_in),
    .out(cond_wire930_out)
);
std_reg # (
    .WIDTH(1)
) cond931 (
    .clk(cond931_clk),
    .done(cond931_done),
    .in(cond931_in),
    .out(cond931_out),
    .reset(cond931_reset),
    .write_en(cond931_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire931 (
    .in(cond_wire931_in),
    .out(cond_wire931_out)
);
std_reg # (
    .WIDTH(1)
) cond932 (
    .clk(cond932_clk),
    .done(cond932_done),
    .in(cond932_in),
    .out(cond932_out),
    .reset(cond932_reset),
    .write_en(cond932_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire932 (
    .in(cond_wire932_in),
    .out(cond_wire932_out)
);
std_reg # (
    .WIDTH(1)
) cond933 (
    .clk(cond933_clk),
    .done(cond933_done),
    .in(cond933_in),
    .out(cond933_out),
    .reset(cond933_reset),
    .write_en(cond933_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire933 (
    .in(cond_wire933_in),
    .out(cond_wire933_out)
);
std_reg # (
    .WIDTH(1)
) cond934 (
    .clk(cond934_clk),
    .done(cond934_done),
    .in(cond934_in),
    .out(cond934_out),
    .reset(cond934_reset),
    .write_en(cond934_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire934 (
    .in(cond_wire934_in),
    .out(cond_wire934_out)
);
std_reg # (
    .WIDTH(1)
) cond935 (
    .clk(cond935_clk),
    .done(cond935_done),
    .in(cond935_in),
    .out(cond935_out),
    .reset(cond935_reset),
    .write_en(cond935_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire935 (
    .in(cond_wire935_in),
    .out(cond_wire935_out)
);
std_reg # (
    .WIDTH(1)
) cond936 (
    .clk(cond936_clk),
    .done(cond936_done),
    .in(cond936_in),
    .out(cond936_out),
    .reset(cond936_reset),
    .write_en(cond936_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire936 (
    .in(cond_wire936_in),
    .out(cond_wire936_out)
);
std_reg # (
    .WIDTH(1)
) cond937 (
    .clk(cond937_clk),
    .done(cond937_done),
    .in(cond937_in),
    .out(cond937_out),
    .reset(cond937_reset),
    .write_en(cond937_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire937 (
    .in(cond_wire937_in),
    .out(cond_wire937_out)
);
std_reg # (
    .WIDTH(1)
) cond938 (
    .clk(cond938_clk),
    .done(cond938_done),
    .in(cond938_in),
    .out(cond938_out),
    .reset(cond938_reset),
    .write_en(cond938_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire938 (
    .in(cond_wire938_in),
    .out(cond_wire938_out)
);
std_reg # (
    .WIDTH(1)
) cond939 (
    .clk(cond939_clk),
    .done(cond939_done),
    .in(cond939_in),
    .out(cond939_out),
    .reset(cond939_reset),
    .write_en(cond939_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire939 (
    .in(cond_wire939_in),
    .out(cond_wire939_out)
);
std_reg # (
    .WIDTH(1)
) cond940 (
    .clk(cond940_clk),
    .done(cond940_done),
    .in(cond940_in),
    .out(cond940_out),
    .reset(cond940_reset),
    .write_en(cond940_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire940 (
    .in(cond_wire940_in),
    .out(cond_wire940_out)
);
std_reg # (
    .WIDTH(1)
) cond941 (
    .clk(cond941_clk),
    .done(cond941_done),
    .in(cond941_in),
    .out(cond941_out),
    .reset(cond941_reset),
    .write_en(cond941_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire941 (
    .in(cond_wire941_in),
    .out(cond_wire941_out)
);
std_reg # (
    .WIDTH(1)
) cond942 (
    .clk(cond942_clk),
    .done(cond942_done),
    .in(cond942_in),
    .out(cond942_out),
    .reset(cond942_reset),
    .write_en(cond942_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire942 (
    .in(cond_wire942_in),
    .out(cond_wire942_out)
);
std_reg # (
    .WIDTH(1)
) cond943 (
    .clk(cond943_clk),
    .done(cond943_done),
    .in(cond943_in),
    .out(cond943_out),
    .reset(cond943_reset),
    .write_en(cond943_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire943 (
    .in(cond_wire943_in),
    .out(cond_wire943_out)
);
std_reg # (
    .WIDTH(1)
) cond944 (
    .clk(cond944_clk),
    .done(cond944_done),
    .in(cond944_in),
    .out(cond944_out),
    .reset(cond944_reset),
    .write_en(cond944_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire944 (
    .in(cond_wire944_in),
    .out(cond_wire944_out)
);
std_reg # (
    .WIDTH(1)
) cond945 (
    .clk(cond945_clk),
    .done(cond945_done),
    .in(cond945_in),
    .out(cond945_out),
    .reset(cond945_reset),
    .write_en(cond945_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire945 (
    .in(cond_wire945_in),
    .out(cond_wire945_out)
);
std_reg # (
    .WIDTH(1)
) cond946 (
    .clk(cond946_clk),
    .done(cond946_done),
    .in(cond946_in),
    .out(cond946_out),
    .reset(cond946_reset),
    .write_en(cond946_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire946 (
    .in(cond_wire946_in),
    .out(cond_wire946_out)
);
std_reg # (
    .WIDTH(1)
) cond947 (
    .clk(cond947_clk),
    .done(cond947_done),
    .in(cond947_in),
    .out(cond947_out),
    .reset(cond947_reset),
    .write_en(cond947_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire947 (
    .in(cond_wire947_in),
    .out(cond_wire947_out)
);
std_reg # (
    .WIDTH(1)
) cond948 (
    .clk(cond948_clk),
    .done(cond948_done),
    .in(cond948_in),
    .out(cond948_out),
    .reset(cond948_reset),
    .write_en(cond948_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire948 (
    .in(cond_wire948_in),
    .out(cond_wire948_out)
);
std_reg # (
    .WIDTH(1)
) cond949 (
    .clk(cond949_clk),
    .done(cond949_done),
    .in(cond949_in),
    .out(cond949_out),
    .reset(cond949_reset),
    .write_en(cond949_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire949 (
    .in(cond_wire949_in),
    .out(cond_wire949_out)
);
std_reg # (
    .WIDTH(1)
) cond950 (
    .clk(cond950_clk),
    .done(cond950_done),
    .in(cond950_in),
    .out(cond950_out),
    .reset(cond950_reset),
    .write_en(cond950_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire950 (
    .in(cond_wire950_in),
    .out(cond_wire950_out)
);
std_reg # (
    .WIDTH(1)
) cond951 (
    .clk(cond951_clk),
    .done(cond951_done),
    .in(cond951_in),
    .out(cond951_out),
    .reset(cond951_reset),
    .write_en(cond951_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire951 (
    .in(cond_wire951_in),
    .out(cond_wire951_out)
);
std_reg # (
    .WIDTH(1)
) cond952 (
    .clk(cond952_clk),
    .done(cond952_done),
    .in(cond952_in),
    .out(cond952_out),
    .reset(cond952_reset),
    .write_en(cond952_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire952 (
    .in(cond_wire952_in),
    .out(cond_wire952_out)
);
std_reg # (
    .WIDTH(1)
) cond953 (
    .clk(cond953_clk),
    .done(cond953_done),
    .in(cond953_in),
    .out(cond953_out),
    .reset(cond953_reset),
    .write_en(cond953_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire953 (
    .in(cond_wire953_in),
    .out(cond_wire953_out)
);
std_reg # (
    .WIDTH(1)
) cond954 (
    .clk(cond954_clk),
    .done(cond954_done),
    .in(cond954_in),
    .out(cond954_out),
    .reset(cond954_reset),
    .write_en(cond954_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire954 (
    .in(cond_wire954_in),
    .out(cond_wire954_out)
);
std_reg # (
    .WIDTH(1)
) cond955 (
    .clk(cond955_clk),
    .done(cond955_done),
    .in(cond955_in),
    .out(cond955_out),
    .reset(cond955_reset),
    .write_en(cond955_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire955 (
    .in(cond_wire955_in),
    .out(cond_wire955_out)
);
std_reg # (
    .WIDTH(1)
) cond956 (
    .clk(cond956_clk),
    .done(cond956_done),
    .in(cond956_in),
    .out(cond956_out),
    .reset(cond956_reset),
    .write_en(cond956_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire956 (
    .in(cond_wire956_in),
    .out(cond_wire956_out)
);
std_reg # (
    .WIDTH(1)
) cond957 (
    .clk(cond957_clk),
    .done(cond957_done),
    .in(cond957_in),
    .out(cond957_out),
    .reset(cond957_reset),
    .write_en(cond957_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire957 (
    .in(cond_wire957_in),
    .out(cond_wire957_out)
);
std_reg # (
    .WIDTH(1)
) cond958 (
    .clk(cond958_clk),
    .done(cond958_done),
    .in(cond958_in),
    .out(cond958_out),
    .reset(cond958_reset),
    .write_en(cond958_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire958 (
    .in(cond_wire958_in),
    .out(cond_wire958_out)
);
std_reg # (
    .WIDTH(1)
) cond959 (
    .clk(cond959_clk),
    .done(cond959_done),
    .in(cond959_in),
    .out(cond959_out),
    .reset(cond959_reset),
    .write_en(cond959_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire959 (
    .in(cond_wire959_in),
    .out(cond_wire959_out)
);
std_reg # (
    .WIDTH(1)
) cond960 (
    .clk(cond960_clk),
    .done(cond960_done),
    .in(cond960_in),
    .out(cond960_out),
    .reset(cond960_reset),
    .write_en(cond960_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire960 (
    .in(cond_wire960_in),
    .out(cond_wire960_out)
);
std_reg # (
    .WIDTH(1)
) cond961 (
    .clk(cond961_clk),
    .done(cond961_done),
    .in(cond961_in),
    .out(cond961_out),
    .reset(cond961_reset),
    .write_en(cond961_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire961 (
    .in(cond_wire961_in),
    .out(cond_wire961_out)
);
std_reg # (
    .WIDTH(1)
) cond962 (
    .clk(cond962_clk),
    .done(cond962_done),
    .in(cond962_in),
    .out(cond962_out),
    .reset(cond962_reset),
    .write_en(cond962_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire962 (
    .in(cond_wire962_in),
    .out(cond_wire962_out)
);
std_reg # (
    .WIDTH(1)
) cond963 (
    .clk(cond963_clk),
    .done(cond963_done),
    .in(cond963_in),
    .out(cond963_out),
    .reset(cond963_reset),
    .write_en(cond963_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire963 (
    .in(cond_wire963_in),
    .out(cond_wire963_out)
);
std_reg # (
    .WIDTH(1)
) cond964 (
    .clk(cond964_clk),
    .done(cond964_done),
    .in(cond964_in),
    .out(cond964_out),
    .reset(cond964_reset),
    .write_en(cond964_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire964 (
    .in(cond_wire964_in),
    .out(cond_wire964_out)
);
std_reg # (
    .WIDTH(1)
) cond965 (
    .clk(cond965_clk),
    .done(cond965_done),
    .in(cond965_in),
    .out(cond965_out),
    .reset(cond965_reset),
    .write_en(cond965_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire965 (
    .in(cond_wire965_in),
    .out(cond_wire965_out)
);
std_reg # (
    .WIDTH(1)
) cond966 (
    .clk(cond966_clk),
    .done(cond966_done),
    .in(cond966_in),
    .out(cond966_out),
    .reset(cond966_reset),
    .write_en(cond966_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire966 (
    .in(cond_wire966_in),
    .out(cond_wire966_out)
);
std_reg # (
    .WIDTH(1)
) cond967 (
    .clk(cond967_clk),
    .done(cond967_done),
    .in(cond967_in),
    .out(cond967_out),
    .reset(cond967_reset),
    .write_en(cond967_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire967 (
    .in(cond_wire967_in),
    .out(cond_wire967_out)
);
std_reg # (
    .WIDTH(1)
) cond968 (
    .clk(cond968_clk),
    .done(cond968_done),
    .in(cond968_in),
    .out(cond968_out),
    .reset(cond968_reset),
    .write_en(cond968_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire968 (
    .in(cond_wire968_in),
    .out(cond_wire968_out)
);
std_reg # (
    .WIDTH(1)
) cond969 (
    .clk(cond969_clk),
    .done(cond969_done),
    .in(cond969_in),
    .out(cond969_out),
    .reset(cond969_reset),
    .write_en(cond969_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire969 (
    .in(cond_wire969_in),
    .out(cond_wire969_out)
);
std_reg # (
    .WIDTH(1)
) cond970 (
    .clk(cond970_clk),
    .done(cond970_done),
    .in(cond970_in),
    .out(cond970_out),
    .reset(cond970_reset),
    .write_en(cond970_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire970 (
    .in(cond_wire970_in),
    .out(cond_wire970_out)
);
std_reg # (
    .WIDTH(1)
) cond971 (
    .clk(cond971_clk),
    .done(cond971_done),
    .in(cond971_in),
    .out(cond971_out),
    .reset(cond971_reset),
    .write_en(cond971_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire971 (
    .in(cond_wire971_in),
    .out(cond_wire971_out)
);
std_reg # (
    .WIDTH(1)
) cond972 (
    .clk(cond972_clk),
    .done(cond972_done),
    .in(cond972_in),
    .out(cond972_out),
    .reset(cond972_reset),
    .write_en(cond972_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire972 (
    .in(cond_wire972_in),
    .out(cond_wire972_out)
);
std_reg # (
    .WIDTH(1)
) cond973 (
    .clk(cond973_clk),
    .done(cond973_done),
    .in(cond973_in),
    .out(cond973_out),
    .reset(cond973_reset),
    .write_en(cond973_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire973 (
    .in(cond_wire973_in),
    .out(cond_wire973_out)
);
std_reg # (
    .WIDTH(1)
) cond974 (
    .clk(cond974_clk),
    .done(cond974_done),
    .in(cond974_in),
    .out(cond974_out),
    .reset(cond974_reset),
    .write_en(cond974_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire974 (
    .in(cond_wire974_in),
    .out(cond_wire974_out)
);
std_reg # (
    .WIDTH(1)
) cond975 (
    .clk(cond975_clk),
    .done(cond975_done),
    .in(cond975_in),
    .out(cond975_out),
    .reset(cond975_reset),
    .write_en(cond975_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire975 (
    .in(cond_wire975_in),
    .out(cond_wire975_out)
);
std_reg # (
    .WIDTH(1)
) cond976 (
    .clk(cond976_clk),
    .done(cond976_done),
    .in(cond976_in),
    .out(cond976_out),
    .reset(cond976_reset),
    .write_en(cond976_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire976 (
    .in(cond_wire976_in),
    .out(cond_wire976_out)
);
std_reg # (
    .WIDTH(1)
) cond977 (
    .clk(cond977_clk),
    .done(cond977_done),
    .in(cond977_in),
    .out(cond977_out),
    .reset(cond977_reset),
    .write_en(cond977_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire977 (
    .in(cond_wire977_in),
    .out(cond_wire977_out)
);
std_reg # (
    .WIDTH(1)
) cond978 (
    .clk(cond978_clk),
    .done(cond978_done),
    .in(cond978_in),
    .out(cond978_out),
    .reset(cond978_reset),
    .write_en(cond978_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire978 (
    .in(cond_wire978_in),
    .out(cond_wire978_out)
);
std_reg # (
    .WIDTH(1)
) cond979 (
    .clk(cond979_clk),
    .done(cond979_done),
    .in(cond979_in),
    .out(cond979_out),
    .reset(cond979_reset),
    .write_en(cond979_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire979 (
    .in(cond_wire979_in),
    .out(cond_wire979_out)
);
std_reg # (
    .WIDTH(1)
) cond980 (
    .clk(cond980_clk),
    .done(cond980_done),
    .in(cond980_in),
    .out(cond980_out),
    .reset(cond980_reset),
    .write_en(cond980_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire980 (
    .in(cond_wire980_in),
    .out(cond_wire980_out)
);
std_reg # (
    .WIDTH(1)
) cond981 (
    .clk(cond981_clk),
    .done(cond981_done),
    .in(cond981_in),
    .out(cond981_out),
    .reset(cond981_reset),
    .write_en(cond981_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire981 (
    .in(cond_wire981_in),
    .out(cond_wire981_out)
);
std_reg # (
    .WIDTH(1)
) cond982 (
    .clk(cond982_clk),
    .done(cond982_done),
    .in(cond982_in),
    .out(cond982_out),
    .reset(cond982_reset),
    .write_en(cond982_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire982 (
    .in(cond_wire982_in),
    .out(cond_wire982_out)
);
std_reg # (
    .WIDTH(1)
) cond983 (
    .clk(cond983_clk),
    .done(cond983_done),
    .in(cond983_in),
    .out(cond983_out),
    .reset(cond983_reset),
    .write_en(cond983_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire983 (
    .in(cond_wire983_in),
    .out(cond_wire983_out)
);
std_reg # (
    .WIDTH(1)
) cond984 (
    .clk(cond984_clk),
    .done(cond984_done),
    .in(cond984_in),
    .out(cond984_out),
    .reset(cond984_reset),
    .write_en(cond984_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire984 (
    .in(cond_wire984_in),
    .out(cond_wire984_out)
);
std_reg # (
    .WIDTH(1)
) cond985 (
    .clk(cond985_clk),
    .done(cond985_done),
    .in(cond985_in),
    .out(cond985_out),
    .reset(cond985_reset),
    .write_en(cond985_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire985 (
    .in(cond_wire985_in),
    .out(cond_wire985_out)
);
std_reg # (
    .WIDTH(1)
) cond986 (
    .clk(cond986_clk),
    .done(cond986_done),
    .in(cond986_in),
    .out(cond986_out),
    .reset(cond986_reset),
    .write_en(cond986_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire986 (
    .in(cond_wire986_in),
    .out(cond_wire986_out)
);
std_reg # (
    .WIDTH(1)
) cond987 (
    .clk(cond987_clk),
    .done(cond987_done),
    .in(cond987_in),
    .out(cond987_out),
    .reset(cond987_reset),
    .write_en(cond987_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire987 (
    .in(cond_wire987_in),
    .out(cond_wire987_out)
);
std_reg # (
    .WIDTH(1)
) cond988 (
    .clk(cond988_clk),
    .done(cond988_done),
    .in(cond988_in),
    .out(cond988_out),
    .reset(cond988_reset),
    .write_en(cond988_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire988 (
    .in(cond_wire988_in),
    .out(cond_wire988_out)
);
std_reg # (
    .WIDTH(1)
) cond989 (
    .clk(cond989_clk),
    .done(cond989_done),
    .in(cond989_in),
    .out(cond989_out),
    .reset(cond989_reset),
    .write_en(cond989_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire989 (
    .in(cond_wire989_in),
    .out(cond_wire989_out)
);
std_reg # (
    .WIDTH(1)
) cond990 (
    .clk(cond990_clk),
    .done(cond990_done),
    .in(cond990_in),
    .out(cond990_out),
    .reset(cond990_reset),
    .write_en(cond990_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire990 (
    .in(cond_wire990_in),
    .out(cond_wire990_out)
);
std_reg # (
    .WIDTH(1)
) cond991 (
    .clk(cond991_clk),
    .done(cond991_done),
    .in(cond991_in),
    .out(cond991_out),
    .reset(cond991_reset),
    .write_en(cond991_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire991 (
    .in(cond_wire991_in),
    .out(cond_wire991_out)
);
std_reg # (
    .WIDTH(1)
) cond992 (
    .clk(cond992_clk),
    .done(cond992_done),
    .in(cond992_in),
    .out(cond992_out),
    .reset(cond992_reset),
    .write_en(cond992_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire992 (
    .in(cond_wire992_in),
    .out(cond_wire992_out)
);
std_reg # (
    .WIDTH(1)
) cond993 (
    .clk(cond993_clk),
    .done(cond993_done),
    .in(cond993_in),
    .out(cond993_out),
    .reset(cond993_reset),
    .write_en(cond993_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire993 (
    .in(cond_wire993_in),
    .out(cond_wire993_out)
);
std_reg # (
    .WIDTH(1)
) cond994 (
    .clk(cond994_clk),
    .done(cond994_done),
    .in(cond994_in),
    .out(cond994_out),
    .reset(cond994_reset),
    .write_en(cond994_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire994 (
    .in(cond_wire994_in),
    .out(cond_wire994_out)
);
std_reg # (
    .WIDTH(1)
) cond995 (
    .clk(cond995_clk),
    .done(cond995_done),
    .in(cond995_in),
    .out(cond995_out),
    .reset(cond995_reset),
    .write_en(cond995_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire995 (
    .in(cond_wire995_in),
    .out(cond_wire995_out)
);
std_reg # (
    .WIDTH(1)
) cond996 (
    .clk(cond996_clk),
    .done(cond996_done),
    .in(cond996_in),
    .out(cond996_out),
    .reset(cond996_reset),
    .write_en(cond996_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire996 (
    .in(cond_wire996_in),
    .out(cond_wire996_out)
);
std_reg # (
    .WIDTH(1)
) cond997 (
    .clk(cond997_clk),
    .done(cond997_done),
    .in(cond997_in),
    .out(cond997_out),
    .reset(cond997_reset),
    .write_en(cond997_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire997 (
    .in(cond_wire997_in),
    .out(cond_wire997_out)
);
std_reg # (
    .WIDTH(1)
) cond998 (
    .clk(cond998_clk),
    .done(cond998_done),
    .in(cond998_in),
    .out(cond998_out),
    .reset(cond998_reset),
    .write_en(cond998_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire998 (
    .in(cond_wire998_in),
    .out(cond_wire998_out)
);
std_reg # (
    .WIDTH(1)
) cond999 (
    .clk(cond999_clk),
    .done(cond999_done),
    .in(cond999_in),
    .out(cond999_out),
    .reset(cond999_reset),
    .write_en(cond999_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire999 (
    .in(cond_wire999_in),
    .out(cond_wire999_out)
);
std_reg # (
    .WIDTH(1)
) cond1000 (
    .clk(cond1000_clk),
    .done(cond1000_done),
    .in(cond1000_in),
    .out(cond1000_out),
    .reset(cond1000_reset),
    .write_en(cond1000_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1000 (
    .in(cond_wire1000_in),
    .out(cond_wire1000_out)
);
std_reg # (
    .WIDTH(1)
) cond1001 (
    .clk(cond1001_clk),
    .done(cond1001_done),
    .in(cond1001_in),
    .out(cond1001_out),
    .reset(cond1001_reset),
    .write_en(cond1001_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1001 (
    .in(cond_wire1001_in),
    .out(cond_wire1001_out)
);
std_reg # (
    .WIDTH(1)
) cond1002 (
    .clk(cond1002_clk),
    .done(cond1002_done),
    .in(cond1002_in),
    .out(cond1002_out),
    .reset(cond1002_reset),
    .write_en(cond1002_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1002 (
    .in(cond_wire1002_in),
    .out(cond_wire1002_out)
);
std_reg # (
    .WIDTH(1)
) cond1003 (
    .clk(cond1003_clk),
    .done(cond1003_done),
    .in(cond1003_in),
    .out(cond1003_out),
    .reset(cond1003_reset),
    .write_en(cond1003_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1003 (
    .in(cond_wire1003_in),
    .out(cond_wire1003_out)
);
std_reg # (
    .WIDTH(1)
) cond1004 (
    .clk(cond1004_clk),
    .done(cond1004_done),
    .in(cond1004_in),
    .out(cond1004_out),
    .reset(cond1004_reset),
    .write_en(cond1004_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1004 (
    .in(cond_wire1004_in),
    .out(cond_wire1004_out)
);
std_reg # (
    .WIDTH(1)
) cond1005 (
    .clk(cond1005_clk),
    .done(cond1005_done),
    .in(cond1005_in),
    .out(cond1005_out),
    .reset(cond1005_reset),
    .write_en(cond1005_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1005 (
    .in(cond_wire1005_in),
    .out(cond_wire1005_out)
);
std_reg # (
    .WIDTH(1)
) cond1006 (
    .clk(cond1006_clk),
    .done(cond1006_done),
    .in(cond1006_in),
    .out(cond1006_out),
    .reset(cond1006_reset),
    .write_en(cond1006_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1006 (
    .in(cond_wire1006_in),
    .out(cond_wire1006_out)
);
std_reg # (
    .WIDTH(1)
) cond1007 (
    .clk(cond1007_clk),
    .done(cond1007_done),
    .in(cond1007_in),
    .out(cond1007_out),
    .reset(cond1007_reset),
    .write_en(cond1007_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1007 (
    .in(cond_wire1007_in),
    .out(cond_wire1007_out)
);
std_reg # (
    .WIDTH(1)
) cond1008 (
    .clk(cond1008_clk),
    .done(cond1008_done),
    .in(cond1008_in),
    .out(cond1008_out),
    .reset(cond1008_reset),
    .write_en(cond1008_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1008 (
    .in(cond_wire1008_in),
    .out(cond_wire1008_out)
);
std_reg # (
    .WIDTH(1)
) cond1009 (
    .clk(cond1009_clk),
    .done(cond1009_done),
    .in(cond1009_in),
    .out(cond1009_out),
    .reset(cond1009_reset),
    .write_en(cond1009_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1009 (
    .in(cond_wire1009_in),
    .out(cond_wire1009_out)
);
std_reg # (
    .WIDTH(1)
) cond1010 (
    .clk(cond1010_clk),
    .done(cond1010_done),
    .in(cond1010_in),
    .out(cond1010_out),
    .reset(cond1010_reset),
    .write_en(cond1010_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1010 (
    .in(cond_wire1010_in),
    .out(cond_wire1010_out)
);
std_reg # (
    .WIDTH(1)
) cond1011 (
    .clk(cond1011_clk),
    .done(cond1011_done),
    .in(cond1011_in),
    .out(cond1011_out),
    .reset(cond1011_reset),
    .write_en(cond1011_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1011 (
    .in(cond_wire1011_in),
    .out(cond_wire1011_out)
);
std_reg # (
    .WIDTH(1)
) cond1012 (
    .clk(cond1012_clk),
    .done(cond1012_done),
    .in(cond1012_in),
    .out(cond1012_out),
    .reset(cond1012_reset),
    .write_en(cond1012_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1012 (
    .in(cond_wire1012_in),
    .out(cond_wire1012_out)
);
std_reg # (
    .WIDTH(1)
) cond1013 (
    .clk(cond1013_clk),
    .done(cond1013_done),
    .in(cond1013_in),
    .out(cond1013_out),
    .reset(cond1013_reset),
    .write_en(cond1013_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1013 (
    .in(cond_wire1013_in),
    .out(cond_wire1013_out)
);
std_reg # (
    .WIDTH(1)
) cond1014 (
    .clk(cond1014_clk),
    .done(cond1014_done),
    .in(cond1014_in),
    .out(cond1014_out),
    .reset(cond1014_reset),
    .write_en(cond1014_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1014 (
    .in(cond_wire1014_in),
    .out(cond_wire1014_out)
);
std_reg # (
    .WIDTH(1)
) cond1015 (
    .clk(cond1015_clk),
    .done(cond1015_done),
    .in(cond1015_in),
    .out(cond1015_out),
    .reset(cond1015_reset),
    .write_en(cond1015_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1015 (
    .in(cond_wire1015_in),
    .out(cond_wire1015_out)
);
std_reg # (
    .WIDTH(1)
) cond1016 (
    .clk(cond1016_clk),
    .done(cond1016_done),
    .in(cond1016_in),
    .out(cond1016_out),
    .reset(cond1016_reset),
    .write_en(cond1016_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1016 (
    .in(cond_wire1016_in),
    .out(cond_wire1016_out)
);
std_reg # (
    .WIDTH(1)
) cond1017 (
    .clk(cond1017_clk),
    .done(cond1017_done),
    .in(cond1017_in),
    .out(cond1017_out),
    .reset(cond1017_reset),
    .write_en(cond1017_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1017 (
    .in(cond_wire1017_in),
    .out(cond_wire1017_out)
);
std_reg # (
    .WIDTH(1)
) cond1018 (
    .clk(cond1018_clk),
    .done(cond1018_done),
    .in(cond1018_in),
    .out(cond1018_out),
    .reset(cond1018_reset),
    .write_en(cond1018_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1018 (
    .in(cond_wire1018_in),
    .out(cond_wire1018_out)
);
std_reg # (
    .WIDTH(1)
) cond1019 (
    .clk(cond1019_clk),
    .done(cond1019_done),
    .in(cond1019_in),
    .out(cond1019_out),
    .reset(cond1019_reset),
    .write_en(cond1019_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1019 (
    .in(cond_wire1019_in),
    .out(cond_wire1019_out)
);
std_reg # (
    .WIDTH(1)
) cond1020 (
    .clk(cond1020_clk),
    .done(cond1020_done),
    .in(cond1020_in),
    .out(cond1020_out),
    .reset(cond1020_reset),
    .write_en(cond1020_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1020 (
    .in(cond_wire1020_in),
    .out(cond_wire1020_out)
);
std_reg # (
    .WIDTH(1)
) cond1021 (
    .clk(cond1021_clk),
    .done(cond1021_done),
    .in(cond1021_in),
    .out(cond1021_out),
    .reset(cond1021_reset),
    .write_en(cond1021_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1021 (
    .in(cond_wire1021_in),
    .out(cond_wire1021_out)
);
std_reg # (
    .WIDTH(1)
) cond1022 (
    .clk(cond1022_clk),
    .done(cond1022_done),
    .in(cond1022_in),
    .out(cond1022_out),
    .reset(cond1022_reset),
    .write_en(cond1022_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1022 (
    .in(cond_wire1022_in),
    .out(cond_wire1022_out)
);
std_reg # (
    .WIDTH(1)
) cond1023 (
    .clk(cond1023_clk),
    .done(cond1023_done),
    .in(cond1023_in),
    .out(cond1023_out),
    .reset(cond1023_reset),
    .write_en(cond1023_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1023 (
    .in(cond_wire1023_in),
    .out(cond_wire1023_out)
);
std_reg # (
    .WIDTH(1)
) cond1024 (
    .clk(cond1024_clk),
    .done(cond1024_done),
    .in(cond1024_in),
    .out(cond1024_out),
    .reset(cond1024_reset),
    .write_en(cond1024_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1024 (
    .in(cond_wire1024_in),
    .out(cond_wire1024_out)
);
std_reg # (
    .WIDTH(1)
) cond1025 (
    .clk(cond1025_clk),
    .done(cond1025_done),
    .in(cond1025_in),
    .out(cond1025_out),
    .reset(cond1025_reset),
    .write_en(cond1025_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1025 (
    .in(cond_wire1025_in),
    .out(cond_wire1025_out)
);
std_reg # (
    .WIDTH(1)
) cond1026 (
    .clk(cond1026_clk),
    .done(cond1026_done),
    .in(cond1026_in),
    .out(cond1026_out),
    .reset(cond1026_reset),
    .write_en(cond1026_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1026 (
    .in(cond_wire1026_in),
    .out(cond_wire1026_out)
);
std_reg # (
    .WIDTH(1)
) cond1027 (
    .clk(cond1027_clk),
    .done(cond1027_done),
    .in(cond1027_in),
    .out(cond1027_out),
    .reset(cond1027_reset),
    .write_en(cond1027_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1027 (
    .in(cond_wire1027_in),
    .out(cond_wire1027_out)
);
std_reg # (
    .WIDTH(1)
) cond1028 (
    .clk(cond1028_clk),
    .done(cond1028_done),
    .in(cond1028_in),
    .out(cond1028_out),
    .reset(cond1028_reset),
    .write_en(cond1028_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1028 (
    .in(cond_wire1028_in),
    .out(cond_wire1028_out)
);
std_reg # (
    .WIDTH(1)
) cond1029 (
    .clk(cond1029_clk),
    .done(cond1029_done),
    .in(cond1029_in),
    .out(cond1029_out),
    .reset(cond1029_reset),
    .write_en(cond1029_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1029 (
    .in(cond_wire1029_in),
    .out(cond_wire1029_out)
);
std_reg # (
    .WIDTH(1)
) cond1030 (
    .clk(cond1030_clk),
    .done(cond1030_done),
    .in(cond1030_in),
    .out(cond1030_out),
    .reset(cond1030_reset),
    .write_en(cond1030_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1030 (
    .in(cond_wire1030_in),
    .out(cond_wire1030_out)
);
std_reg # (
    .WIDTH(1)
) cond1031 (
    .clk(cond1031_clk),
    .done(cond1031_done),
    .in(cond1031_in),
    .out(cond1031_out),
    .reset(cond1031_reset),
    .write_en(cond1031_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1031 (
    .in(cond_wire1031_in),
    .out(cond_wire1031_out)
);
std_reg # (
    .WIDTH(1)
) cond1032 (
    .clk(cond1032_clk),
    .done(cond1032_done),
    .in(cond1032_in),
    .out(cond1032_out),
    .reset(cond1032_reset),
    .write_en(cond1032_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1032 (
    .in(cond_wire1032_in),
    .out(cond_wire1032_out)
);
std_reg # (
    .WIDTH(1)
) cond1033 (
    .clk(cond1033_clk),
    .done(cond1033_done),
    .in(cond1033_in),
    .out(cond1033_out),
    .reset(cond1033_reset),
    .write_en(cond1033_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1033 (
    .in(cond_wire1033_in),
    .out(cond_wire1033_out)
);
std_reg # (
    .WIDTH(1)
) cond1034 (
    .clk(cond1034_clk),
    .done(cond1034_done),
    .in(cond1034_in),
    .out(cond1034_out),
    .reset(cond1034_reset),
    .write_en(cond1034_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1034 (
    .in(cond_wire1034_in),
    .out(cond_wire1034_out)
);
std_reg # (
    .WIDTH(1)
) cond1035 (
    .clk(cond1035_clk),
    .done(cond1035_done),
    .in(cond1035_in),
    .out(cond1035_out),
    .reset(cond1035_reset),
    .write_en(cond1035_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1035 (
    .in(cond_wire1035_in),
    .out(cond_wire1035_out)
);
std_reg # (
    .WIDTH(1)
) cond1036 (
    .clk(cond1036_clk),
    .done(cond1036_done),
    .in(cond1036_in),
    .out(cond1036_out),
    .reset(cond1036_reset),
    .write_en(cond1036_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1036 (
    .in(cond_wire1036_in),
    .out(cond_wire1036_out)
);
std_reg # (
    .WIDTH(1)
) cond1037 (
    .clk(cond1037_clk),
    .done(cond1037_done),
    .in(cond1037_in),
    .out(cond1037_out),
    .reset(cond1037_reset),
    .write_en(cond1037_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1037 (
    .in(cond_wire1037_in),
    .out(cond_wire1037_out)
);
std_reg # (
    .WIDTH(1)
) cond1038 (
    .clk(cond1038_clk),
    .done(cond1038_done),
    .in(cond1038_in),
    .out(cond1038_out),
    .reset(cond1038_reset),
    .write_en(cond1038_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1038 (
    .in(cond_wire1038_in),
    .out(cond_wire1038_out)
);
std_reg # (
    .WIDTH(1)
) cond1039 (
    .clk(cond1039_clk),
    .done(cond1039_done),
    .in(cond1039_in),
    .out(cond1039_out),
    .reset(cond1039_reset),
    .write_en(cond1039_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1039 (
    .in(cond_wire1039_in),
    .out(cond_wire1039_out)
);
std_reg # (
    .WIDTH(1)
) cond1040 (
    .clk(cond1040_clk),
    .done(cond1040_done),
    .in(cond1040_in),
    .out(cond1040_out),
    .reset(cond1040_reset),
    .write_en(cond1040_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1040 (
    .in(cond_wire1040_in),
    .out(cond_wire1040_out)
);
std_reg # (
    .WIDTH(1)
) cond1041 (
    .clk(cond1041_clk),
    .done(cond1041_done),
    .in(cond1041_in),
    .out(cond1041_out),
    .reset(cond1041_reset),
    .write_en(cond1041_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1041 (
    .in(cond_wire1041_in),
    .out(cond_wire1041_out)
);
std_reg # (
    .WIDTH(1)
) cond1042 (
    .clk(cond1042_clk),
    .done(cond1042_done),
    .in(cond1042_in),
    .out(cond1042_out),
    .reset(cond1042_reset),
    .write_en(cond1042_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1042 (
    .in(cond_wire1042_in),
    .out(cond_wire1042_out)
);
std_reg # (
    .WIDTH(1)
) cond1043 (
    .clk(cond1043_clk),
    .done(cond1043_done),
    .in(cond1043_in),
    .out(cond1043_out),
    .reset(cond1043_reset),
    .write_en(cond1043_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1043 (
    .in(cond_wire1043_in),
    .out(cond_wire1043_out)
);
std_reg # (
    .WIDTH(1)
) cond1044 (
    .clk(cond1044_clk),
    .done(cond1044_done),
    .in(cond1044_in),
    .out(cond1044_out),
    .reset(cond1044_reset),
    .write_en(cond1044_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1044 (
    .in(cond_wire1044_in),
    .out(cond_wire1044_out)
);
std_reg # (
    .WIDTH(1)
) cond1045 (
    .clk(cond1045_clk),
    .done(cond1045_done),
    .in(cond1045_in),
    .out(cond1045_out),
    .reset(cond1045_reset),
    .write_en(cond1045_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1045 (
    .in(cond_wire1045_in),
    .out(cond_wire1045_out)
);
std_reg # (
    .WIDTH(1)
) cond1046 (
    .clk(cond1046_clk),
    .done(cond1046_done),
    .in(cond1046_in),
    .out(cond1046_out),
    .reset(cond1046_reset),
    .write_en(cond1046_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1046 (
    .in(cond_wire1046_in),
    .out(cond_wire1046_out)
);
std_reg # (
    .WIDTH(1)
) cond1047 (
    .clk(cond1047_clk),
    .done(cond1047_done),
    .in(cond1047_in),
    .out(cond1047_out),
    .reset(cond1047_reset),
    .write_en(cond1047_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1047 (
    .in(cond_wire1047_in),
    .out(cond_wire1047_out)
);
std_reg # (
    .WIDTH(1)
) cond1048 (
    .clk(cond1048_clk),
    .done(cond1048_done),
    .in(cond1048_in),
    .out(cond1048_out),
    .reset(cond1048_reset),
    .write_en(cond1048_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1048 (
    .in(cond_wire1048_in),
    .out(cond_wire1048_out)
);
std_reg # (
    .WIDTH(1)
) cond1049 (
    .clk(cond1049_clk),
    .done(cond1049_done),
    .in(cond1049_in),
    .out(cond1049_out),
    .reset(cond1049_reset),
    .write_en(cond1049_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1049 (
    .in(cond_wire1049_in),
    .out(cond_wire1049_out)
);
std_reg # (
    .WIDTH(1)
) cond1050 (
    .clk(cond1050_clk),
    .done(cond1050_done),
    .in(cond1050_in),
    .out(cond1050_out),
    .reset(cond1050_reset),
    .write_en(cond1050_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1050 (
    .in(cond_wire1050_in),
    .out(cond_wire1050_out)
);
std_reg # (
    .WIDTH(1)
) cond1051 (
    .clk(cond1051_clk),
    .done(cond1051_done),
    .in(cond1051_in),
    .out(cond1051_out),
    .reset(cond1051_reset),
    .write_en(cond1051_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1051 (
    .in(cond_wire1051_in),
    .out(cond_wire1051_out)
);
std_reg # (
    .WIDTH(1)
) cond1052 (
    .clk(cond1052_clk),
    .done(cond1052_done),
    .in(cond1052_in),
    .out(cond1052_out),
    .reset(cond1052_reset),
    .write_en(cond1052_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1052 (
    .in(cond_wire1052_in),
    .out(cond_wire1052_out)
);
std_reg # (
    .WIDTH(1)
) fsm (
    .clk(fsm_clk),
    .done(fsm_done),
    .in(fsm_in),
    .out(fsm_out),
    .reset(fsm_reset),
    .write_en(fsm_write_en)
);
std_reg # (
    .WIDTH(6)
) fsm0 (
    .clk(fsm0_clk),
    .done(fsm0_done),
    .in(fsm0_in),
    .out(fsm0_out),
    .reset(fsm0_reset),
    .write_en(fsm0_write_en)
);
undef # (
    .WIDTH(1)
) ud (
    .out(ud_out)
);
std_add # (
    .WIDTH(6)
) adder (
    .left(adder_left),
    .out(adder_out),
    .right(adder_right)
);
undef # (
    .WIDTH(1)
) ud0 (
    .out(ud0_out)
);
std_add # (
    .WIDTH(1)
) adder0 (
    .left(adder0_left),
    .out(adder0_out),
    .right(adder0_right)
);
std_reg # (
    .WIDTH(1)
) signal_reg (
    .clk(signal_reg_clk),
    .done(signal_reg_done),
    .in(signal_reg_in),
    .out(signal_reg_out),
    .reset(signal_reg_reset),
    .write_en(signal_reg_write_en)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_seq_go (
    .in(early_reset_static_seq_go_in),
    .out(early_reset_static_seq_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_seq_done (
    .in(early_reset_static_seq_done_in),
    .out(early_reset_static_seq_done_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par0_go (
    .in(early_reset_static_par0_go_in),
    .out(early_reset_static_par0_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par0_done (
    .in(early_reset_static_par0_done_in),
    .out(early_reset_static_par0_done_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_seq_go (
    .in(wrapper_early_reset_static_seq_go_in),
    .out(wrapper_early_reset_static_seq_go_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_seq_done (
    .in(wrapper_early_reset_static_seq_done_in),
    .out(wrapper_early_reset_static_seq_done_out)
);
wire _guard0 = 1;
wire _guard1 = cond_wire98_out;
wire _guard2 = early_reset_static_par0_go_out;
wire _guard3 = _guard1 & _guard2;
wire _guard4 = cond_wire96_out;
wire _guard5 = early_reset_static_par0_go_out;
wire _guard6 = _guard4 & _guard5;
wire _guard7 = fsm_out == 1'd0;
wire _guard8 = cond_wire96_out;
wire _guard9 = _guard7 & _guard8;
wire _guard10 = fsm_out == 1'd0;
wire _guard11 = _guard9 & _guard10;
wire _guard12 = fsm_out == 1'd0;
wire _guard13 = cond_wire98_out;
wire _guard14 = _guard12 & _guard13;
wire _guard15 = fsm_out == 1'd0;
wire _guard16 = _guard14 & _guard15;
wire _guard17 = _guard11 | _guard16;
wire _guard18 = early_reset_static_par0_go_out;
wire _guard19 = _guard17 & _guard18;
wire _guard20 = fsm_out == 1'd0;
wire _guard21 = cond_wire96_out;
wire _guard22 = _guard20 & _guard21;
wire _guard23 = fsm_out == 1'd0;
wire _guard24 = _guard22 & _guard23;
wire _guard25 = fsm_out == 1'd0;
wire _guard26 = cond_wire98_out;
wire _guard27 = _guard25 & _guard26;
wire _guard28 = fsm_out == 1'd0;
wire _guard29 = _guard27 & _guard28;
wire _guard30 = _guard24 | _guard29;
wire _guard31 = early_reset_static_par0_go_out;
wire _guard32 = _guard30 & _guard31;
wire _guard33 = fsm_out == 1'd0;
wire _guard34 = cond_wire96_out;
wire _guard35 = _guard33 & _guard34;
wire _guard36 = fsm_out == 1'd0;
wire _guard37 = _guard35 & _guard36;
wire _guard38 = fsm_out == 1'd0;
wire _guard39 = cond_wire98_out;
wire _guard40 = _guard38 & _guard39;
wire _guard41 = fsm_out == 1'd0;
wire _guard42 = _guard40 & _guard41;
wire _guard43 = _guard37 | _guard42;
wire _guard44 = early_reset_static_par0_go_out;
wire _guard45 = _guard43 & _guard44;
wire _guard46 = cond_wire110_out;
wire _guard47 = early_reset_static_par0_go_out;
wire _guard48 = _guard46 & _guard47;
wire _guard49 = cond_wire108_out;
wire _guard50 = early_reset_static_par0_go_out;
wire _guard51 = _guard49 & _guard50;
wire _guard52 = fsm_out == 1'd0;
wire _guard53 = cond_wire108_out;
wire _guard54 = _guard52 & _guard53;
wire _guard55 = fsm_out == 1'd0;
wire _guard56 = _guard54 & _guard55;
wire _guard57 = fsm_out == 1'd0;
wire _guard58 = cond_wire110_out;
wire _guard59 = _guard57 & _guard58;
wire _guard60 = fsm_out == 1'd0;
wire _guard61 = _guard59 & _guard60;
wire _guard62 = _guard56 | _guard61;
wire _guard63 = early_reset_static_par0_go_out;
wire _guard64 = _guard62 & _guard63;
wire _guard65 = fsm_out == 1'd0;
wire _guard66 = cond_wire108_out;
wire _guard67 = _guard65 & _guard66;
wire _guard68 = fsm_out == 1'd0;
wire _guard69 = _guard67 & _guard68;
wire _guard70 = fsm_out == 1'd0;
wire _guard71 = cond_wire110_out;
wire _guard72 = _guard70 & _guard71;
wire _guard73 = fsm_out == 1'd0;
wire _guard74 = _guard72 & _guard73;
wire _guard75 = _guard69 | _guard74;
wire _guard76 = early_reset_static_par0_go_out;
wire _guard77 = _guard75 & _guard76;
wire _guard78 = fsm_out == 1'd0;
wire _guard79 = cond_wire108_out;
wire _guard80 = _guard78 & _guard79;
wire _guard81 = fsm_out == 1'd0;
wire _guard82 = _guard80 & _guard81;
wire _guard83 = fsm_out == 1'd0;
wire _guard84 = cond_wire110_out;
wire _guard85 = _guard83 & _guard84;
wire _guard86 = fsm_out == 1'd0;
wire _guard87 = _guard85 & _guard86;
wire _guard88 = _guard82 | _guard87;
wire _guard89 = early_reset_static_par0_go_out;
wire _guard90 = _guard88 & _guard89;
wire _guard91 = cond_wire129_out;
wire _guard92 = early_reset_static_par0_go_out;
wire _guard93 = _guard91 & _guard92;
wire _guard94 = cond_wire129_out;
wire _guard95 = early_reset_static_par0_go_out;
wire _guard96 = _guard94 & _guard95;
wire _guard97 = cond_wire97_out;
wire _guard98 = early_reset_static_par0_go_out;
wire _guard99 = _guard97 & _guard98;
wire _guard100 = cond_wire97_out;
wire _guard101 = early_reset_static_par0_go_out;
wire _guard102 = _guard100 & _guard101;
wire _guard103 = cond_wire158_out;
wire _guard104 = early_reset_static_par0_go_out;
wire _guard105 = _guard103 & _guard104;
wire _guard106 = cond_wire158_out;
wire _guard107 = early_reset_static_par0_go_out;
wire _guard108 = _guard106 & _guard107;
wire _guard109 = cond_wire195_out;
wire _guard110 = early_reset_static_par0_go_out;
wire _guard111 = _guard109 & _guard110;
wire _guard112 = cond_wire193_out;
wire _guard113 = early_reset_static_par0_go_out;
wire _guard114 = _guard112 & _guard113;
wire _guard115 = fsm_out == 1'd0;
wire _guard116 = cond_wire193_out;
wire _guard117 = _guard115 & _guard116;
wire _guard118 = fsm_out == 1'd0;
wire _guard119 = _guard117 & _guard118;
wire _guard120 = fsm_out == 1'd0;
wire _guard121 = cond_wire195_out;
wire _guard122 = _guard120 & _guard121;
wire _guard123 = fsm_out == 1'd0;
wire _guard124 = _guard122 & _guard123;
wire _guard125 = _guard119 | _guard124;
wire _guard126 = early_reset_static_par0_go_out;
wire _guard127 = _guard125 & _guard126;
wire _guard128 = fsm_out == 1'd0;
wire _guard129 = cond_wire193_out;
wire _guard130 = _guard128 & _guard129;
wire _guard131 = fsm_out == 1'd0;
wire _guard132 = _guard130 & _guard131;
wire _guard133 = fsm_out == 1'd0;
wire _guard134 = cond_wire195_out;
wire _guard135 = _guard133 & _guard134;
wire _guard136 = fsm_out == 1'd0;
wire _guard137 = _guard135 & _guard136;
wire _guard138 = _guard132 | _guard137;
wire _guard139 = early_reset_static_par0_go_out;
wire _guard140 = _guard138 & _guard139;
wire _guard141 = fsm_out == 1'd0;
wire _guard142 = cond_wire193_out;
wire _guard143 = _guard141 & _guard142;
wire _guard144 = fsm_out == 1'd0;
wire _guard145 = _guard143 & _guard144;
wire _guard146 = fsm_out == 1'd0;
wire _guard147 = cond_wire195_out;
wire _guard148 = _guard146 & _guard147;
wire _guard149 = fsm_out == 1'd0;
wire _guard150 = _guard148 & _guard149;
wire _guard151 = _guard145 | _guard150;
wire _guard152 = early_reset_static_par0_go_out;
wire _guard153 = _guard151 & _guard152;
wire _guard154 = cond_wire166_out;
wire _guard155 = early_reset_static_par0_go_out;
wire _guard156 = _guard154 & _guard155;
wire _guard157 = cond_wire166_out;
wire _guard158 = early_reset_static_par0_go_out;
wire _guard159 = _guard157 & _guard158;
wire _guard160 = cond_wire170_out;
wire _guard161 = early_reset_static_par0_go_out;
wire _guard162 = _guard160 & _guard161;
wire _guard163 = cond_wire170_out;
wire _guard164 = early_reset_static_par0_go_out;
wire _guard165 = _guard163 & _guard164;
wire _guard166 = cond_wire244_out;
wire _guard167 = early_reset_static_par0_go_out;
wire _guard168 = _guard166 & _guard167;
wire _guard169 = cond_wire242_out;
wire _guard170 = early_reset_static_par0_go_out;
wire _guard171 = _guard169 & _guard170;
wire _guard172 = fsm_out == 1'd0;
wire _guard173 = cond_wire242_out;
wire _guard174 = _guard172 & _guard173;
wire _guard175 = fsm_out == 1'd0;
wire _guard176 = _guard174 & _guard175;
wire _guard177 = fsm_out == 1'd0;
wire _guard178 = cond_wire244_out;
wire _guard179 = _guard177 & _guard178;
wire _guard180 = fsm_out == 1'd0;
wire _guard181 = _guard179 & _guard180;
wire _guard182 = _guard176 | _guard181;
wire _guard183 = early_reset_static_par0_go_out;
wire _guard184 = _guard182 & _guard183;
wire _guard185 = fsm_out == 1'd0;
wire _guard186 = cond_wire242_out;
wire _guard187 = _guard185 & _guard186;
wire _guard188 = fsm_out == 1'd0;
wire _guard189 = _guard187 & _guard188;
wire _guard190 = fsm_out == 1'd0;
wire _guard191 = cond_wire244_out;
wire _guard192 = _guard190 & _guard191;
wire _guard193 = fsm_out == 1'd0;
wire _guard194 = _guard192 & _guard193;
wire _guard195 = _guard189 | _guard194;
wire _guard196 = early_reset_static_par0_go_out;
wire _guard197 = _guard195 & _guard196;
wire _guard198 = fsm_out == 1'd0;
wire _guard199 = cond_wire242_out;
wire _guard200 = _guard198 & _guard199;
wire _guard201 = fsm_out == 1'd0;
wire _guard202 = _guard200 & _guard201;
wire _guard203 = fsm_out == 1'd0;
wire _guard204 = cond_wire244_out;
wire _guard205 = _guard203 & _guard204;
wire _guard206 = fsm_out == 1'd0;
wire _guard207 = _guard205 & _guard206;
wire _guard208 = _guard202 | _guard207;
wire _guard209 = early_reset_static_par0_go_out;
wire _guard210 = _guard208 & _guard209;
wire _guard211 = cond_wire274_out;
wire _guard212 = early_reset_static_par0_go_out;
wire _guard213 = _guard211 & _guard212;
wire _guard214 = cond_wire274_out;
wire _guard215 = early_reset_static_par0_go_out;
wire _guard216 = _guard214 & _guard215;
wire _guard217 = cond_wire227_out;
wire _guard218 = early_reset_static_par0_go_out;
wire _guard219 = _guard217 & _guard218;
wire _guard220 = cond_wire227_out;
wire _guard221 = early_reset_static_par0_go_out;
wire _guard222 = _guard220 & _guard221;
wire _guard223 = cond_wire313_out;
wire _guard224 = early_reset_static_par0_go_out;
wire _guard225 = _guard223 & _guard224;
wire _guard226 = cond_wire311_out;
wire _guard227 = early_reset_static_par0_go_out;
wire _guard228 = _guard226 & _guard227;
wire _guard229 = fsm_out == 1'd0;
wire _guard230 = cond_wire311_out;
wire _guard231 = _guard229 & _guard230;
wire _guard232 = fsm_out == 1'd0;
wire _guard233 = _guard231 & _guard232;
wire _guard234 = fsm_out == 1'd0;
wire _guard235 = cond_wire313_out;
wire _guard236 = _guard234 & _guard235;
wire _guard237 = fsm_out == 1'd0;
wire _guard238 = _guard236 & _guard237;
wire _guard239 = _guard233 | _guard238;
wire _guard240 = early_reset_static_par0_go_out;
wire _guard241 = _guard239 & _guard240;
wire _guard242 = fsm_out == 1'd0;
wire _guard243 = cond_wire311_out;
wire _guard244 = _guard242 & _guard243;
wire _guard245 = fsm_out == 1'd0;
wire _guard246 = _guard244 & _guard245;
wire _guard247 = fsm_out == 1'd0;
wire _guard248 = cond_wire313_out;
wire _guard249 = _guard247 & _guard248;
wire _guard250 = fsm_out == 1'd0;
wire _guard251 = _guard249 & _guard250;
wire _guard252 = _guard246 | _guard251;
wire _guard253 = early_reset_static_par0_go_out;
wire _guard254 = _guard252 & _guard253;
wire _guard255 = fsm_out == 1'd0;
wire _guard256 = cond_wire311_out;
wire _guard257 = _guard255 & _guard256;
wire _guard258 = fsm_out == 1'd0;
wire _guard259 = _guard257 & _guard258;
wire _guard260 = fsm_out == 1'd0;
wire _guard261 = cond_wire313_out;
wire _guard262 = _guard260 & _guard261;
wire _guard263 = fsm_out == 1'd0;
wire _guard264 = _guard262 & _guard263;
wire _guard265 = _guard259 | _guard264;
wire _guard266 = early_reset_static_par0_go_out;
wire _guard267 = _guard265 & _guard266;
wire _guard268 = cond_wire350_out;
wire _guard269 = early_reset_static_par0_go_out;
wire _guard270 = _guard268 & _guard269;
wire _guard271 = cond_wire348_out;
wire _guard272 = early_reset_static_par0_go_out;
wire _guard273 = _guard271 & _guard272;
wire _guard274 = fsm_out == 1'd0;
wire _guard275 = cond_wire348_out;
wire _guard276 = _guard274 & _guard275;
wire _guard277 = fsm_out == 1'd0;
wire _guard278 = _guard276 & _guard277;
wire _guard279 = fsm_out == 1'd0;
wire _guard280 = cond_wire350_out;
wire _guard281 = _guard279 & _guard280;
wire _guard282 = fsm_out == 1'd0;
wire _guard283 = _guard281 & _guard282;
wire _guard284 = _guard278 | _guard283;
wire _guard285 = early_reset_static_par0_go_out;
wire _guard286 = _guard284 & _guard285;
wire _guard287 = fsm_out == 1'd0;
wire _guard288 = cond_wire348_out;
wire _guard289 = _guard287 & _guard288;
wire _guard290 = fsm_out == 1'd0;
wire _guard291 = _guard289 & _guard290;
wire _guard292 = fsm_out == 1'd0;
wire _guard293 = cond_wire350_out;
wire _guard294 = _guard292 & _guard293;
wire _guard295 = fsm_out == 1'd0;
wire _guard296 = _guard294 & _guard295;
wire _guard297 = _guard291 | _guard296;
wire _guard298 = early_reset_static_par0_go_out;
wire _guard299 = _guard297 & _guard298;
wire _guard300 = fsm_out == 1'd0;
wire _guard301 = cond_wire348_out;
wire _guard302 = _guard300 & _guard301;
wire _guard303 = fsm_out == 1'd0;
wire _guard304 = _guard302 & _guard303;
wire _guard305 = fsm_out == 1'd0;
wire _guard306 = cond_wire350_out;
wire _guard307 = _guard305 & _guard306;
wire _guard308 = fsm_out == 1'd0;
wire _guard309 = _guard307 & _guard308;
wire _guard310 = _guard304 | _guard309;
wire _guard311 = early_reset_static_par0_go_out;
wire _guard312 = _guard310 & _guard311;
wire _guard313 = cond_wire308_out;
wire _guard314 = early_reset_static_par0_go_out;
wire _guard315 = _guard313 & _guard314;
wire _guard316 = cond_wire308_out;
wire _guard317 = early_reset_static_par0_go_out;
wire _guard318 = _guard316 & _guard317;
wire _guard319 = cond_wire345_out;
wire _guard320 = early_reset_static_par0_go_out;
wire _guard321 = _guard319 & _guard320;
wire _guard322 = cond_wire345_out;
wire _guard323 = early_reset_static_par0_go_out;
wire _guard324 = _guard322 & _guard323;
wire _guard325 = cond_wire410_out;
wire _guard326 = early_reset_static_par0_go_out;
wire _guard327 = _guard325 & _guard326;
wire _guard328 = cond_wire410_out;
wire _guard329 = early_reset_static_par0_go_out;
wire _guard330 = _guard328 & _guard329;
wire _guard331 = cond_wire353_out;
wire _guard332 = early_reset_static_par0_go_out;
wire _guard333 = _guard331 & _guard332;
wire _guard334 = cond_wire353_out;
wire _guard335 = early_reset_static_par0_go_out;
wire _guard336 = _guard334 & _guard335;
wire _guard337 = cond_wire418_out;
wire _guard338 = early_reset_static_par0_go_out;
wire _guard339 = _guard337 & _guard338;
wire _guard340 = cond_wire418_out;
wire _guard341 = early_reset_static_par0_go_out;
wire _guard342 = _guard340 & _guard341;
wire _guard343 = cond_wire393_out;
wire _guard344 = early_reset_static_par0_go_out;
wire _guard345 = _guard343 & _guard344;
wire _guard346 = cond_wire393_out;
wire _guard347 = early_reset_static_par0_go_out;
wire _guard348 = _guard346 & _guard347;
wire _guard349 = cond_wire406_out;
wire _guard350 = early_reset_static_par0_go_out;
wire _guard351 = _guard349 & _guard350;
wire _guard352 = cond_wire406_out;
wire _guard353 = early_reset_static_par0_go_out;
wire _guard354 = _guard352 & _guard353;
wire _guard355 = cond_wire508_out;
wire _guard356 = early_reset_static_par0_go_out;
wire _guard357 = _guard355 & _guard356;
wire _guard358 = cond_wire506_out;
wire _guard359 = early_reset_static_par0_go_out;
wire _guard360 = _guard358 & _guard359;
wire _guard361 = fsm_out == 1'd0;
wire _guard362 = cond_wire506_out;
wire _guard363 = _guard361 & _guard362;
wire _guard364 = fsm_out == 1'd0;
wire _guard365 = _guard363 & _guard364;
wire _guard366 = fsm_out == 1'd0;
wire _guard367 = cond_wire508_out;
wire _guard368 = _guard366 & _guard367;
wire _guard369 = fsm_out == 1'd0;
wire _guard370 = _guard368 & _guard369;
wire _guard371 = _guard365 | _guard370;
wire _guard372 = early_reset_static_par0_go_out;
wire _guard373 = _guard371 & _guard372;
wire _guard374 = fsm_out == 1'd0;
wire _guard375 = cond_wire506_out;
wire _guard376 = _guard374 & _guard375;
wire _guard377 = fsm_out == 1'd0;
wire _guard378 = _guard376 & _guard377;
wire _guard379 = fsm_out == 1'd0;
wire _guard380 = cond_wire508_out;
wire _guard381 = _guard379 & _guard380;
wire _guard382 = fsm_out == 1'd0;
wire _guard383 = _guard381 & _guard382;
wire _guard384 = _guard378 | _guard383;
wire _guard385 = early_reset_static_par0_go_out;
wire _guard386 = _guard384 & _guard385;
wire _guard387 = fsm_out == 1'd0;
wire _guard388 = cond_wire506_out;
wire _guard389 = _guard387 & _guard388;
wire _guard390 = fsm_out == 1'd0;
wire _guard391 = _guard389 & _guard390;
wire _guard392 = fsm_out == 1'd0;
wire _guard393 = cond_wire508_out;
wire _guard394 = _guard392 & _guard393;
wire _guard395 = fsm_out == 1'd0;
wire _guard396 = _guard394 & _guard395;
wire _guard397 = _guard391 | _guard396;
wire _guard398 = early_reset_static_par0_go_out;
wire _guard399 = _guard397 & _guard398;
wire _guard400 = cond_wire523_out;
wire _guard401 = early_reset_static_par0_go_out;
wire _guard402 = _guard400 & _guard401;
wire _guard403 = cond_wire523_out;
wire _guard404 = early_reset_static_par0_go_out;
wire _guard405 = _guard403 & _guard404;
wire _guard406 = cond_wire487_out;
wire _guard407 = early_reset_static_par0_go_out;
wire _guard408 = _guard406 & _guard407;
wire _guard409 = cond_wire487_out;
wire _guard410 = early_reset_static_par0_go_out;
wire _guard411 = _guard409 & _guard410;
wire _guard412 = cond_wire576_out;
wire _guard413 = early_reset_static_par0_go_out;
wire _guard414 = _guard412 & _guard413;
wire _guard415 = cond_wire576_out;
wire _guard416 = early_reset_static_par0_go_out;
wire _guard417 = _guard415 & _guard416;
wire _guard418 = cond_wire617_out;
wire _guard419 = early_reset_static_par0_go_out;
wire _guard420 = _guard418 & _guard419;
wire _guard421 = cond_wire617_out;
wire _guard422 = early_reset_static_par0_go_out;
wire _guard423 = _guard421 & _guard422;
wire _guard424 = cond_wire662_out;
wire _guard425 = early_reset_static_par0_go_out;
wire _guard426 = _guard424 & _guard425;
wire _guard427 = cond_wire660_out;
wire _guard428 = early_reset_static_par0_go_out;
wire _guard429 = _guard427 & _guard428;
wire _guard430 = fsm_out == 1'd0;
wire _guard431 = cond_wire660_out;
wire _guard432 = _guard430 & _guard431;
wire _guard433 = fsm_out == 1'd0;
wire _guard434 = _guard432 & _guard433;
wire _guard435 = fsm_out == 1'd0;
wire _guard436 = cond_wire662_out;
wire _guard437 = _guard435 & _guard436;
wire _guard438 = fsm_out == 1'd0;
wire _guard439 = _guard437 & _guard438;
wire _guard440 = _guard434 | _guard439;
wire _guard441 = early_reset_static_par0_go_out;
wire _guard442 = _guard440 & _guard441;
wire _guard443 = fsm_out == 1'd0;
wire _guard444 = cond_wire660_out;
wire _guard445 = _guard443 & _guard444;
wire _guard446 = fsm_out == 1'd0;
wire _guard447 = _guard445 & _guard446;
wire _guard448 = fsm_out == 1'd0;
wire _guard449 = cond_wire662_out;
wire _guard450 = _guard448 & _guard449;
wire _guard451 = fsm_out == 1'd0;
wire _guard452 = _guard450 & _guard451;
wire _guard453 = _guard447 | _guard452;
wire _guard454 = early_reset_static_par0_go_out;
wire _guard455 = _guard453 & _guard454;
wire _guard456 = fsm_out == 1'd0;
wire _guard457 = cond_wire660_out;
wire _guard458 = _guard456 & _guard457;
wire _guard459 = fsm_out == 1'd0;
wire _guard460 = _guard458 & _guard459;
wire _guard461 = fsm_out == 1'd0;
wire _guard462 = cond_wire662_out;
wire _guard463 = _guard461 & _guard462;
wire _guard464 = fsm_out == 1'd0;
wire _guard465 = _guard463 & _guard464;
wire _guard466 = _guard460 | _guard465;
wire _guard467 = early_reset_static_par0_go_out;
wire _guard468 = _guard466 & _guard467;
wire _guard469 = cond_wire687_out;
wire _guard470 = early_reset_static_par0_go_out;
wire _guard471 = _guard469 & _guard470;
wire _guard472 = cond_wire685_out;
wire _guard473 = early_reset_static_par0_go_out;
wire _guard474 = _guard472 & _guard473;
wire _guard475 = fsm_out == 1'd0;
wire _guard476 = cond_wire685_out;
wire _guard477 = _guard475 & _guard476;
wire _guard478 = fsm_out == 1'd0;
wire _guard479 = _guard477 & _guard478;
wire _guard480 = fsm_out == 1'd0;
wire _guard481 = cond_wire687_out;
wire _guard482 = _guard480 & _guard481;
wire _guard483 = fsm_out == 1'd0;
wire _guard484 = _guard482 & _guard483;
wire _guard485 = _guard479 | _guard484;
wire _guard486 = early_reset_static_par0_go_out;
wire _guard487 = _guard485 & _guard486;
wire _guard488 = fsm_out == 1'd0;
wire _guard489 = cond_wire685_out;
wire _guard490 = _guard488 & _guard489;
wire _guard491 = fsm_out == 1'd0;
wire _guard492 = _guard490 & _guard491;
wire _guard493 = fsm_out == 1'd0;
wire _guard494 = cond_wire687_out;
wire _guard495 = _guard493 & _guard494;
wire _guard496 = fsm_out == 1'd0;
wire _guard497 = _guard495 & _guard496;
wire _guard498 = _guard492 | _guard497;
wire _guard499 = early_reset_static_par0_go_out;
wire _guard500 = _guard498 & _guard499;
wire _guard501 = fsm_out == 1'd0;
wire _guard502 = cond_wire685_out;
wire _guard503 = _guard501 & _guard502;
wire _guard504 = fsm_out == 1'd0;
wire _guard505 = _guard503 & _guard504;
wire _guard506 = fsm_out == 1'd0;
wire _guard507 = cond_wire687_out;
wire _guard508 = _guard506 & _guard507;
wire _guard509 = fsm_out == 1'd0;
wire _guard510 = _guard508 & _guard509;
wire _guard511 = _guard505 | _guard510;
wire _guard512 = early_reset_static_par0_go_out;
wire _guard513 = _guard511 & _guard512;
wire _guard514 = cond_wire633_out;
wire _guard515 = early_reset_static_par0_go_out;
wire _guard516 = _guard514 & _guard515;
wire _guard517 = cond_wire633_out;
wire _guard518 = early_reset_static_par0_go_out;
wire _guard519 = _guard517 & _guard518;
wire _guard520 = cond_wire653_out;
wire _guard521 = early_reset_static_par0_go_out;
wire _guard522 = _guard520 & _guard521;
wire _guard523 = cond_wire653_out;
wire _guard524 = early_reset_static_par0_go_out;
wire _guard525 = _guard523 & _guard524;
wire _guard526 = cond_wire726_out;
wire _guard527 = early_reset_static_par0_go_out;
wire _guard528 = _guard526 & _guard527;
wire _guard529 = cond_wire726_out;
wire _guard530 = early_reset_static_par0_go_out;
wire _guard531 = _guard529 & _guard530;
wire _guard532 = cond_wire743_out;
wire _guard533 = early_reset_static_par0_go_out;
wire _guard534 = _guard532 & _guard533;
wire _guard535 = cond_wire743_out;
wire _guard536 = early_reset_static_par0_go_out;
wire _guard537 = _guard535 & _guard536;
wire _guard538 = cond_wire808_out;
wire _guard539 = early_reset_static_par0_go_out;
wire _guard540 = _guard538 & _guard539;
wire _guard541 = cond_wire808_out;
wire _guard542 = early_reset_static_par0_go_out;
wire _guard543 = _guard541 & _guard542;
wire _guard544 = cond_wire837_out;
wire _guard545 = early_reset_static_par0_go_out;
wire _guard546 = _guard544 & _guard545;
wire _guard547 = cond_wire835_out;
wire _guard548 = early_reset_static_par0_go_out;
wire _guard549 = _guard547 & _guard548;
wire _guard550 = fsm_out == 1'd0;
wire _guard551 = cond_wire835_out;
wire _guard552 = _guard550 & _guard551;
wire _guard553 = fsm_out == 1'd0;
wire _guard554 = _guard552 & _guard553;
wire _guard555 = fsm_out == 1'd0;
wire _guard556 = cond_wire837_out;
wire _guard557 = _guard555 & _guard556;
wire _guard558 = fsm_out == 1'd0;
wire _guard559 = _guard557 & _guard558;
wire _guard560 = _guard554 | _guard559;
wire _guard561 = early_reset_static_par0_go_out;
wire _guard562 = _guard560 & _guard561;
wire _guard563 = fsm_out == 1'd0;
wire _guard564 = cond_wire835_out;
wire _guard565 = _guard563 & _guard564;
wire _guard566 = fsm_out == 1'd0;
wire _guard567 = _guard565 & _guard566;
wire _guard568 = fsm_out == 1'd0;
wire _guard569 = cond_wire837_out;
wire _guard570 = _guard568 & _guard569;
wire _guard571 = fsm_out == 1'd0;
wire _guard572 = _guard570 & _guard571;
wire _guard573 = _guard567 | _guard572;
wire _guard574 = early_reset_static_par0_go_out;
wire _guard575 = _guard573 & _guard574;
wire _guard576 = fsm_out == 1'd0;
wire _guard577 = cond_wire835_out;
wire _guard578 = _guard576 & _guard577;
wire _guard579 = fsm_out == 1'd0;
wire _guard580 = _guard578 & _guard579;
wire _guard581 = fsm_out == 1'd0;
wire _guard582 = cond_wire837_out;
wire _guard583 = _guard581 & _guard582;
wire _guard584 = fsm_out == 1'd0;
wire _guard585 = _guard583 & _guard584;
wire _guard586 = _guard580 | _guard585;
wire _guard587 = early_reset_static_par0_go_out;
wire _guard588 = _guard586 & _guard587;
wire _guard589 = cond_wire865_out;
wire _guard590 = early_reset_static_par0_go_out;
wire _guard591 = _guard589 & _guard590;
wire _guard592 = cond_wire865_out;
wire _guard593 = early_reset_static_par0_go_out;
wire _guard594 = _guard592 & _guard593;
wire _guard595 = cond_wire824_out;
wire _guard596 = early_reset_static_par0_go_out;
wire _guard597 = _guard595 & _guard596;
wire _guard598 = cond_wire824_out;
wire _guard599 = early_reset_static_par0_go_out;
wire _guard600 = _guard598 & _guard599;
wire _guard601 = cond_wire844_out;
wire _guard602 = early_reset_static_par0_go_out;
wire _guard603 = _guard601 & _guard602;
wire _guard604 = cond_wire844_out;
wire _guard605 = early_reset_static_par0_go_out;
wire _guard606 = _guard604 & _guard605;
wire _guard607 = cond_wire918_out;
wire _guard608 = early_reset_static_par0_go_out;
wire _guard609 = _guard607 & _guard608;
wire _guard610 = cond_wire916_out;
wire _guard611 = early_reset_static_par0_go_out;
wire _guard612 = _guard610 & _guard611;
wire _guard613 = fsm_out == 1'd0;
wire _guard614 = cond_wire916_out;
wire _guard615 = _guard613 & _guard614;
wire _guard616 = fsm_out == 1'd0;
wire _guard617 = _guard615 & _guard616;
wire _guard618 = fsm_out == 1'd0;
wire _guard619 = cond_wire918_out;
wire _guard620 = _guard618 & _guard619;
wire _guard621 = fsm_out == 1'd0;
wire _guard622 = _guard620 & _guard621;
wire _guard623 = _guard617 | _guard622;
wire _guard624 = early_reset_static_par0_go_out;
wire _guard625 = _guard623 & _guard624;
wire _guard626 = fsm_out == 1'd0;
wire _guard627 = cond_wire916_out;
wire _guard628 = _guard626 & _guard627;
wire _guard629 = fsm_out == 1'd0;
wire _guard630 = _guard628 & _guard629;
wire _guard631 = fsm_out == 1'd0;
wire _guard632 = cond_wire918_out;
wire _guard633 = _guard631 & _guard632;
wire _guard634 = fsm_out == 1'd0;
wire _guard635 = _guard633 & _guard634;
wire _guard636 = _guard630 | _guard635;
wire _guard637 = early_reset_static_par0_go_out;
wire _guard638 = _guard636 & _guard637;
wire _guard639 = fsm_out == 1'd0;
wire _guard640 = cond_wire916_out;
wire _guard641 = _guard639 & _guard640;
wire _guard642 = fsm_out == 1'd0;
wire _guard643 = _guard641 & _guard642;
wire _guard644 = fsm_out == 1'd0;
wire _guard645 = cond_wire918_out;
wire _guard646 = _guard644 & _guard645;
wire _guard647 = fsm_out == 1'd0;
wire _guard648 = _guard646 & _guard647;
wire _guard649 = _guard643 | _guard648;
wire _guard650 = early_reset_static_par0_go_out;
wire _guard651 = _guard649 & _guard650;
wire _guard652 = cond_wire861_out;
wire _guard653 = early_reset_static_par0_go_out;
wire _guard654 = _guard652 & _guard653;
wire _guard655 = cond_wire861_out;
wire _guard656 = early_reset_static_par0_go_out;
wire _guard657 = _guard655 & _guard656;
wire _guard658 = cond_wire921_out;
wire _guard659 = early_reset_static_par0_go_out;
wire _guard660 = _guard658 & _guard659;
wire _guard661 = cond_wire921_out;
wire _guard662 = early_reset_static_par0_go_out;
wire _guard663 = _guard661 & _guard662;
wire _guard664 = cond_wire926_out;
wire _guard665 = early_reset_static_par0_go_out;
wire _guard666 = _guard664 & _guard665;
wire _guard667 = cond_wire926_out;
wire _guard668 = early_reset_static_par0_go_out;
wire _guard669 = _guard667 & _guard668;
wire _guard670 = cond_wire954_out;
wire _guard671 = early_reset_static_par0_go_out;
wire _guard672 = _guard670 & _guard671;
wire _guard673 = cond_wire954_out;
wire _guard674 = early_reset_static_par0_go_out;
wire _guard675 = _guard673 & _guard674;
wire _guard676 = cond_wire14_out;
wire _guard677 = early_reset_static_par0_go_out;
wire _guard678 = _guard676 & _guard677;
wire _guard679 = cond_wire14_out;
wire _guard680 = early_reset_static_par0_go_out;
wire _guard681 = _guard679 & _guard680;
wire _guard682 = fsm0_out == 6'd0;
wire _guard683 = early_reset_static_seq_go_out;
wire _guard684 = _guard682 & _guard683;
wire _guard685 = cond_wire74_out;
wire _guard686 = early_reset_static_par0_go_out;
wire _guard687 = _guard685 & _guard686;
wire _guard688 = _guard684 | _guard687;
wire _guard689 = fsm0_out == 6'd0;
wire _guard690 = early_reset_static_seq_go_out;
wire _guard691 = _guard689 & _guard690;
wire _guard692 = cond_wire74_out;
wire _guard693 = early_reset_static_par0_go_out;
wire _guard694 = _guard692 & _guard693;
wire _guard695 = cond_wire79_out;
wire _guard696 = early_reset_static_par0_go_out;
wire _guard697 = _guard695 & _guard696;
wire _guard698 = cond_wire79_out;
wire _guard699 = early_reset_static_par0_go_out;
wire _guard700 = _guard698 & _guard699;
wire _guard701 = fsm0_out == 6'd0;
wire _guard702 = early_reset_static_seq_go_out;
wire _guard703 = _guard701 & _guard702;
wire _guard704 = cond_wire794_out;
wire _guard705 = early_reset_static_par0_go_out;
wire _guard706 = _guard704 & _guard705;
wire _guard707 = _guard703 | _guard706;
wire _guard708 = fsm0_out == 6'd0;
wire _guard709 = early_reset_static_seq_go_out;
wire _guard710 = _guard708 & _guard709;
wire _guard711 = cond_wire794_out;
wire _guard712 = early_reset_static_par0_go_out;
wire _guard713 = _guard711 & _guard712;
wire _guard714 = fsm0_out == 6'd0;
wire _guard715 = early_reset_static_seq_go_out;
wire _guard716 = _guard714 & _guard715;
wire _guard717 = cond_wire859_out;
wire _guard718 = early_reset_static_par0_go_out;
wire _guard719 = _guard717 & _guard718;
wire _guard720 = _guard716 | _guard719;
wire _guard721 = fsm0_out == 6'd0;
wire _guard722 = early_reset_static_seq_go_out;
wire _guard723 = _guard721 & _guard722;
wire _guard724 = cond_wire859_out;
wire _guard725 = early_reset_static_par0_go_out;
wire _guard726 = _guard724 & _guard725;
wire _guard727 = early_reset_static_par0_go_out;
wire _guard728 = early_reset_static_par0_go_out;
wire _guard729 = early_reset_static_par0_go_out;
wire _guard730 = early_reset_static_par0_go_out;
wire _guard731 = early_reset_static_par0_go_out;
wire _guard732 = early_reset_static_par0_go_out;
wire _guard733 = early_reset_static_par0_go_out;
wire _guard734 = early_reset_static_par0_go_out;
wire _guard735 = fsm0_out == 6'd0;
wire _guard736 = early_reset_static_seq_go_out;
wire _guard737 = _guard735 & _guard736;
wire _guard738 = early_reset_static_par0_go_out;
wire _guard739 = _guard737 | _guard738;
wire _guard740 = early_reset_static_par0_go_out;
wire _guard741 = fsm0_out == 6'd0;
wire _guard742 = early_reset_static_seq_go_out;
wire _guard743 = _guard741 & _guard742;
wire _guard744 = fsm0_out == 6'd0;
wire _guard745 = early_reset_static_seq_go_out;
wire _guard746 = _guard744 & _guard745;
wire _guard747 = early_reset_static_par0_go_out;
wire _guard748 = _guard746 | _guard747;
wire _guard749 = fsm0_out == 6'd0;
wire _guard750 = early_reset_static_seq_go_out;
wire _guard751 = _guard749 & _guard750;
wire _guard752 = early_reset_static_par0_go_out;
wire _guard753 = early_reset_static_par0_go_out;
wire _guard754 = early_reset_static_par0_go_out;
wire _guard755 = early_reset_static_par0_go_out;
wire _guard756 = early_reset_static_par0_go_out;
wire _guard757 = fsm0_out == 6'd0;
wire _guard758 = early_reset_static_seq_go_out;
wire _guard759 = _guard757 & _guard758;
wire _guard760 = early_reset_static_par0_go_out;
wire _guard761 = _guard759 | _guard760;
wire _guard762 = early_reset_static_par0_go_out;
wire _guard763 = fsm0_out == 6'd0;
wire _guard764 = early_reset_static_seq_go_out;
wire _guard765 = _guard763 & _guard764;
wire _guard766 = early_reset_static_par0_go_out;
wire _guard767 = early_reset_static_par0_go_out;
wire _guard768 = early_reset_static_par0_go_out;
wire _guard769 = early_reset_static_par0_go_out;
wire _guard770 = early_reset_static_par0_go_out;
wire _guard771 = early_reset_static_par0_go_out;
wire _guard772 = early_reset_static_par0_go_out;
wire _guard773 = early_reset_static_par0_go_out;
wire _guard774 = early_reset_static_par0_go_out;
wire _guard775 = early_reset_static_par0_go_out;
wire _guard776 = fsm0_out == 6'd0;
wire _guard777 = early_reset_static_seq_go_out;
wire _guard778 = _guard776 & _guard777;
wire _guard779 = early_reset_static_par0_go_out;
wire _guard780 = _guard778 | _guard779;
wire _guard781 = early_reset_static_par0_go_out;
wire _guard782 = fsm0_out == 6'd0;
wire _guard783 = early_reset_static_seq_go_out;
wire _guard784 = _guard782 & _guard783;
wire _guard785 = fsm0_out == 6'd0;
wire _guard786 = early_reset_static_seq_go_out;
wire _guard787 = _guard785 & _guard786;
wire _guard788 = early_reset_static_par0_go_out;
wire _guard789 = _guard787 | _guard788;
wire _guard790 = early_reset_static_par0_go_out;
wire _guard791 = fsm0_out == 6'd0;
wire _guard792 = early_reset_static_seq_go_out;
wire _guard793 = _guard791 & _guard792;
wire _guard794 = early_reset_static_par0_go_out;
wire _guard795 = early_reset_static_par0_go_out;
wire _guard796 = fsm0_out == 6'd0;
wire _guard797 = early_reset_static_seq_go_out;
wire _guard798 = _guard796 & _guard797;
wire _guard799 = early_reset_static_par0_go_out;
wire _guard800 = _guard798 | _guard799;
wire _guard801 = early_reset_static_par0_go_out;
wire _guard802 = fsm0_out == 6'd0;
wire _guard803 = early_reset_static_seq_go_out;
wire _guard804 = _guard802 & _guard803;
wire _guard805 = fsm0_out == 6'd0;
wire _guard806 = early_reset_static_seq_go_out;
wire _guard807 = _guard805 & _guard806;
wire _guard808 = early_reset_static_par0_go_out;
wire _guard809 = _guard807 | _guard808;
wire _guard810 = early_reset_static_par0_go_out;
wire _guard811 = fsm0_out == 6'd0;
wire _guard812 = early_reset_static_seq_go_out;
wire _guard813 = _guard811 & _guard812;
wire _guard814 = fsm0_out == 6'd0;
wire _guard815 = early_reset_static_seq_go_out;
wire _guard816 = _guard814 & _guard815;
wire _guard817 = early_reset_static_par0_go_out;
wire _guard818 = _guard816 | _guard817;
wire _guard819 = early_reset_static_par0_go_out;
wire _guard820 = fsm0_out == 6'd0;
wire _guard821 = early_reset_static_seq_go_out;
wire _guard822 = _guard820 & _guard821;
wire _guard823 = early_reset_static_par0_go_out;
wire _guard824 = ~_guard0;
wire _guard825 = early_reset_static_par0_go_out;
wire _guard826 = _guard824 & _guard825;
wire _guard827 = ~_guard0;
wire _guard828 = early_reset_static_par0_go_out;
wire _guard829 = _guard827 & _guard828;
wire _guard830 = early_reset_static_par0_go_out;
wire _guard831 = early_reset_static_par0_go_out;
wire _guard832 = ~_guard0;
wire _guard833 = early_reset_static_par0_go_out;
wire _guard834 = _guard832 & _guard833;
wire _guard835 = early_reset_static_par0_go_out;
wire _guard836 = ~_guard0;
wire _guard837 = early_reset_static_par0_go_out;
wire _guard838 = _guard836 & _guard837;
wire _guard839 = early_reset_static_par0_go_out;
wire _guard840 = ~_guard0;
wire _guard841 = early_reset_static_par0_go_out;
wire _guard842 = _guard840 & _guard841;
wire _guard843 = early_reset_static_par0_go_out;
wire _guard844 = early_reset_static_par0_go_out;
wire _guard845 = early_reset_static_par0_go_out;
wire _guard846 = ~_guard0;
wire _guard847 = early_reset_static_par0_go_out;
wire _guard848 = _guard846 & _guard847;
wire _guard849 = early_reset_static_par0_go_out;
wire _guard850 = early_reset_static_par0_go_out;
wire _guard851 = early_reset_static_par0_go_out;
wire _guard852 = early_reset_static_par0_go_out;
wire _guard853 = early_reset_static_par0_go_out;
wire _guard854 = early_reset_static_par0_go_out;
wire _guard855 = ~_guard0;
wire _guard856 = early_reset_static_par0_go_out;
wire _guard857 = _guard855 & _guard856;
wire _guard858 = early_reset_static_par0_go_out;
wire _guard859 = ~_guard0;
wire _guard860 = early_reset_static_par0_go_out;
wire _guard861 = _guard859 & _guard860;
wire _guard862 = early_reset_static_par0_go_out;
wire _guard863 = ~_guard0;
wire _guard864 = early_reset_static_par0_go_out;
wire _guard865 = _guard863 & _guard864;
wire _guard866 = early_reset_static_par0_go_out;
wire _guard867 = early_reset_static_par0_go_out;
wire _guard868 = ~_guard0;
wire _guard869 = early_reset_static_par0_go_out;
wire _guard870 = _guard868 & _guard869;
wire _guard871 = ~_guard0;
wire _guard872 = early_reset_static_par0_go_out;
wire _guard873 = _guard871 & _guard872;
wire _guard874 = early_reset_static_par0_go_out;
wire _guard875 = early_reset_static_par0_go_out;
wire _guard876 = early_reset_static_par0_go_out;
wire _guard877 = early_reset_static_par0_go_out;
wire _guard878 = early_reset_static_par0_go_out;
wire _guard879 = early_reset_static_par0_go_out;
wire _guard880 = ~_guard0;
wire _guard881 = early_reset_static_par0_go_out;
wire _guard882 = _guard880 & _guard881;
wire _guard883 = early_reset_static_par0_go_out;
wire _guard884 = ~_guard0;
wire _guard885 = early_reset_static_par0_go_out;
wire _guard886 = _guard884 & _guard885;
wire _guard887 = early_reset_static_par0_go_out;
wire _guard888 = early_reset_static_par0_go_out;
wire _guard889 = ~_guard0;
wire _guard890 = early_reset_static_par0_go_out;
wire _guard891 = _guard889 & _guard890;
wire _guard892 = early_reset_static_par0_go_out;
wire _guard893 = early_reset_static_par0_go_out;
wire _guard894 = ~_guard0;
wire _guard895 = early_reset_static_par0_go_out;
wire _guard896 = _guard894 & _guard895;
wire _guard897 = early_reset_static_par0_go_out;
wire _guard898 = early_reset_static_par0_go_out;
wire _guard899 = early_reset_static_par0_go_out;
wire _guard900 = early_reset_static_par0_go_out;
wire _guard901 = early_reset_static_par0_go_out;
wire _guard902 = ~_guard0;
wire _guard903 = early_reset_static_par0_go_out;
wire _guard904 = _guard902 & _guard903;
wire _guard905 = early_reset_static_par0_go_out;
wire _guard906 = early_reset_static_par0_go_out;
wire _guard907 = ~_guard0;
wire _guard908 = early_reset_static_par0_go_out;
wire _guard909 = _guard907 & _guard908;
wire _guard910 = early_reset_static_par0_go_out;
wire _guard911 = early_reset_static_par0_go_out;
wire _guard912 = early_reset_static_par0_go_out;
wire _guard913 = early_reset_static_par0_go_out;
wire _guard914 = early_reset_static_par0_go_out;
wire _guard915 = early_reset_static_par0_go_out;
wire _guard916 = early_reset_static_par0_go_out;
wire _guard917 = ~_guard0;
wire _guard918 = early_reset_static_par0_go_out;
wire _guard919 = _guard917 & _guard918;
wire _guard920 = early_reset_static_par0_go_out;
wire _guard921 = ~_guard0;
wire _guard922 = early_reset_static_par0_go_out;
wire _guard923 = _guard921 & _guard922;
wire _guard924 = early_reset_static_par0_go_out;
wire _guard925 = early_reset_static_par0_go_out;
wire _guard926 = ~_guard0;
wire _guard927 = early_reset_static_par0_go_out;
wire _guard928 = _guard926 & _guard927;
wire _guard929 = ~_guard0;
wire _guard930 = early_reset_static_par0_go_out;
wire _guard931 = _guard929 & _guard930;
wire _guard932 = early_reset_static_par0_go_out;
wire _guard933 = early_reset_static_par0_go_out;
wire _guard934 = ~_guard0;
wire _guard935 = early_reset_static_par0_go_out;
wire _guard936 = _guard934 & _guard935;
wire _guard937 = early_reset_static_par0_go_out;
wire _guard938 = ~_guard0;
wire _guard939 = early_reset_static_par0_go_out;
wire _guard940 = _guard938 & _guard939;
wire _guard941 = early_reset_static_par0_go_out;
wire _guard942 = ~_guard0;
wire _guard943 = early_reset_static_par0_go_out;
wire _guard944 = _guard942 & _guard943;
wire _guard945 = early_reset_static_par0_go_out;
wire _guard946 = early_reset_static_par0_go_out;
wire _guard947 = early_reset_static_par0_go_out;
wire _guard948 = early_reset_static_par0_go_out;
wire _guard949 = early_reset_static_par0_go_out;
wire _guard950 = early_reset_static_par0_go_out;
wire _guard951 = early_reset_static_par0_go_out;
wire _guard952 = early_reset_static_par0_go_out;
wire _guard953 = early_reset_static_par0_go_out;
wire _guard954 = early_reset_static_par0_go_out;
wire _guard955 = early_reset_static_par0_go_out;
wire _guard956 = ~_guard0;
wire _guard957 = early_reset_static_par0_go_out;
wire _guard958 = _guard956 & _guard957;
wire _guard959 = early_reset_static_par0_go_out;
wire _guard960 = ~_guard0;
wire _guard961 = early_reset_static_par0_go_out;
wire _guard962 = _guard960 & _guard961;
wire _guard963 = early_reset_static_par0_go_out;
wire _guard964 = ~_guard0;
wire _guard965 = early_reset_static_par0_go_out;
wire _guard966 = _guard964 & _guard965;
wire _guard967 = early_reset_static_par0_go_out;
wire _guard968 = ~_guard0;
wire _guard969 = early_reset_static_par0_go_out;
wire _guard970 = _guard968 & _guard969;
wire _guard971 = ~_guard0;
wire _guard972 = early_reset_static_par0_go_out;
wire _guard973 = _guard971 & _guard972;
wire _guard974 = early_reset_static_par0_go_out;
wire _guard975 = early_reset_static_par0_go_out;
wire _guard976 = early_reset_static_par0_go_out;
wire _guard977 = early_reset_static_par0_go_out;
wire _guard978 = ~_guard0;
wire _guard979 = early_reset_static_par0_go_out;
wire _guard980 = _guard978 & _guard979;
wire _guard981 = early_reset_static_par0_go_out;
wire _guard982 = ~_guard0;
wire _guard983 = early_reset_static_par0_go_out;
wire _guard984 = _guard982 & _guard983;
wire _guard985 = early_reset_static_par0_go_out;
wire _guard986 = early_reset_static_par0_go_out;
wire _guard987 = ~_guard0;
wire _guard988 = early_reset_static_par0_go_out;
wire _guard989 = _guard987 & _guard988;
wire _guard990 = early_reset_static_par0_go_out;
wire _guard991 = early_reset_static_par0_go_out;
wire _guard992 = early_reset_static_par0_go_out;
wire _guard993 = ~_guard0;
wire _guard994 = early_reset_static_par0_go_out;
wire _guard995 = _guard993 & _guard994;
wire _guard996 = early_reset_static_par0_go_out;
wire _guard997 = early_reset_static_par0_go_out;
wire _guard998 = early_reset_static_par0_go_out;
wire _guard999 = early_reset_static_par0_go_out;
wire _guard1000 = early_reset_static_par0_go_out;
wire _guard1001 = early_reset_static_par0_go_out;
wire _guard1002 = early_reset_static_par0_go_out;
wire _guard1003 = early_reset_static_par0_go_out;
wire _guard1004 = ~_guard0;
wire _guard1005 = early_reset_static_par0_go_out;
wire _guard1006 = _guard1004 & _guard1005;
wire _guard1007 = early_reset_static_par0_go_out;
wire _guard1008 = ~_guard0;
wire _guard1009 = early_reset_static_par0_go_out;
wire _guard1010 = _guard1008 & _guard1009;
wire _guard1011 = early_reset_static_par0_go_out;
wire _guard1012 = early_reset_static_par0_go_out;
wire _guard1013 = ~_guard0;
wire _guard1014 = early_reset_static_par0_go_out;
wire _guard1015 = _guard1013 & _guard1014;
wire _guard1016 = early_reset_static_par0_go_out;
wire _guard1017 = ~_guard0;
wire _guard1018 = early_reset_static_par0_go_out;
wire _guard1019 = _guard1017 & _guard1018;
wire _guard1020 = early_reset_static_par0_go_out;
wire _guard1021 = ~_guard0;
wire _guard1022 = early_reset_static_par0_go_out;
wire _guard1023 = _guard1021 & _guard1022;
wire _guard1024 = early_reset_static_par0_go_out;
wire _guard1025 = early_reset_static_par0_go_out;
wire _guard1026 = early_reset_static_par0_go_out;
wire _guard1027 = ~_guard0;
wire _guard1028 = early_reset_static_par0_go_out;
wire _guard1029 = _guard1027 & _guard1028;
wire _guard1030 = early_reset_static_par0_go_out;
wire _guard1031 = early_reset_static_par0_go_out;
wire _guard1032 = ~_guard0;
wire _guard1033 = early_reset_static_par0_go_out;
wire _guard1034 = _guard1032 & _guard1033;
wire _guard1035 = early_reset_static_par0_go_out;
wire _guard1036 = early_reset_static_par0_go_out;
wire _guard1037 = ~_guard0;
wire _guard1038 = early_reset_static_par0_go_out;
wire _guard1039 = _guard1037 & _guard1038;
wire _guard1040 = early_reset_static_par0_go_out;
wire _guard1041 = ~_guard0;
wire _guard1042 = early_reset_static_par0_go_out;
wire _guard1043 = _guard1041 & _guard1042;
wire _guard1044 = early_reset_static_par0_go_out;
wire _guard1045 = ~_guard0;
wire _guard1046 = early_reset_static_par0_go_out;
wire _guard1047 = _guard1045 & _guard1046;
wire _guard1048 = early_reset_static_par0_go_out;
wire _guard1049 = early_reset_static_par0_go_out;
wire _guard1050 = ~_guard0;
wire _guard1051 = early_reset_static_par0_go_out;
wire _guard1052 = _guard1050 & _guard1051;
wire _guard1053 = early_reset_static_par0_go_out;
wire _guard1054 = ~_guard0;
wire _guard1055 = early_reset_static_par0_go_out;
wire _guard1056 = _guard1054 & _guard1055;
wire _guard1057 = early_reset_static_par0_go_out;
wire _guard1058 = early_reset_static_par0_go_out;
wire _guard1059 = early_reset_static_par0_go_out;
wire _guard1060 = ~_guard0;
wire _guard1061 = early_reset_static_par0_go_out;
wire _guard1062 = _guard1060 & _guard1061;
wire _guard1063 = early_reset_static_par0_go_out;
wire _guard1064 = early_reset_static_par0_go_out;
wire _guard1065 = early_reset_static_par0_go_out;
wire _guard1066 = early_reset_static_par0_go_out;
wire _guard1067 = early_reset_static_par0_go_out;
wire _guard1068 = early_reset_static_par0_go_out;
wire _guard1069 = early_reset_static_par0_go_out;
wire _guard1070 = early_reset_static_par0_go_out;
wire _guard1071 = ~_guard0;
wire _guard1072 = early_reset_static_par0_go_out;
wire _guard1073 = _guard1071 & _guard1072;
wire _guard1074 = early_reset_static_par0_go_out;
wire _guard1075 = early_reset_static_par0_go_out;
wire _guard1076 = early_reset_static_par0_go_out;
wire _guard1077 = ~_guard0;
wire _guard1078 = early_reset_static_par0_go_out;
wire _guard1079 = _guard1077 & _guard1078;
wire _guard1080 = early_reset_static_par0_go_out;
wire _guard1081 = early_reset_static_par0_go_out;
wire _guard1082 = early_reset_static_par0_go_out;
wire _guard1083 = ~_guard0;
wire _guard1084 = early_reset_static_par0_go_out;
wire _guard1085 = _guard1083 & _guard1084;
wire _guard1086 = early_reset_static_par0_go_out;
wire _guard1087 = ~_guard0;
wire _guard1088 = early_reset_static_par0_go_out;
wire _guard1089 = _guard1087 & _guard1088;
wire _guard1090 = early_reset_static_par0_go_out;
wire _guard1091 = early_reset_static_par0_go_out;
wire _guard1092 = ~_guard0;
wire _guard1093 = early_reset_static_par0_go_out;
wire _guard1094 = _guard1092 & _guard1093;
wire _guard1095 = early_reset_static_par0_go_out;
wire _guard1096 = early_reset_static_par0_go_out;
wire _guard1097 = early_reset_static_par0_go_out;
wire _guard1098 = early_reset_static_par0_go_out;
wire _guard1099 = early_reset_static_par0_go_out;
wire _guard1100 = early_reset_static_par0_go_out;
wire _guard1101 = early_reset_static_par0_go_out;
wire _guard1102 = ~_guard0;
wire _guard1103 = early_reset_static_par0_go_out;
wire _guard1104 = _guard1102 & _guard1103;
wire _guard1105 = early_reset_static_par0_go_out;
wire _guard1106 = ~_guard0;
wire _guard1107 = early_reset_static_par0_go_out;
wire _guard1108 = _guard1106 & _guard1107;
wire _guard1109 = early_reset_static_par0_go_out;
wire _guard1110 = early_reset_static_par0_go_out;
wire _guard1111 = early_reset_static_par0_go_out;
wire _guard1112 = ~_guard0;
wire _guard1113 = early_reset_static_par0_go_out;
wire _guard1114 = _guard1112 & _guard1113;
wire _guard1115 = early_reset_static_par0_go_out;
wire _guard1116 = ~_guard0;
wire _guard1117 = early_reset_static_par0_go_out;
wire _guard1118 = _guard1116 & _guard1117;
wire _guard1119 = early_reset_static_par0_go_out;
wire _guard1120 = ~_guard0;
wire _guard1121 = early_reset_static_par0_go_out;
wire _guard1122 = _guard1120 & _guard1121;
wire _guard1123 = early_reset_static_par0_go_out;
wire _guard1124 = early_reset_static_par0_go_out;
wire _guard1125 = early_reset_static_par0_go_out;
wire _guard1126 = ~_guard0;
wire _guard1127 = early_reset_static_par0_go_out;
wire _guard1128 = _guard1126 & _guard1127;
wire _guard1129 = ~_guard0;
wire _guard1130 = early_reset_static_par0_go_out;
wire _guard1131 = _guard1129 & _guard1130;
wire _guard1132 = early_reset_static_par0_go_out;
wire _guard1133 = ~_guard0;
wire _guard1134 = early_reset_static_par0_go_out;
wire _guard1135 = _guard1133 & _guard1134;
wire _guard1136 = early_reset_static_par0_go_out;
wire _guard1137 = early_reset_static_par0_go_out;
wire _guard1138 = ~_guard0;
wire _guard1139 = early_reset_static_par0_go_out;
wire _guard1140 = _guard1138 & _guard1139;
wire _guard1141 = ~_guard0;
wire _guard1142 = early_reset_static_par0_go_out;
wire _guard1143 = _guard1141 & _guard1142;
wire _guard1144 = early_reset_static_par0_go_out;
wire _guard1145 = ~_guard0;
wire _guard1146 = early_reset_static_par0_go_out;
wire _guard1147 = _guard1145 & _guard1146;
wire _guard1148 = early_reset_static_par0_go_out;
wire _guard1149 = early_reset_static_par0_go_out;
wire _guard1150 = ~_guard0;
wire _guard1151 = early_reset_static_par0_go_out;
wire _guard1152 = _guard1150 & _guard1151;
wire _guard1153 = early_reset_static_par0_go_out;
wire _guard1154 = early_reset_static_par0_go_out;
wire _guard1155 = ~_guard0;
wire _guard1156 = early_reset_static_par0_go_out;
wire _guard1157 = _guard1155 & _guard1156;
wire _guard1158 = early_reset_static_par0_go_out;
wire _guard1159 = early_reset_static_par0_go_out;
wire _guard1160 = early_reset_static_par0_go_out;
wire _guard1161 = early_reset_static_par0_go_out;
wire _guard1162 = early_reset_static_par0_go_out;
wire _guard1163 = early_reset_static_par0_go_out;
wire _guard1164 = early_reset_static_par0_go_out;
wire _guard1165 = early_reset_static_par0_go_out;
wire _guard1166 = early_reset_static_par0_go_out;
wire _guard1167 = early_reset_static_par0_go_out;
wire _guard1168 = early_reset_static_par0_go_out;
wire _guard1169 = early_reset_static_par0_go_out;
wire _guard1170 = early_reset_static_par0_go_out;
wire _guard1171 = early_reset_static_par0_go_out;
wire _guard1172 = ~_guard0;
wire _guard1173 = early_reset_static_par0_go_out;
wire _guard1174 = _guard1172 & _guard1173;
wire _guard1175 = early_reset_static_par0_go_out;
wire _guard1176 = ~_guard0;
wire _guard1177 = early_reset_static_par0_go_out;
wire _guard1178 = _guard1176 & _guard1177;
wire _guard1179 = early_reset_static_par0_go_out;
wire _guard1180 = ~_guard0;
wire _guard1181 = early_reset_static_par0_go_out;
wire _guard1182 = _guard1180 & _guard1181;
wire _guard1183 = early_reset_static_par0_go_out;
wire _guard1184 = ~_guard0;
wire _guard1185 = early_reset_static_par0_go_out;
wire _guard1186 = _guard1184 & _guard1185;
wire _guard1187 = early_reset_static_par0_go_out;
wire _guard1188 = ~_guard0;
wire _guard1189 = early_reset_static_par0_go_out;
wire _guard1190 = _guard1188 & _guard1189;
wire _guard1191 = early_reset_static_par0_go_out;
wire _guard1192 = ~_guard0;
wire _guard1193 = early_reset_static_par0_go_out;
wire _guard1194 = _guard1192 & _guard1193;
wire _guard1195 = early_reset_static_par0_go_out;
wire _guard1196 = ~_guard0;
wire _guard1197 = early_reset_static_par0_go_out;
wire _guard1198 = _guard1196 & _guard1197;
wire _guard1199 = cond_wire11_out;
wire _guard1200 = early_reset_static_par0_go_out;
wire _guard1201 = _guard1199 & _guard1200;
wire _guard1202 = cond_wire11_out;
wire _guard1203 = early_reset_static_par0_go_out;
wire _guard1204 = _guard1202 & _guard1203;
wire _guard1205 = cond_wire16_out;
wire _guard1206 = early_reset_static_par0_go_out;
wire _guard1207 = _guard1205 & _guard1206;
wire _guard1208 = cond_wire16_out;
wire _guard1209 = early_reset_static_par0_go_out;
wire _guard1210 = _guard1208 & _guard1209;
wire _guard1211 = cond_wire52_out;
wire _guard1212 = early_reset_static_par0_go_out;
wire _guard1213 = _guard1211 & _guard1212;
wire _guard1214 = cond_wire50_out;
wire _guard1215 = early_reset_static_par0_go_out;
wire _guard1216 = _guard1214 & _guard1215;
wire _guard1217 = fsm_out == 1'd0;
wire _guard1218 = cond_wire50_out;
wire _guard1219 = _guard1217 & _guard1218;
wire _guard1220 = fsm_out == 1'd0;
wire _guard1221 = _guard1219 & _guard1220;
wire _guard1222 = fsm_out == 1'd0;
wire _guard1223 = cond_wire52_out;
wire _guard1224 = _guard1222 & _guard1223;
wire _guard1225 = fsm_out == 1'd0;
wire _guard1226 = _guard1224 & _guard1225;
wire _guard1227 = _guard1221 | _guard1226;
wire _guard1228 = early_reset_static_par0_go_out;
wire _guard1229 = _guard1227 & _guard1228;
wire _guard1230 = fsm_out == 1'd0;
wire _guard1231 = cond_wire50_out;
wire _guard1232 = _guard1230 & _guard1231;
wire _guard1233 = fsm_out == 1'd0;
wire _guard1234 = _guard1232 & _guard1233;
wire _guard1235 = fsm_out == 1'd0;
wire _guard1236 = cond_wire52_out;
wire _guard1237 = _guard1235 & _guard1236;
wire _guard1238 = fsm_out == 1'd0;
wire _guard1239 = _guard1237 & _guard1238;
wire _guard1240 = _guard1234 | _guard1239;
wire _guard1241 = early_reset_static_par0_go_out;
wire _guard1242 = _guard1240 & _guard1241;
wire _guard1243 = fsm_out == 1'd0;
wire _guard1244 = cond_wire50_out;
wire _guard1245 = _guard1243 & _guard1244;
wire _guard1246 = fsm_out == 1'd0;
wire _guard1247 = _guard1245 & _guard1246;
wire _guard1248 = fsm_out == 1'd0;
wire _guard1249 = cond_wire52_out;
wire _guard1250 = _guard1248 & _guard1249;
wire _guard1251 = fsm_out == 1'd0;
wire _guard1252 = _guard1250 & _guard1251;
wire _guard1253 = _guard1247 | _guard1252;
wire _guard1254 = early_reset_static_par0_go_out;
wire _guard1255 = _guard1253 & _guard1254;
wire _guard1256 = cond_wire1_out;
wire _guard1257 = early_reset_static_par0_go_out;
wire _guard1258 = _guard1256 & _guard1257;
wire _guard1259 = cond_wire1_out;
wire _guard1260 = early_reset_static_par0_go_out;
wire _guard1261 = _guard1259 & _guard1260;
wire _guard1262 = cond_wire90_out;
wire _guard1263 = early_reset_static_par0_go_out;
wire _guard1264 = _guard1262 & _guard1263;
wire _guard1265 = cond_wire88_out;
wire _guard1266 = early_reset_static_par0_go_out;
wire _guard1267 = _guard1265 & _guard1266;
wire _guard1268 = fsm_out == 1'd0;
wire _guard1269 = cond_wire88_out;
wire _guard1270 = _guard1268 & _guard1269;
wire _guard1271 = fsm_out == 1'd0;
wire _guard1272 = _guard1270 & _guard1271;
wire _guard1273 = fsm_out == 1'd0;
wire _guard1274 = cond_wire90_out;
wire _guard1275 = _guard1273 & _guard1274;
wire _guard1276 = fsm_out == 1'd0;
wire _guard1277 = _guard1275 & _guard1276;
wire _guard1278 = _guard1272 | _guard1277;
wire _guard1279 = early_reset_static_par0_go_out;
wire _guard1280 = _guard1278 & _guard1279;
wire _guard1281 = fsm_out == 1'd0;
wire _guard1282 = cond_wire88_out;
wire _guard1283 = _guard1281 & _guard1282;
wire _guard1284 = fsm_out == 1'd0;
wire _guard1285 = _guard1283 & _guard1284;
wire _guard1286 = fsm_out == 1'd0;
wire _guard1287 = cond_wire90_out;
wire _guard1288 = _guard1286 & _guard1287;
wire _guard1289 = fsm_out == 1'd0;
wire _guard1290 = _guard1288 & _guard1289;
wire _guard1291 = _guard1285 | _guard1290;
wire _guard1292 = early_reset_static_par0_go_out;
wire _guard1293 = _guard1291 & _guard1292;
wire _guard1294 = fsm_out == 1'd0;
wire _guard1295 = cond_wire88_out;
wire _guard1296 = _guard1294 & _guard1295;
wire _guard1297 = fsm_out == 1'd0;
wire _guard1298 = _guard1296 & _guard1297;
wire _guard1299 = fsm_out == 1'd0;
wire _guard1300 = cond_wire90_out;
wire _guard1301 = _guard1299 & _guard1300;
wire _guard1302 = fsm_out == 1'd0;
wire _guard1303 = _guard1301 & _guard1302;
wire _guard1304 = _guard1298 | _guard1303;
wire _guard1305 = early_reset_static_par0_go_out;
wire _guard1306 = _guard1304 & _guard1305;
wire _guard1307 = cond_wire94_out;
wire _guard1308 = early_reset_static_par0_go_out;
wire _guard1309 = _guard1307 & _guard1308;
wire _guard1310 = cond_wire92_out;
wire _guard1311 = early_reset_static_par0_go_out;
wire _guard1312 = _guard1310 & _guard1311;
wire _guard1313 = fsm_out == 1'd0;
wire _guard1314 = cond_wire92_out;
wire _guard1315 = _guard1313 & _guard1314;
wire _guard1316 = fsm_out == 1'd0;
wire _guard1317 = _guard1315 & _guard1316;
wire _guard1318 = fsm_out == 1'd0;
wire _guard1319 = cond_wire94_out;
wire _guard1320 = _guard1318 & _guard1319;
wire _guard1321 = fsm_out == 1'd0;
wire _guard1322 = _guard1320 & _guard1321;
wire _guard1323 = _guard1317 | _guard1322;
wire _guard1324 = early_reset_static_par0_go_out;
wire _guard1325 = _guard1323 & _guard1324;
wire _guard1326 = fsm_out == 1'd0;
wire _guard1327 = cond_wire92_out;
wire _guard1328 = _guard1326 & _guard1327;
wire _guard1329 = fsm_out == 1'd0;
wire _guard1330 = _guard1328 & _guard1329;
wire _guard1331 = fsm_out == 1'd0;
wire _guard1332 = cond_wire94_out;
wire _guard1333 = _guard1331 & _guard1332;
wire _guard1334 = fsm_out == 1'd0;
wire _guard1335 = _guard1333 & _guard1334;
wire _guard1336 = _guard1330 | _guard1335;
wire _guard1337 = early_reset_static_par0_go_out;
wire _guard1338 = _guard1336 & _guard1337;
wire _guard1339 = fsm_out == 1'd0;
wire _guard1340 = cond_wire92_out;
wire _guard1341 = _guard1339 & _guard1340;
wire _guard1342 = fsm_out == 1'd0;
wire _guard1343 = _guard1341 & _guard1342;
wire _guard1344 = fsm_out == 1'd0;
wire _guard1345 = cond_wire94_out;
wire _guard1346 = _guard1344 & _guard1345;
wire _guard1347 = fsm_out == 1'd0;
wire _guard1348 = _guard1346 & _guard1347;
wire _guard1349 = _guard1343 | _guard1348;
wire _guard1350 = early_reset_static_par0_go_out;
wire _guard1351 = _guard1349 & _guard1350;
wire _guard1352 = cond_wire89_out;
wire _guard1353 = early_reset_static_par0_go_out;
wire _guard1354 = _guard1352 & _guard1353;
wire _guard1355 = cond_wire89_out;
wire _guard1356 = early_reset_static_par0_go_out;
wire _guard1357 = _guard1355 & _guard1356;
wire _guard1358 = cond_wire66_out;
wire _guard1359 = early_reset_static_par0_go_out;
wire _guard1360 = _guard1358 & _guard1359;
wire _guard1361 = cond_wire66_out;
wire _guard1362 = early_reset_static_par0_go_out;
wire _guard1363 = _guard1361 & _guard1362;
wire _guard1364 = cond_wire133_out;
wire _guard1365 = early_reset_static_par0_go_out;
wire _guard1366 = _guard1364 & _guard1365;
wire _guard1367 = cond_wire133_out;
wire _guard1368 = early_reset_static_par0_go_out;
wire _guard1369 = _guard1367 & _guard1368;
wire _guard1370 = cond_wire166_out;
wire _guard1371 = early_reset_static_par0_go_out;
wire _guard1372 = _guard1370 & _guard1371;
wire _guard1373 = cond_wire166_out;
wire _guard1374 = early_reset_static_par0_go_out;
wire _guard1375 = _guard1373 & _guard1374;
wire _guard1376 = cond_wire174_out;
wire _guard1377 = early_reset_static_par0_go_out;
wire _guard1378 = _guard1376 & _guard1377;
wire _guard1379 = cond_wire174_out;
wire _guard1380 = early_reset_static_par0_go_out;
wire _guard1381 = _guard1379 & _guard1380;
wire _guard1382 = cond_wire191_out;
wire _guard1383 = early_reset_static_par0_go_out;
wire _guard1384 = _guard1382 & _guard1383;
wire _guard1385 = cond_wire189_out;
wire _guard1386 = early_reset_static_par0_go_out;
wire _guard1387 = _guard1385 & _guard1386;
wire _guard1388 = fsm_out == 1'd0;
wire _guard1389 = cond_wire189_out;
wire _guard1390 = _guard1388 & _guard1389;
wire _guard1391 = fsm_out == 1'd0;
wire _guard1392 = _guard1390 & _guard1391;
wire _guard1393 = fsm_out == 1'd0;
wire _guard1394 = cond_wire191_out;
wire _guard1395 = _guard1393 & _guard1394;
wire _guard1396 = fsm_out == 1'd0;
wire _guard1397 = _guard1395 & _guard1396;
wire _guard1398 = _guard1392 | _guard1397;
wire _guard1399 = early_reset_static_par0_go_out;
wire _guard1400 = _guard1398 & _guard1399;
wire _guard1401 = fsm_out == 1'd0;
wire _guard1402 = cond_wire189_out;
wire _guard1403 = _guard1401 & _guard1402;
wire _guard1404 = fsm_out == 1'd0;
wire _guard1405 = _guard1403 & _guard1404;
wire _guard1406 = fsm_out == 1'd0;
wire _guard1407 = cond_wire191_out;
wire _guard1408 = _guard1406 & _guard1407;
wire _guard1409 = fsm_out == 1'd0;
wire _guard1410 = _guard1408 & _guard1409;
wire _guard1411 = _guard1405 | _guard1410;
wire _guard1412 = early_reset_static_par0_go_out;
wire _guard1413 = _guard1411 & _guard1412;
wire _guard1414 = fsm_out == 1'd0;
wire _guard1415 = cond_wire189_out;
wire _guard1416 = _guard1414 & _guard1415;
wire _guard1417 = fsm_out == 1'd0;
wire _guard1418 = _guard1416 & _guard1417;
wire _guard1419 = fsm_out == 1'd0;
wire _guard1420 = cond_wire191_out;
wire _guard1421 = _guard1419 & _guard1420;
wire _guard1422 = fsm_out == 1'd0;
wire _guard1423 = _guard1421 & _guard1422;
wire _guard1424 = _guard1418 | _guard1423;
wire _guard1425 = early_reset_static_par0_go_out;
wire _guard1426 = _guard1424 & _guard1425;
wire _guard1427 = cond_wire239_out;
wire _guard1428 = early_reset_static_par0_go_out;
wire _guard1429 = _guard1427 & _guard1428;
wire _guard1430 = cond_wire239_out;
wire _guard1431 = early_reset_static_par0_go_out;
wire _guard1432 = _guard1430 & _guard1431;
wire _guard1433 = cond_wire341_out;
wire _guard1434 = early_reset_static_par0_go_out;
wire _guard1435 = _guard1433 & _guard1434;
wire _guard1436 = cond_wire341_out;
wire _guard1437 = early_reset_static_par0_go_out;
wire _guard1438 = _guard1436 & _guard1437;
wire _guard1439 = cond_wire349_out;
wire _guard1440 = early_reset_static_par0_go_out;
wire _guard1441 = _guard1439 & _guard1440;
wire _guard1442 = cond_wire349_out;
wire _guard1443 = early_reset_static_par0_go_out;
wire _guard1444 = _guard1442 & _guard1443;
wire _guard1445 = cond_wire374_out;
wire _guard1446 = early_reset_static_par0_go_out;
wire _guard1447 = _guard1445 & _guard1446;
wire _guard1448 = cond_wire372_out;
wire _guard1449 = early_reset_static_par0_go_out;
wire _guard1450 = _guard1448 & _guard1449;
wire _guard1451 = fsm_out == 1'd0;
wire _guard1452 = cond_wire372_out;
wire _guard1453 = _guard1451 & _guard1452;
wire _guard1454 = fsm_out == 1'd0;
wire _guard1455 = _guard1453 & _guard1454;
wire _guard1456 = fsm_out == 1'd0;
wire _guard1457 = cond_wire374_out;
wire _guard1458 = _guard1456 & _guard1457;
wire _guard1459 = fsm_out == 1'd0;
wire _guard1460 = _guard1458 & _guard1459;
wire _guard1461 = _guard1455 | _guard1460;
wire _guard1462 = early_reset_static_par0_go_out;
wire _guard1463 = _guard1461 & _guard1462;
wire _guard1464 = fsm_out == 1'd0;
wire _guard1465 = cond_wire372_out;
wire _guard1466 = _guard1464 & _guard1465;
wire _guard1467 = fsm_out == 1'd0;
wire _guard1468 = _guard1466 & _guard1467;
wire _guard1469 = fsm_out == 1'd0;
wire _guard1470 = cond_wire374_out;
wire _guard1471 = _guard1469 & _guard1470;
wire _guard1472 = fsm_out == 1'd0;
wire _guard1473 = _guard1471 & _guard1472;
wire _guard1474 = _guard1468 | _guard1473;
wire _guard1475 = early_reset_static_par0_go_out;
wire _guard1476 = _guard1474 & _guard1475;
wire _guard1477 = fsm_out == 1'd0;
wire _guard1478 = cond_wire372_out;
wire _guard1479 = _guard1477 & _guard1478;
wire _guard1480 = fsm_out == 1'd0;
wire _guard1481 = _guard1479 & _guard1480;
wire _guard1482 = fsm_out == 1'd0;
wire _guard1483 = cond_wire374_out;
wire _guard1484 = _guard1482 & _guard1483;
wire _guard1485 = fsm_out == 1'd0;
wire _guard1486 = _guard1484 & _guard1485;
wire _guard1487 = _guard1481 | _guard1486;
wire _guard1488 = early_reset_static_par0_go_out;
wire _guard1489 = _guard1487 & _guard1488;
wire _guard1490 = cond_wire394_out;
wire _guard1491 = early_reset_static_par0_go_out;
wire _guard1492 = _guard1490 & _guard1491;
wire _guard1493 = cond_wire392_out;
wire _guard1494 = early_reset_static_par0_go_out;
wire _guard1495 = _guard1493 & _guard1494;
wire _guard1496 = fsm_out == 1'd0;
wire _guard1497 = cond_wire392_out;
wire _guard1498 = _guard1496 & _guard1497;
wire _guard1499 = fsm_out == 1'd0;
wire _guard1500 = _guard1498 & _guard1499;
wire _guard1501 = fsm_out == 1'd0;
wire _guard1502 = cond_wire394_out;
wire _guard1503 = _guard1501 & _guard1502;
wire _guard1504 = fsm_out == 1'd0;
wire _guard1505 = _guard1503 & _guard1504;
wire _guard1506 = _guard1500 | _guard1505;
wire _guard1507 = early_reset_static_par0_go_out;
wire _guard1508 = _guard1506 & _guard1507;
wire _guard1509 = fsm_out == 1'd0;
wire _guard1510 = cond_wire392_out;
wire _guard1511 = _guard1509 & _guard1510;
wire _guard1512 = fsm_out == 1'd0;
wire _guard1513 = _guard1511 & _guard1512;
wire _guard1514 = fsm_out == 1'd0;
wire _guard1515 = cond_wire394_out;
wire _guard1516 = _guard1514 & _guard1515;
wire _guard1517 = fsm_out == 1'd0;
wire _guard1518 = _guard1516 & _guard1517;
wire _guard1519 = _guard1513 | _guard1518;
wire _guard1520 = early_reset_static_par0_go_out;
wire _guard1521 = _guard1519 & _guard1520;
wire _guard1522 = fsm_out == 1'd0;
wire _guard1523 = cond_wire392_out;
wire _guard1524 = _guard1522 & _guard1523;
wire _guard1525 = fsm_out == 1'd0;
wire _guard1526 = _guard1524 & _guard1525;
wire _guard1527 = fsm_out == 1'd0;
wire _guard1528 = cond_wire394_out;
wire _guard1529 = _guard1527 & _guard1528;
wire _guard1530 = fsm_out == 1'd0;
wire _guard1531 = _guard1529 & _guard1530;
wire _guard1532 = _guard1526 | _guard1531;
wire _guard1533 = early_reset_static_par0_go_out;
wire _guard1534 = _guard1532 & _guard1533;
wire _guard1535 = cond_wire332_out;
wire _guard1536 = early_reset_static_par0_go_out;
wire _guard1537 = _guard1535 & _guard1536;
wire _guard1538 = cond_wire332_out;
wire _guard1539 = early_reset_static_par0_go_out;
wire _guard1540 = _guard1538 & _guard1539;
wire _guard1541 = cond_wire423_out;
wire _guard1542 = early_reset_static_par0_go_out;
wire _guard1543 = _guard1541 & _guard1542;
wire _guard1544 = cond_wire421_out;
wire _guard1545 = early_reset_static_par0_go_out;
wire _guard1546 = _guard1544 & _guard1545;
wire _guard1547 = fsm_out == 1'd0;
wire _guard1548 = cond_wire421_out;
wire _guard1549 = _guard1547 & _guard1548;
wire _guard1550 = fsm_out == 1'd0;
wire _guard1551 = _guard1549 & _guard1550;
wire _guard1552 = fsm_out == 1'd0;
wire _guard1553 = cond_wire423_out;
wire _guard1554 = _guard1552 & _guard1553;
wire _guard1555 = fsm_out == 1'd0;
wire _guard1556 = _guard1554 & _guard1555;
wire _guard1557 = _guard1551 | _guard1556;
wire _guard1558 = early_reset_static_par0_go_out;
wire _guard1559 = _guard1557 & _guard1558;
wire _guard1560 = fsm_out == 1'd0;
wire _guard1561 = cond_wire421_out;
wire _guard1562 = _guard1560 & _guard1561;
wire _guard1563 = fsm_out == 1'd0;
wire _guard1564 = _guard1562 & _guard1563;
wire _guard1565 = fsm_out == 1'd0;
wire _guard1566 = cond_wire423_out;
wire _guard1567 = _guard1565 & _guard1566;
wire _guard1568 = fsm_out == 1'd0;
wire _guard1569 = _guard1567 & _guard1568;
wire _guard1570 = _guard1564 | _guard1569;
wire _guard1571 = early_reset_static_par0_go_out;
wire _guard1572 = _guard1570 & _guard1571;
wire _guard1573 = fsm_out == 1'd0;
wire _guard1574 = cond_wire421_out;
wire _guard1575 = _guard1573 & _guard1574;
wire _guard1576 = fsm_out == 1'd0;
wire _guard1577 = _guard1575 & _guard1576;
wire _guard1578 = fsm_out == 1'd0;
wire _guard1579 = cond_wire423_out;
wire _guard1580 = _guard1578 & _guard1579;
wire _guard1581 = fsm_out == 1'd0;
wire _guard1582 = _guard1580 & _guard1581;
wire _guard1583 = _guard1577 | _guard1582;
wire _guard1584 = early_reset_static_par0_go_out;
wire _guard1585 = _guard1583 & _guard1584;
wire _guard1586 = cond_wire369_out;
wire _guard1587 = early_reset_static_par0_go_out;
wire _guard1588 = _guard1586 & _guard1587;
wire _guard1589 = cond_wire369_out;
wire _guard1590 = early_reset_static_par0_go_out;
wire _guard1591 = _guard1589 & _guard1590;
wire _guard1592 = cond_wire450_out;
wire _guard1593 = early_reset_static_par0_go_out;
wire _guard1594 = _guard1592 & _guard1593;
wire _guard1595 = cond_wire450_out;
wire _guard1596 = early_reset_static_par0_go_out;
wire _guard1597 = _guard1595 & _guard1596;
wire _guard1598 = cond_wire484_out;
wire _guard1599 = early_reset_static_par0_go_out;
wire _guard1600 = _guard1598 & _guard1599;
wire _guard1601 = cond_wire482_out;
wire _guard1602 = early_reset_static_par0_go_out;
wire _guard1603 = _guard1601 & _guard1602;
wire _guard1604 = fsm_out == 1'd0;
wire _guard1605 = cond_wire482_out;
wire _guard1606 = _guard1604 & _guard1605;
wire _guard1607 = fsm_out == 1'd0;
wire _guard1608 = _guard1606 & _guard1607;
wire _guard1609 = fsm_out == 1'd0;
wire _guard1610 = cond_wire484_out;
wire _guard1611 = _guard1609 & _guard1610;
wire _guard1612 = fsm_out == 1'd0;
wire _guard1613 = _guard1611 & _guard1612;
wire _guard1614 = _guard1608 | _guard1613;
wire _guard1615 = early_reset_static_par0_go_out;
wire _guard1616 = _guard1614 & _guard1615;
wire _guard1617 = fsm_out == 1'd0;
wire _guard1618 = cond_wire482_out;
wire _guard1619 = _guard1617 & _guard1618;
wire _guard1620 = fsm_out == 1'd0;
wire _guard1621 = _guard1619 & _guard1620;
wire _guard1622 = fsm_out == 1'd0;
wire _guard1623 = cond_wire484_out;
wire _guard1624 = _guard1622 & _guard1623;
wire _guard1625 = fsm_out == 1'd0;
wire _guard1626 = _guard1624 & _guard1625;
wire _guard1627 = _guard1621 | _guard1626;
wire _guard1628 = early_reset_static_par0_go_out;
wire _guard1629 = _guard1627 & _guard1628;
wire _guard1630 = fsm_out == 1'd0;
wire _guard1631 = cond_wire482_out;
wire _guard1632 = _guard1630 & _guard1631;
wire _guard1633 = fsm_out == 1'd0;
wire _guard1634 = _guard1632 & _guard1633;
wire _guard1635 = fsm_out == 1'd0;
wire _guard1636 = cond_wire484_out;
wire _guard1637 = _guard1635 & _guard1636;
wire _guard1638 = fsm_out == 1'd0;
wire _guard1639 = _guard1637 & _guard1638;
wire _guard1640 = _guard1634 | _guard1639;
wire _guard1641 = early_reset_static_par0_go_out;
wire _guard1642 = _guard1640 & _guard1641;
wire _guard1643 = cond_wire483_out;
wire _guard1644 = early_reset_static_par0_go_out;
wire _guard1645 = _guard1643 & _guard1644;
wire _guard1646 = cond_wire483_out;
wire _guard1647 = early_reset_static_par0_go_out;
wire _guard1648 = _guard1646 & _guard1647;
wire _guard1649 = cond_wire491_out;
wire _guard1650 = early_reset_static_par0_go_out;
wire _guard1651 = _guard1649 & _guard1650;
wire _guard1652 = cond_wire491_out;
wire _guard1653 = early_reset_static_par0_go_out;
wire _guard1654 = _guard1652 & _guard1653;
wire _guard1655 = cond_wire434_out;
wire _guard1656 = early_reset_static_par0_go_out;
wire _guard1657 = _guard1655 & _guard1656;
wire _guard1658 = cond_wire434_out;
wire _guard1659 = early_reset_static_par0_go_out;
wire _guard1660 = _guard1658 & _guard1659;
wire _guard1661 = cond_wire503_out;
wire _guard1662 = early_reset_static_par0_go_out;
wire _guard1663 = _guard1661 & _guard1662;
wire _guard1664 = cond_wire503_out;
wire _guard1665 = early_reset_static_par0_go_out;
wire _guard1666 = _guard1664 & _guard1665;
wire _guard1667 = cond_wire479_out;
wire _guard1668 = early_reset_static_par0_go_out;
wire _guard1669 = _guard1667 & _guard1668;
wire _guard1670 = cond_wire479_out;
wire _guard1671 = early_reset_static_par0_go_out;
wire _guard1672 = _guard1670 & _guard1671;
wire _guard1673 = cond_wire561_out;
wire _guard1674 = early_reset_static_par0_go_out;
wire _guard1675 = _guard1673 & _guard1674;
wire _guard1676 = cond_wire559_out;
wire _guard1677 = early_reset_static_par0_go_out;
wire _guard1678 = _guard1676 & _guard1677;
wire _guard1679 = fsm_out == 1'd0;
wire _guard1680 = cond_wire559_out;
wire _guard1681 = _guard1679 & _guard1680;
wire _guard1682 = fsm_out == 1'd0;
wire _guard1683 = _guard1681 & _guard1682;
wire _guard1684 = fsm_out == 1'd0;
wire _guard1685 = cond_wire561_out;
wire _guard1686 = _guard1684 & _guard1685;
wire _guard1687 = fsm_out == 1'd0;
wire _guard1688 = _guard1686 & _guard1687;
wire _guard1689 = _guard1683 | _guard1688;
wire _guard1690 = early_reset_static_par0_go_out;
wire _guard1691 = _guard1689 & _guard1690;
wire _guard1692 = fsm_out == 1'd0;
wire _guard1693 = cond_wire559_out;
wire _guard1694 = _guard1692 & _guard1693;
wire _guard1695 = fsm_out == 1'd0;
wire _guard1696 = _guard1694 & _guard1695;
wire _guard1697 = fsm_out == 1'd0;
wire _guard1698 = cond_wire561_out;
wire _guard1699 = _guard1697 & _guard1698;
wire _guard1700 = fsm_out == 1'd0;
wire _guard1701 = _guard1699 & _guard1700;
wire _guard1702 = _guard1696 | _guard1701;
wire _guard1703 = early_reset_static_par0_go_out;
wire _guard1704 = _guard1702 & _guard1703;
wire _guard1705 = fsm_out == 1'd0;
wire _guard1706 = cond_wire559_out;
wire _guard1707 = _guard1705 & _guard1706;
wire _guard1708 = fsm_out == 1'd0;
wire _guard1709 = _guard1707 & _guard1708;
wire _guard1710 = fsm_out == 1'd0;
wire _guard1711 = cond_wire561_out;
wire _guard1712 = _guard1710 & _guard1711;
wire _guard1713 = fsm_out == 1'd0;
wire _guard1714 = _guard1712 & _guard1713;
wire _guard1715 = _guard1709 | _guard1714;
wire _guard1716 = early_reset_static_par0_go_out;
wire _guard1717 = _guard1715 & _guard1716;
wire _guard1718 = cond_wire495_out;
wire _guard1719 = early_reset_static_par0_go_out;
wire _guard1720 = _guard1718 & _guard1719;
wire _guard1721 = cond_wire495_out;
wire _guard1722 = early_reset_static_par0_go_out;
wire _guard1723 = _guard1721 & _guard1722;
wire _guard1724 = cond_wire511_out;
wire _guard1725 = early_reset_static_par0_go_out;
wire _guard1726 = _guard1724 & _guard1725;
wire _guard1727 = cond_wire511_out;
wire _guard1728 = early_reset_static_par0_go_out;
wire _guard1729 = _guard1727 & _guard1728;
wire _guard1730 = cond_wire588_out;
wire _guard1731 = early_reset_static_par0_go_out;
wire _guard1732 = _guard1730 & _guard1731;
wire _guard1733 = cond_wire588_out;
wire _guard1734 = early_reset_static_par0_go_out;
wire _guard1735 = _guard1733 & _guard1734;
wire _guard1736 = cond_wire592_out;
wire _guard1737 = early_reset_static_par0_go_out;
wire _guard1738 = _guard1736 & _guard1737;
wire _guard1739 = cond_wire592_out;
wire _guard1740 = early_reset_static_par0_go_out;
wire _guard1741 = _guard1739 & _guard1740;
wire _guard1742 = cond_wire614_out;
wire _guard1743 = early_reset_static_par0_go_out;
wire _guard1744 = _guard1742 & _guard1743;
wire _guard1745 = cond_wire612_out;
wire _guard1746 = early_reset_static_par0_go_out;
wire _guard1747 = _guard1745 & _guard1746;
wire _guard1748 = fsm_out == 1'd0;
wire _guard1749 = cond_wire612_out;
wire _guard1750 = _guard1748 & _guard1749;
wire _guard1751 = fsm_out == 1'd0;
wire _guard1752 = _guard1750 & _guard1751;
wire _guard1753 = fsm_out == 1'd0;
wire _guard1754 = cond_wire614_out;
wire _guard1755 = _guard1753 & _guard1754;
wire _guard1756 = fsm_out == 1'd0;
wire _guard1757 = _guard1755 & _guard1756;
wire _guard1758 = _guard1752 | _guard1757;
wire _guard1759 = early_reset_static_par0_go_out;
wire _guard1760 = _guard1758 & _guard1759;
wire _guard1761 = fsm_out == 1'd0;
wire _guard1762 = cond_wire612_out;
wire _guard1763 = _guard1761 & _guard1762;
wire _guard1764 = fsm_out == 1'd0;
wire _guard1765 = _guard1763 & _guard1764;
wire _guard1766 = fsm_out == 1'd0;
wire _guard1767 = cond_wire614_out;
wire _guard1768 = _guard1766 & _guard1767;
wire _guard1769 = fsm_out == 1'd0;
wire _guard1770 = _guard1768 & _guard1769;
wire _guard1771 = _guard1765 | _guard1770;
wire _guard1772 = early_reset_static_par0_go_out;
wire _guard1773 = _guard1771 & _guard1772;
wire _guard1774 = fsm_out == 1'd0;
wire _guard1775 = cond_wire612_out;
wire _guard1776 = _guard1774 & _guard1775;
wire _guard1777 = fsm_out == 1'd0;
wire _guard1778 = _guard1776 & _guard1777;
wire _guard1779 = fsm_out == 1'd0;
wire _guard1780 = cond_wire614_out;
wire _guard1781 = _guard1779 & _guard1780;
wire _guard1782 = fsm_out == 1'd0;
wire _guard1783 = _guard1781 & _guard1782;
wire _guard1784 = _guard1778 | _guard1783;
wire _guard1785 = early_reset_static_par0_go_out;
wire _guard1786 = _guard1784 & _guard1785;
wire _guard1787 = cond_wire646_out;
wire _guard1788 = early_reset_static_par0_go_out;
wire _guard1789 = _guard1787 & _guard1788;
wire _guard1790 = cond_wire644_out;
wire _guard1791 = early_reset_static_par0_go_out;
wire _guard1792 = _guard1790 & _guard1791;
wire _guard1793 = fsm_out == 1'd0;
wire _guard1794 = cond_wire644_out;
wire _guard1795 = _guard1793 & _guard1794;
wire _guard1796 = fsm_out == 1'd0;
wire _guard1797 = _guard1795 & _guard1796;
wire _guard1798 = fsm_out == 1'd0;
wire _guard1799 = cond_wire646_out;
wire _guard1800 = _guard1798 & _guard1799;
wire _guard1801 = fsm_out == 1'd0;
wire _guard1802 = _guard1800 & _guard1801;
wire _guard1803 = _guard1797 | _guard1802;
wire _guard1804 = early_reset_static_par0_go_out;
wire _guard1805 = _guard1803 & _guard1804;
wire _guard1806 = fsm_out == 1'd0;
wire _guard1807 = cond_wire644_out;
wire _guard1808 = _guard1806 & _guard1807;
wire _guard1809 = fsm_out == 1'd0;
wire _guard1810 = _guard1808 & _guard1809;
wire _guard1811 = fsm_out == 1'd0;
wire _guard1812 = cond_wire646_out;
wire _guard1813 = _guard1811 & _guard1812;
wire _guard1814 = fsm_out == 1'd0;
wire _guard1815 = _guard1813 & _guard1814;
wire _guard1816 = _guard1810 | _guard1815;
wire _guard1817 = early_reset_static_par0_go_out;
wire _guard1818 = _guard1816 & _guard1817;
wire _guard1819 = fsm_out == 1'd0;
wire _guard1820 = cond_wire644_out;
wire _guard1821 = _guard1819 & _guard1820;
wire _guard1822 = fsm_out == 1'd0;
wire _guard1823 = _guard1821 & _guard1822;
wire _guard1824 = fsm_out == 1'd0;
wire _guard1825 = cond_wire646_out;
wire _guard1826 = _guard1824 & _guard1825;
wire _guard1827 = fsm_out == 1'd0;
wire _guard1828 = _guard1826 & _guard1827;
wire _guard1829 = _guard1823 | _guard1828;
wire _guard1830 = early_reset_static_par0_go_out;
wire _guard1831 = _guard1829 & _guard1830;
wire _guard1832 = cond_wire649_out;
wire _guard1833 = early_reset_static_par0_go_out;
wire _guard1834 = _guard1832 & _guard1833;
wire _guard1835 = cond_wire649_out;
wire _guard1836 = early_reset_static_par0_go_out;
wire _guard1837 = _guard1835 & _guard1836;
wire _guard1838 = cond_wire592_out;
wire _guard1839 = early_reset_static_par0_go_out;
wire _guard1840 = _guard1838 & _guard1839;
wire _guard1841 = cond_wire592_out;
wire _guard1842 = early_reset_static_par0_go_out;
wire _guard1843 = _guard1841 & _guard1842;
wire _guard1844 = cond_wire664_out;
wire _guard1845 = early_reset_static_par0_go_out;
wire _guard1846 = _guard1844 & _guard1845;
wire _guard1847 = cond_wire664_out;
wire _guard1848 = early_reset_static_par0_go_out;
wire _guard1849 = _guard1847 & _guard1848;
wire _guard1850 = cond_wire678_out;
wire _guard1851 = early_reset_static_par0_go_out;
wire _guard1852 = _guard1850 & _guard1851;
wire _guard1853 = cond_wire678_out;
wire _guard1854 = early_reset_static_par0_go_out;
wire _guard1855 = _guard1853 & _guard1854;
wire _guard1856 = cond_wire629_out;
wire _guard1857 = early_reset_static_par0_go_out;
wire _guard1858 = _guard1856 & _guard1857;
wire _guard1859 = cond_wire629_out;
wire _guard1860 = early_reset_static_par0_go_out;
wire _guard1861 = _guard1859 & _guard1860;
wire _guard1862 = cond_wire735_out;
wire _guard1863 = early_reset_static_par0_go_out;
wire _guard1864 = _guard1862 & _guard1863;
wire _guard1865 = cond_wire735_out;
wire _guard1866 = early_reset_static_par0_go_out;
wire _guard1867 = _guard1865 & _guard1866;
wire _guard1868 = cond_wire752_out;
wire _guard1869 = early_reset_static_par0_go_out;
wire _guard1870 = _guard1868 & _guard1869;
wire _guard1871 = cond_wire750_out;
wire _guard1872 = early_reset_static_par0_go_out;
wire _guard1873 = _guard1871 & _guard1872;
wire _guard1874 = fsm_out == 1'd0;
wire _guard1875 = cond_wire750_out;
wire _guard1876 = _guard1874 & _guard1875;
wire _guard1877 = fsm_out == 1'd0;
wire _guard1878 = _guard1876 & _guard1877;
wire _guard1879 = fsm_out == 1'd0;
wire _guard1880 = cond_wire752_out;
wire _guard1881 = _guard1879 & _guard1880;
wire _guard1882 = fsm_out == 1'd0;
wire _guard1883 = _guard1881 & _guard1882;
wire _guard1884 = _guard1878 | _guard1883;
wire _guard1885 = early_reset_static_par0_go_out;
wire _guard1886 = _guard1884 & _guard1885;
wire _guard1887 = fsm_out == 1'd0;
wire _guard1888 = cond_wire750_out;
wire _guard1889 = _guard1887 & _guard1888;
wire _guard1890 = fsm_out == 1'd0;
wire _guard1891 = _guard1889 & _guard1890;
wire _guard1892 = fsm_out == 1'd0;
wire _guard1893 = cond_wire752_out;
wire _guard1894 = _guard1892 & _guard1893;
wire _guard1895 = fsm_out == 1'd0;
wire _guard1896 = _guard1894 & _guard1895;
wire _guard1897 = _guard1891 | _guard1896;
wire _guard1898 = early_reset_static_par0_go_out;
wire _guard1899 = _guard1897 & _guard1898;
wire _guard1900 = fsm_out == 1'd0;
wire _guard1901 = cond_wire750_out;
wire _guard1902 = _guard1900 & _guard1901;
wire _guard1903 = fsm_out == 1'd0;
wire _guard1904 = _guard1902 & _guard1903;
wire _guard1905 = fsm_out == 1'd0;
wire _guard1906 = cond_wire752_out;
wire _guard1907 = _guard1905 & _guard1906;
wire _guard1908 = fsm_out == 1'd0;
wire _guard1909 = _guard1907 & _guard1908;
wire _guard1910 = _guard1904 | _guard1909;
wire _guard1911 = early_reset_static_par0_go_out;
wire _guard1912 = _guard1910 & _guard1911;
wire _guard1913 = cond_wire747_out;
wire _guard1914 = early_reset_static_par0_go_out;
wire _guard1915 = _guard1913 & _guard1914;
wire _guard1916 = cond_wire747_out;
wire _guard1917 = early_reset_static_par0_go_out;
wire _guard1918 = _guard1916 & _guard1917;
wire _guard1919 = cond_wire767_out;
wire _guard1920 = early_reset_static_par0_go_out;
wire _guard1921 = _guard1919 & _guard1920;
wire _guard1922 = cond_wire767_out;
wire _guard1923 = early_reset_static_par0_go_out;
wire _guard1924 = _guard1922 & _guard1923;
wire _guard1925 = cond_wire780_out;
wire _guard1926 = early_reset_static_par0_go_out;
wire _guard1927 = _guard1925 & _guard1926;
wire _guard1928 = cond_wire778_out;
wire _guard1929 = early_reset_static_par0_go_out;
wire _guard1930 = _guard1928 & _guard1929;
wire _guard1931 = fsm_out == 1'd0;
wire _guard1932 = cond_wire778_out;
wire _guard1933 = _guard1931 & _guard1932;
wire _guard1934 = fsm_out == 1'd0;
wire _guard1935 = _guard1933 & _guard1934;
wire _guard1936 = fsm_out == 1'd0;
wire _guard1937 = cond_wire780_out;
wire _guard1938 = _guard1936 & _guard1937;
wire _guard1939 = fsm_out == 1'd0;
wire _guard1940 = _guard1938 & _guard1939;
wire _guard1941 = _guard1935 | _guard1940;
wire _guard1942 = early_reset_static_par0_go_out;
wire _guard1943 = _guard1941 & _guard1942;
wire _guard1944 = fsm_out == 1'd0;
wire _guard1945 = cond_wire778_out;
wire _guard1946 = _guard1944 & _guard1945;
wire _guard1947 = fsm_out == 1'd0;
wire _guard1948 = _guard1946 & _guard1947;
wire _guard1949 = fsm_out == 1'd0;
wire _guard1950 = cond_wire780_out;
wire _guard1951 = _guard1949 & _guard1950;
wire _guard1952 = fsm_out == 1'd0;
wire _guard1953 = _guard1951 & _guard1952;
wire _guard1954 = _guard1948 | _guard1953;
wire _guard1955 = early_reset_static_par0_go_out;
wire _guard1956 = _guard1954 & _guard1955;
wire _guard1957 = fsm_out == 1'd0;
wire _guard1958 = cond_wire778_out;
wire _guard1959 = _guard1957 & _guard1958;
wire _guard1960 = fsm_out == 1'd0;
wire _guard1961 = _guard1959 & _guard1960;
wire _guard1962 = fsm_out == 1'd0;
wire _guard1963 = cond_wire780_out;
wire _guard1964 = _guard1962 & _guard1963;
wire _guard1965 = fsm_out == 1'd0;
wire _guard1966 = _guard1964 & _guard1965;
wire _guard1967 = _guard1961 | _guard1966;
wire _guard1968 = early_reset_static_par0_go_out;
wire _guard1969 = _guard1967 & _guard1968;
wire _guard1970 = cond_wire832_out;
wire _guard1971 = early_reset_static_par0_go_out;
wire _guard1972 = _guard1970 & _guard1971;
wire _guard1973 = cond_wire832_out;
wire _guard1974 = early_reset_static_par0_go_out;
wire _guard1975 = _guard1973 & _guard1974;
wire _guard1976 = cond_wire893_out;
wire _guard1977 = early_reset_static_par0_go_out;
wire _guard1978 = _guard1976 & _guard1977;
wire _guard1979 = cond_wire893_out;
wire _guard1980 = early_reset_static_par0_go_out;
wire _guard1981 = _guard1979 & _guard1980;
wire _guard1982 = cond_wire902_out;
wire _guard1983 = early_reset_static_par0_go_out;
wire _guard1984 = _guard1982 & _guard1983;
wire _guard1985 = cond_wire900_out;
wire _guard1986 = early_reset_static_par0_go_out;
wire _guard1987 = _guard1985 & _guard1986;
wire _guard1988 = fsm_out == 1'd0;
wire _guard1989 = cond_wire900_out;
wire _guard1990 = _guard1988 & _guard1989;
wire _guard1991 = fsm_out == 1'd0;
wire _guard1992 = _guard1990 & _guard1991;
wire _guard1993 = fsm_out == 1'd0;
wire _guard1994 = cond_wire902_out;
wire _guard1995 = _guard1993 & _guard1994;
wire _guard1996 = fsm_out == 1'd0;
wire _guard1997 = _guard1995 & _guard1996;
wire _guard1998 = _guard1992 | _guard1997;
wire _guard1999 = early_reset_static_par0_go_out;
wire _guard2000 = _guard1998 & _guard1999;
wire _guard2001 = fsm_out == 1'd0;
wire _guard2002 = cond_wire900_out;
wire _guard2003 = _guard2001 & _guard2002;
wire _guard2004 = fsm_out == 1'd0;
wire _guard2005 = _guard2003 & _guard2004;
wire _guard2006 = fsm_out == 1'd0;
wire _guard2007 = cond_wire902_out;
wire _guard2008 = _guard2006 & _guard2007;
wire _guard2009 = fsm_out == 1'd0;
wire _guard2010 = _guard2008 & _guard2009;
wire _guard2011 = _guard2005 | _guard2010;
wire _guard2012 = early_reset_static_par0_go_out;
wire _guard2013 = _guard2011 & _guard2012;
wire _guard2014 = fsm_out == 1'd0;
wire _guard2015 = cond_wire900_out;
wire _guard2016 = _guard2014 & _guard2015;
wire _guard2017 = fsm_out == 1'd0;
wire _guard2018 = _guard2016 & _guard2017;
wire _guard2019 = fsm_out == 1'd0;
wire _guard2020 = cond_wire902_out;
wire _guard2021 = _guard2019 & _guard2020;
wire _guard2022 = fsm_out == 1'd0;
wire _guard2023 = _guard2021 & _guard2022;
wire _guard2024 = _guard2018 | _guard2023;
wire _guard2025 = early_reset_static_par0_go_out;
wire _guard2026 = _guard2024 & _guard2025;
wire _guard2027 = cond_wire930_out;
wire _guard2028 = early_reset_static_par0_go_out;
wire _guard2029 = _guard2027 & _guard2028;
wire _guard2030 = cond_wire930_out;
wire _guard2031 = early_reset_static_par0_go_out;
wire _guard2032 = _guard2030 & _guard2031;
wire _guard2033 = fsm0_out == 6'd0;
wire _guard2034 = early_reset_static_seq_go_out;
wire _guard2035 = _guard2033 & _guard2034;
wire _guard2036 = cond_wire39_out;
wire _guard2037 = early_reset_static_par0_go_out;
wire _guard2038 = _guard2036 & _guard2037;
wire _guard2039 = _guard2035 | _guard2038;
wire _guard2040 = fsm0_out == 6'd0;
wire _guard2041 = early_reset_static_seq_go_out;
wire _guard2042 = _guard2040 & _guard2041;
wire _guard2043 = cond_wire39_out;
wire _guard2044 = early_reset_static_par0_go_out;
wire _guard2045 = _guard2043 & _guard2044;
wire _guard2046 = fsm0_out == 6'd0;
wire _guard2047 = early_reset_static_seq_go_out;
wire _guard2048 = _guard2046 & _guard2047;
wire _guard2049 = cond_wire54_out;
wire _guard2050 = early_reset_static_par0_go_out;
wire _guard2051 = _guard2049 & _guard2050;
wire _guard2052 = _guard2048 | _guard2051;
wire _guard2053 = fsm0_out == 6'd0;
wire _guard2054 = early_reset_static_seq_go_out;
wire _guard2055 = _guard2053 & _guard2054;
wire _guard2056 = cond_wire54_out;
wire _guard2057 = early_reset_static_par0_go_out;
wire _guard2058 = _guard2056 & _guard2057;
wire _guard2059 = fsm0_out == 6'd0;
wire _guard2060 = early_reset_static_seq_go_out;
wire _guard2061 = _guard2059 & _guard2060;
wire _guard2062 = cond_wire209_out;
wire _guard2063 = early_reset_static_par0_go_out;
wire _guard2064 = _guard2062 & _guard2063;
wire _guard2065 = _guard2061 | _guard2064;
wire _guard2066 = cond_wire209_out;
wire _guard2067 = early_reset_static_par0_go_out;
wire _guard2068 = _guard2066 & _guard2067;
wire _guard2069 = fsm0_out == 6'd0;
wire _guard2070 = early_reset_static_seq_go_out;
wire _guard2071 = _guard2069 & _guard2070;
wire _guard2072 = fsm0_out == 6'd0;
wire _guard2073 = early_reset_static_seq_go_out;
wire _guard2074 = _guard2072 & _guard2073;
wire _guard2075 = cond_wire469_out;
wire _guard2076 = early_reset_static_par0_go_out;
wire _guard2077 = _guard2075 & _guard2076;
wire _guard2078 = _guard2074 | _guard2077;
wire _guard2079 = fsm0_out == 6'd0;
wire _guard2080 = early_reset_static_seq_go_out;
wire _guard2081 = _guard2079 & _guard2080;
wire _guard2082 = cond_wire469_out;
wire _guard2083 = early_reset_static_par0_go_out;
wire _guard2084 = _guard2082 & _guard2083;
wire _guard2085 = fsm0_out == 6'd0;
wire _guard2086 = early_reset_static_seq_go_out;
wire _guard2087 = _guard2085 & _guard2086;
wire _guard2088 = cond_wire664_out;
wire _guard2089 = early_reset_static_par0_go_out;
wire _guard2090 = _guard2088 & _guard2089;
wire _guard2091 = _guard2087 | _guard2090;
wire _guard2092 = fsm0_out == 6'd0;
wire _guard2093 = early_reset_static_seq_go_out;
wire _guard2094 = _guard2092 & _guard2093;
wire _guard2095 = cond_wire664_out;
wire _guard2096 = early_reset_static_par0_go_out;
wire _guard2097 = _guard2095 & _guard2096;
wire _guard2098 = fsm0_out == 6'd0;
wire _guard2099 = early_reset_static_seq_go_out;
wire _guard2100 = _guard2098 & _guard2099;
wire _guard2101 = early_reset_static_par0_go_out;
wire _guard2102 = _guard2100 | _guard2101;
wire _guard2103 = early_reset_static_par0_go_out;
wire _guard2104 = fsm0_out == 6'd0;
wire _guard2105 = early_reset_static_seq_go_out;
wire _guard2106 = _guard2104 & _guard2105;
wire _guard2107 = early_reset_static_par0_go_out;
wire _guard2108 = early_reset_static_par0_go_out;
wire _guard2109 = early_reset_static_par0_go_out;
wire _guard2110 = early_reset_static_par0_go_out;
wire _guard2111 = early_reset_static_par0_go_out;
wire _guard2112 = early_reset_static_par0_go_out;
wire _guard2113 = early_reset_static_par0_go_out;
wire _guard2114 = early_reset_static_par0_go_out;
wire _guard2115 = early_reset_static_par0_go_out;
wire _guard2116 = early_reset_static_par0_go_out;
wire _guard2117 = early_reset_static_par0_go_out;
wire _guard2118 = early_reset_static_par0_go_out;
wire _guard2119 = early_reset_static_par0_go_out;
wire _guard2120 = early_reset_static_par0_go_out;
wire _guard2121 = fsm0_out == 6'd0;
wire _guard2122 = early_reset_static_seq_go_out;
wire _guard2123 = _guard2121 & _guard2122;
wire _guard2124 = early_reset_static_par0_go_out;
wire _guard2125 = _guard2123 | _guard2124;
wire _guard2126 = early_reset_static_par0_go_out;
wire _guard2127 = fsm0_out == 6'd0;
wire _guard2128 = early_reset_static_seq_go_out;
wire _guard2129 = _guard2127 & _guard2128;
wire _guard2130 = early_reset_static_par0_go_out;
wire _guard2131 = early_reset_static_par0_go_out;
wire _guard2132 = fsm0_out == 6'd0;
wire _guard2133 = early_reset_static_seq_go_out;
wire _guard2134 = _guard2132 & _guard2133;
wire _guard2135 = early_reset_static_par0_go_out;
wire _guard2136 = _guard2134 | _guard2135;
wire _guard2137 = fsm0_out == 6'd0;
wire _guard2138 = early_reset_static_seq_go_out;
wire _guard2139 = _guard2137 & _guard2138;
wire _guard2140 = early_reset_static_par0_go_out;
wire _guard2141 = fsm0_out == 6'd0;
wire _guard2142 = early_reset_static_seq_go_out;
wire _guard2143 = _guard2141 & _guard2142;
wire _guard2144 = early_reset_static_par0_go_out;
wire _guard2145 = _guard2143 | _guard2144;
wire _guard2146 = early_reset_static_par0_go_out;
wire _guard2147 = fsm0_out == 6'd0;
wire _guard2148 = early_reset_static_seq_go_out;
wire _guard2149 = _guard2147 & _guard2148;
wire _guard2150 = early_reset_static_par0_go_out;
wire _guard2151 = early_reset_static_par0_go_out;
wire _guard2152 = early_reset_static_par0_go_out;
wire _guard2153 = early_reset_static_par0_go_out;
wire _guard2154 = fsm0_out == 6'd0;
wire _guard2155 = early_reset_static_seq_go_out;
wire _guard2156 = _guard2154 & _guard2155;
wire _guard2157 = early_reset_static_par0_go_out;
wire _guard2158 = _guard2156 | _guard2157;
wire _guard2159 = early_reset_static_par0_go_out;
wire _guard2160 = fsm0_out == 6'd0;
wire _guard2161 = early_reset_static_seq_go_out;
wire _guard2162 = _guard2160 & _guard2161;
wire _guard2163 = fsm0_out == 6'd0;
wire _guard2164 = early_reset_static_seq_go_out;
wire _guard2165 = _guard2163 & _guard2164;
wire _guard2166 = early_reset_static_par0_go_out;
wire _guard2167 = _guard2165 | _guard2166;
wire _guard2168 = early_reset_static_par0_go_out;
wire _guard2169 = fsm0_out == 6'd0;
wire _guard2170 = early_reset_static_seq_go_out;
wire _guard2171 = _guard2169 & _guard2170;
wire _guard2172 = early_reset_static_par0_go_out;
wire _guard2173 = early_reset_static_par0_go_out;
wire _guard2174 = early_reset_static_par0_go_out;
wire _guard2175 = early_reset_static_par0_go_out;
wire _guard2176 = fsm0_out == 6'd0;
wire _guard2177 = early_reset_static_seq_go_out;
wire _guard2178 = _guard2176 & _guard2177;
wire _guard2179 = early_reset_static_par0_go_out;
wire _guard2180 = _guard2178 | _guard2179;
wire _guard2181 = early_reset_static_par0_go_out;
wire _guard2182 = fsm0_out == 6'd0;
wire _guard2183 = early_reset_static_seq_go_out;
wire _guard2184 = _guard2182 & _guard2183;
wire _guard2185 = early_reset_static_par0_go_out;
wire _guard2186 = early_reset_static_par0_go_out;
wire _guard2187 = early_reset_static_par0_go_out;
wire _guard2188 = early_reset_static_par0_go_out;
wire _guard2189 = early_reset_static_par0_go_out;
wire _guard2190 = early_reset_static_par0_go_out;
wire _guard2191 = fsm0_out == 6'd0;
wire _guard2192 = early_reset_static_seq_go_out;
wire _guard2193 = _guard2191 & _guard2192;
wire _guard2194 = early_reset_static_par0_go_out;
wire _guard2195 = _guard2193 | _guard2194;
wire _guard2196 = fsm0_out == 6'd0;
wire _guard2197 = early_reset_static_seq_go_out;
wire _guard2198 = _guard2196 & _guard2197;
wire _guard2199 = early_reset_static_par0_go_out;
wire _guard2200 = wrapper_early_reset_static_seq_done_out;
wire _guard2201 = cond_wire9_out;
wire _guard2202 = early_reset_static_par0_go_out;
wire _guard2203 = _guard2201 & _guard2202;
wire _guard2204 = cond_wire64_out;
wire _guard2205 = early_reset_static_par0_go_out;
wire _guard2206 = _guard2204 & _guard2205;
wire _guard2207 = cond_wire989_out;
wire _guard2208 = early_reset_static_par0_go_out;
wire _guard2209 = _guard2207 & _guard2208;
wire _guard2210 = cond_wire314_out;
wire _guard2211 = early_reset_static_par0_go_out;
wire _guard2212 = _guard2210 & _guard2211;
wire _guard2213 = cond_wire278_out;
wire _guard2214 = early_reset_static_par0_go_out;
wire _guard2215 = _guard2213 & _guard2214;
wire _guard2216 = cond_wire298_out;
wire _guard2217 = early_reset_static_par0_go_out;
wire _guard2218 = _guard2216 & _guard2217;
wire _guard2219 = cond_wire326_out;
wire _guard2220 = early_reset_static_par0_go_out;
wire _guard2221 = _guard2219 & _guard2220;
wire _guard2222 = cond_wire334_out;
wire _guard2223 = early_reset_static_par0_go_out;
wire _guard2224 = _guard2222 & _guard2223;
wire _guard2225 = cond_wire338_out;
wire _guard2226 = early_reset_static_par0_go_out;
wire _guard2227 = _guard2225 & _guard2226;
wire _guard2228 = cond_wire302_out;
wire _guard2229 = early_reset_static_par0_go_out;
wire _guard2230 = _guard2228 & _guard2229;
wire _guard2231 = cond_wire322_out;
wire _guard2232 = early_reset_static_par0_go_out;
wire _guard2233 = _guard2231 & _guard2232;
wire _guard2234 = cond_wire286_out;
wire _guard2235 = early_reset_static_par0_go_out;
wire _guard2236 = _guard2234 & _guard2235;
wire _guard2237 = cond_wire310_out;
wire _guard2238 = early_reset_static_par0_go_out;
wire _guard2239 = _guard2237 & _guard2238;
wire _guard2240 = cond_wire294_out;
wire _guard2241 = early_reset_static_par0_go_out;
wire _guard2242 = _guard2240 & _guard2241;
wire _guard2243 = cond_wire306_out;
wire _guard2244 = early_reset_static_par0_go_out;
wire _guard2245 = _guard2243 & _guard2244;
wire _guard2246 = cond_wire330_out;
wire _guard2247 = early_reset_static_par0_go_out;
wire _guard2248 = _guard2246 & _guard2247;
wire _guard2249 = cond_wire290_out;
wire _guard2250 = early_reset_static_par0_go_out;
wire _guard2251 = _guard2249 & _guard2250;
wire _guard2252 = cond_wire318_out;
wire _guard2253 = early_reset_static_par0_go_out;
wire _guard2254 = _guard2252 & _guard2253;
wire _guard2255 = cond_wire282_out;
wire _guard2256 = early_reset_static_par0_go_out;
wire _guard2257 = _guard2255 & _guard2256;
wire _guard2258 = cond_wire802_out;
wire _guard2259 = early_reset_static_par0_go_out;
wire _guard2260 = _guard2258 & _guard2259;
wire _guard2261 = cond_wire858_out;
wire _guard2262 = early_reset_static_par0_go_out;
wire _guard2263 = _guard2261 & _guard2262;
wire _guard2264 = cond_wire798_out;
wire _guard2265 = early_reset_static_par0_go_out;
wire _guard2266 = _guard2264 & _guard2265;
wire _guard2267 = cond_wire810_out;
wire _guard2268 = early_reset_static_par0_go_out;
wire _guard2269 = _guard2267 & _guard2268;
wire _guard2270 = cond_wire850_out;
wire _guard2271 = early_reset_static_par0_go_out;
wire _guard2272 = _guard2270 & _guard2271;
wire _guard2273 = cond_wire854_out;
wire _guard2274 = early_reset_static_par0_go_out;
wire _guard2275 = _guard2273 & _guard2274;
wire _guard2276 = cond_wire818_out;
wire _guard2277 = early_reset_static_par0_go_out;
wire _guard2278 = _guard2276 & _guard2277;
wire _guard2279 = cond_wire846_out;
wire _guard2280 = early_reset_static_par0_go_out;
wire _guard2281 = _guard2279 & _guard2280;
wire _guard2282 = cond_wire806_out;
wire _guard2283 = early_reset_static_par0_go_out;
wire _guard2284 = _guard2282 & _guard2283;
wire _guard2285 = cond_wire830_out;
wire _guard2286 = early_reset_static_par0_go_out;
wire _guard2287 = _guard2285 & _guard2286;
wire _guard2288 = cond_wire838_out;
wire _guard2289 = early_reset_static_par0_go_out;
wire _guard2290 = _guard2288 & _guard2289;
wire _guard2291 = cond_wire826_out;
wire _guard2292 = early_reset_static_par0_go_out;
wire _guard2293 = _guard2291 & _guard2292;
wire _guard2294 = cond_wire842_out;
wire _guard2295 = early_reset_static_par0_go_out;
wire _guard2296 = _guard2294 & _guard2295;
wire _guard2297 = cond_wire814_out;
wire _guard2298 = early_reset_static_par0_go_out;
wire _guard2299 = _guard2297 & _guard2298;
wire _guard2300 = cond_wire822_out;
wire _guard2301 = early_reset_static_par0_go_out;
wire _guard2302 = _guard2300 & _guard2301;
wire _guard2303 = cond_wire834_out;
wire _guard2304 = early_reset_static_par0_go_out;
wire _guard2305 = _guard2303 & _guard2304;
wire _guard2306 = cond_wire339_out;
wire _guard2307 = early_reset_static_par0_go_out;
wire _guard2308 = _guard2306 & _guard2307;
wire _guard2309 = cond_wire997_out;
wire _guard2310 = early_reset_static_par0_go_out;
wire _guard2311 = _guard2309 & _guard2310;
wire _guard2312 = cond_wire1052_out;
wire _guard2313 = early_reset_static_par0_go_out;
wire _guard2314 = _guard2312 & _guard2313;
wire _guard2315 = cond_wire993_out;
wire _guard2316 = early_reset_static_par0_go_out;
wire _guard2317 = _guard2315 & _guard2316;
wire _guard2318 = cond_wire1005_out;
wire _guard2319 = early_reset_static_par0_go_out;
wire _guard2320 = _guard2318 & _guard2319;
wire _guard2321 = cond_wire1045_out;
wire _guard2322 = early_reset_static_par0_go_out;
wire _guard2323 = _guard2321 & _guard2322;
wire _guard2324 = cond_wire1049_out;
wire _guard2325 = early_reset_static_par0_go_out;
wire _guard2326 = _guard2324 & _guard2325;
wire _guard2327 = cond_wire1013_out;
wire _guard2328 = early_reset_static_par0_go_out;
wire _guard2329 = _guard2327 & _guard2328;
wire _guard2330 = cond_wire1041_out;
wire _guard2331 = early_reset_static_par0_go_out;
wire _guard2332 = _guard2330 & _guard2331;
wire _guard2333 = cond_wire1001_out;
wire _guard2334 = early_reset_static_par0_go_out;
wire _guard2335 = _guard2333 & _guard2334;
wire _guard2336 = cond_wire1025_out;
wire _guard2337 = early_reset_static_par0_go_out;
wire _guard2338 = _guard2336 & _guard2337;
wire _guard2339 = cond_wire1033_out;
wire _guard2340 = early_reset_static_par0_go_out;
wire _guard2341 = _guard2339 & _guard2340;
wire _guard2342 = cond_wire1021_out;
wire _guard2343 = early_reset_static_par0_go_out;
wire _guard2344 = _guard2342 & _guard2343;
wire _guard2345 = cond_wire1037_out;
wire _guard2346 = early_reset_static_par0_go_out;
wire _guard2347 = _guard2345 & _guard2346;
wire _guard2348 = cond_wire1009_out;
wire _guard2349 = early_reset_static_par0_go_out;
wire _guard2350 = _guard2348 & _guard2349;
wire _guard2351 = cond_wire1017_out;
wire _guard2352 = early_reset_static_par0_go_out;
wire _guard2353 = _guard2351 & _guard2352;
wire _guard2354 = cond_wire1029_out;
wire _guard2355 = early_reset_static_par0_go_out;
wire _guard2356 = _guard2354 & _guard2355;
wire _guard2357 = cond_wire_out;
wire _guard2358 = early_reset_static_par0_go_out;
wire _guard2359 = _guard2357 & _guard2358;
wire _guard2360 = cond_wire87_out;
wire _guard2361 = early_reset_static_par0_go_out;
wire _guard2362 = _guard2360 & _guard2361;
wire _guard2363 = cond_wire143_out;
wire _guard2364 = early_reset_static_par0_go_out;
wire _guard2365 = _guard2363 & _guard2364;
wire _guard2366 = cond_wire83_out;
wire _guard2367 = early_reset_static_par0_go_out;
wire _guard2368 = _guard2366 & _guard2367;
wire _guard2369 = cond_wire95_out;
wire _guard2370 = early_reset_static_par0_go_out;
wire _guard2371 = _guard2369 & _guard2370;
wire _guard2372 = cond_wire135_out;
wire _guard2373 = early_reset_static_par0_go_out;
wire _guard2374 = _guard2372 & _guard2373;
wire _guard2375 = cond_wire139_out;
wire _guard2376 = early_reset_static_par0_go_out;
wire _guard2377 = _guard2375 & _guard2376;
wire _guard2378 = cond_wire103_out;
wire _guard2379 = early_reset_static_par0_go_out;
wire _guard2380 = _guard2378 & _guard2379;
wire _guard2381 = cond_wire131_out;
wire _guard2382 = early_reset_static_par0_go_out;
wire _guard2383 = _guard2381 & _guard2382;
wire _guard2384 = cond_wire91_out;
wire _guard2385 = early_reset_static_par0_go_out;
wire _guard2386 = _guard2384 & _guard2385;
wire _guard2387 = cond_wire115_out;
wire _guard2388 = early_reset_static_par0_go_out;
wire _guard2389 = _guard2387 & _guard2388;
wire _guard2390 = cond_wire123_out;
wire _guard2391 = early_reset_static_par0_go_out;
wire _guard2392 = _guard2390 & _guard2391;
wire _guard2393 = cond_wire111_out;
wire _guard2394 = early_reset_static_par0_go_out;
wire _guard2395 = _guard2393 & _guard2394;
wire _guard2396 = cond_wire127_out;
wire _guard2397 = early_reset_static_par0_go_out;
wire _guard2398 = _guard2396 & _guard2397;
wire _guard2399 = cond_wire99_out;
wire _guard2400 = early_reset_static_par0_go_out;
wire _guard2401 = _guard2399 & _guard2400;
wire _guard2402 = cond_wire107_out;
wire _guard2403 = early_reset_static_par0_go_out;
wire _guard2404 = _guard2402 & _guard2403;
wire _guard2405 = cond_wire119_out;
wire _guard2406 = early_reset_static_par0_go_out;
wire _guard2407 = _guard2405 & _guard2406;
wire _guard2408 = cond_wire347_out;
wire _guard2409 = early_reset_static_par0_go_out;
wire _guard2410 = _guard2408 & _guard2409;
wire _guard2411 = cond_wire403_out;
wire _guard2412 = early_reset_static_par0_go_out;
wire _guard2413 = _guard2411 & _guard2412;
wire _guard2414 = cond_wire343_out;
wire _guard2415 = early_reset_static_par0_go_out;
wire _guard2416 = _guard2414 & _guard2415;
wire _guard2417 = cond_wire355_out;
wire _guard2418 = early_reset_static_par0_go_out;
wire _guard2419 = _guard2417 & _guard2418;
wire _guard2420 = cond_wire395_out;
wire _guard2421 = early_reset_static_par0_go_out;
wire _guard2422 = _guard2420 & _guard2421;
wire _guard2423 = cond_wire399_out;
wire _guard2424 = early_reset_static_par0_go_out;
wire _guard2425 = _guard2423 & _guard2424;
wire _guard2426 = cond_wire363_out;
wire _guard2427 = early_reset_static_par0_go_out;
wire _guard2428 = _guard2426 & _guard2427;
wire _guard2429 = cond_wire391_out;
wire _guard2430 = early_reset_static_par0_go_out;
wire _guard2431 = _guard2429 & _guard2430;
wire _guard2432 = cond_wire351_out;
wire _guard2433 = early_reset_static_par0_go_out;
wire _guard2434 = _guard2432 & _guard2433;
wire _guard2435 = cond_wire375_out;
wire _guard2436 = early_reset_static_par0_go_out;
wire _guard2437 = _guard2435 & _guard2436;
wire _guard2438 = cond_wire383_out;
wire _guard2439 = early_reset_static_par0_go_out;
wire _guard2440 = _guard2438 & _guard2439;
wire _guard2441 = cond_wire371_out;
wire _guard2442 = early_reset_static_par0_go_out;
wire _guard2443 = _guard2441 & _guard2442;
wire _guard2444 = cond_wire387_out;
wire _guard2445 = early_reset_static_par0_go_out;
wire _guard2446 = _guard2444 & _guard2445;
wire _guard2447 = cond_wire359_out;
wire _guard2448 = early_reset_static_par0_go_out;
wire _guard2449 = _guard2447 & _guard2448;
wire _guard2450 = cond_wire367_out;
wire _guard2451 = early_reset_static_par0_go_out;
wire _guard2452 = _guard2450 & _guard2451;
wire _guard2453 = cond_wire379_out;
wire _guard2454 = early_reset_static_par0_go_out;
wire _guard2455 = _guard2453 & _guard2454;
wire _guard2456 = cond_wire351_out;
wire _guard2457 = early_reset_static_par0_go_out;
wire _guard2458 = _guard2456 & _guard2457;
wire _guard2459 = cond_wire375_out;
wire _guard2460 = early_reset_static_par0_go_out;
wire _guard2461 = _guard2459 & _guard2460;
wire _guard2462 = cond_wire395_out;
wire _guard2463 = early_reset_static_par0_go_out;
wire _guard2464 = _guard2462 & _guard2463;
wire _guard2465 = cond_wire343_out;
wire _guard2466 = early_reset_static_par0_go_out;
wire _guard2467 = _guard2465 & _guard2466;
wire _guard2468 = cond_wire359_out;
wire _guard2469 = early_reset_static_par0_go_out;
wire _guard2470 = _guard2468 & _guard2469;
wire _guard2471 = cond_wire347_out;
wire _guard2472 = early_reset_static_par0_go_out;
wire _guard2473 = _guard2471 & _guard2472;
wire _guard2474 = cond_wire371_out;
wire _guard2475 = early_reset_static_par0_go_out;
wire _guard2476 = _guard2474 & _guard2475;
wire _guard2477 = cond_wire379_out;
wire _guard2478 = early_reset_static_par0_go_out;
wire _guard2479 = _guard2477 & _guard2478;
wire _guard2480 = cond_wire383_out;
wire _guard2481 = early_reset_static_par0_go_out;
wire _guard2482 = _guard2480 & _guard2481;
wire _guard2483 = cond_wire355_out;
wire _guard2484 = early_reset_static_par0_go_out;
wire _guard2485 = _guard2483 & _guard2484;
wire _guard2486 = cond_wire363_out;
wire _guard2487 = early_reset_static_par0_go_out;
wire _guard2488 = _guard2486 & _guard2487;
wire _guard2489 = cond_wire399_out;
wire _guard2490 = early_reset_static_par0_go_out;
wire _guard2491 = _guard2489 & _guard2490;
wire _guard2492 = cond_wire367_out;
wire _guard2493 = early_reset_static_par0_go_out;
wire _guard2494 = _guard2492 & _guard2493;
wire _guard2495 = cond_wire387_out;
wire _guard2496 = early_reset_static_par0_go_out;
wire _guard2497 = _guard2495 & _guard2496;
wire _guard2498 = cond_wire403_out;
wire _guard2499 = early_reset_static_par0_go_out;
wire _guard2500 = _guard2498 & _guard2499;
wire _guard2501 = cond_wire391_out;
wire _guard2502 = early_reset_static_par0_go_out;
wire _guard2503 = _guard2501 & _guard2502;
wire _guard2504 = cond_wire737_out;
wire _guard2505 = early_reset_static_par0_go_out;
wire _guard2506 = _guard2504 & _guard2505;
wire _guard2507 = cond_wire793_out;
wire _guard2508 = early_reset_static_par0_go_out;
wire _guard2509 = _guard2507 & _guard2508;
wire _guard2510 = cond_wire733_out;
wire _guard2511 = early_reset_static_par0_go_out;
wire _guard2512 = _guard2510 & _guard2511;
wire _guard2513 = cond_wire745_out;
wire _guard2514 = early_reset_static_par0_go_out;
wire _guard2515 = _guard2513 & _guard2514;
wire _guard2516 = cond_wire785_out;
wire _guard2517 = early_reset_static_par0_go_out;
wire _guard2518 = _guard2516 & _guard2517;
wire _guard2519 = cond_wire789_out;
wire _guard2520 = early_reset_static_par0_go_out;
wire _guard2521 = _guard2519 & _guard2520;
wire _guard2522 = cond_wire753_out;
wire _guard2523 = early_reset_static_par0_go_out;
wire _guard2524 = _guard2522 & _guard2523;
wire _guard2525 = cond_wire781_out;
wire _guard2526 = early_reset_static_par0_go_out;
wire _guard2527 = _guard2525 & _guard2526;
wire _guard2528 = cond_wire741_out;
wire _guard2529 = early_reset_static_par0_go_out;
wire _guard2530 = _guard2528 & _guard2529;
wire _guard2531 = cond_wire765_out;
wire _guard2532 = early_reset_static_par0_go_out;
wire _guard2533 = _guard2531 & _guard2532;
wire _guard2534 = cond_wire773_out;
wire _guard2535 = early_reset_static_par0_go_out;
wire _guard2536 = _guard2534 & _guard2535;
wire _guard2537 = cond_wire761_out;
wire _guard2538 = early_reset_static_par0_go_out;
wire _guard2539 = _guard2537 & _guard2538;
wire _guard2540 = cond_wire777_out;
wire _guard2541 = early_reset_static_par0_go_out;
wire _guard2542 = _guard2540 & _guard2541;
wire _guard2543 = cond_wire749_out;
wire _guard2544 = early_reset_static_par0_go_out;
wire _guard2545 = _guard2543 & _guard2544;
wire _guard2546 = cond_wire757_out;
wire _guard2547 = early_reset_static_par0_go_out;
wire _guard2548 = _guard2546 & _guard2547;
wire _guard2549 = cond_wire769_out;
wire _guard2550 = early_reset_static_par0_go_out;
wire _guard2551 = _guard2549 & _guard2550;
wire _guard2552 = cond_wire404_out;
wire _guard2553 = early_reset_static_par0_go_out;
wire _guard2554 = _guard2552 & _guard2553;
wire _guard2555 = cond_wire53_out;
wire _guard2556 = early_reset_static_par0_go_out;
wire _guard2557 = _guard2555 & _guard2556;
wire _guard2558 = cond_wire8_out;
wire _guard2559 = early_reset_static_par0_go_out;
wire _guard2560 = _guard2558 & _guard2559;
wire _guard2561 = cond_wire38_out;
wire _guard2562 = early_reset_static_par0_go_out;
wire _guard2563 = _guard2561 & _guard2562;
wire _guard2564 = cond_wire18_out;
wire _guard2565 = early_reset_static_par0_go_out;
wire _guard2566 = _guard2564 & _guard2565;
wire _guard2567 = cond_wire28_out;
wire _guard2568 = early_reset_static_par0_go_out;
wire _guard2569 = _guard2567 & _guard2568;
wire _guard2570 = cond_wire43_out;
wire _guard2571 = early_reset_static_par0_go_out;
wire _guard2572 = _guard2570 & _guard2571;
wire _guard2573 = cond_wire48_out;
wire _guard2574 = early_reset_static_par0_go_out;
wire _guard2575 = _guard2573 & _guard2574;
wire _guard2576 = cond_wire13_out;
wire _guard2577 = early_reset_static_par0_go_out;
wire _guard2578 = _guard2576 & _guard2577;
wire _guard2579 = cond_wire63_out;
wire _guard2580 = early_reset_static_par0_go_out;
wire _guard2581 = _guard2579 & _guard2580;
wire _guard2582 = cond_wire78_out;
wire _guard2583 = early_reset_static_par0_go_out;
wire _guard2584 = _guard2582 & _guard2583;
wire _guard2585 = cond_wire23_out;
wire _guard2586 = early_reset_static_par0_go_out;
wire _guard2587 = _guard2585 & _guard2586;
wire _guard2588 = cond_wire73_out;
wire _guard2589 = early_reset_static_par0_go_out;
wire _guard2590 = _guard2588 & _guard2589;
wire _guard2591 = cond_wire58_out;
wire _guard2592 = early_reset_static_par0_go_out;
wire _guard2593 = _guard2591 & _guard2592;
wire _guard2594 = cond_wire3_out;
wire _guard2595 = early_reset_static_par0_go_out;
wire _guard2596 = _guard2594 & _guard2595;
wire _guard2597 = cond_wire33_out;
wire _guard2598 = early_reset_static_par0_go_out;
wire _guard2599 = _guard2597 & _guard2598;
wire _guard2600 = cond_wire68_out;
wire _guard2601 = early_reset_static_par0_go_out;
wire _guard2602 = _guard2600 & _guard2601;
wire _guard2603 = cond_wire838_out;
wire _guard2604 = early_reset_static_par0_go_out;
wire _guard2605 = _guard2603 & _guard2604;
wire _guard2606 = cond_wire834_out;
wire _guard2607 = early_reset_static_par0_go_out;
wire _guard2608 = _guard2606 & _guard2607;
wire _guard2609 = cond_wire846_out;
wire _guard2610 = early_reset_static_par0_go_out;
wire _guard2611 = _guard2609 & _guard2610;
wire _guard2612 = cond_wire810_out;
wire _guard2613 = early_reset_static_par0_go_out;
wire _guard2614 = _guard2612 & _guard2613;
wire _guard2615 = cond_wire814_out;
wire _guard2616 = early_reset_static_par0_go_out;
wire _guard2617 = _guard2615 & _guard2616;
wire _guard2618 = cond_wire802_out;
wire _guard2619 = early_reset_static_par0_go_out;
wire _guard2620 = _guard2618 & _guard2619;
wire _guard2621 = cond_wire826_out;
wire _guard2622 = early_reset_static_par0_go_out;
wire _guard2623 = _guard2621 & _guard2622;
wire _guard2624 = cond_wire842_out;
wire _guard2625 = early_reset_static_par0_go_out;
wire _guard2626 = _guard2624 & _guard2625;
wire _guard2627 = cond_wire822_out;
wire _guard2628 = early_reset_static_par0_go_out;
wire _guard2629 = _guard2627 & _guard2628;
wire _guard2630 = cond_wire818_out;
wire _guard2631 = early_reset_static_par0_go_out;
wire _guard2632 = _guard2630 & _guard2631;
wire _guard2633 = cond_wire850_out;
wire _guard2634 = early_reset_static_par0_go_out;
wire _guard2635 = _guard2633 & _guard2634;
wire _guard2636 = cond_wire858_out;
wire _guard2637 = early_reset_static_par0_go_out;
wire _guard2638 = _guard2636 & _guard2637;
wire _guard2639 = cond_wire798_out;
wire _guard2640 = early_reset_static_par0_go_out;
wire _guard2641 = _guard2639 & _guard2640;
wire _guard2642 = cond_wire806_out;
wire _guard2643 = early_reset_static_par0_go_out;
wire _guard2644 = _guard2642 & _guard2643;
wire _guard2645 = cond_wire830_out;
wire _guard2646 = early_reset_static_par0_go_out;
wire _guard2647 = _guard2645 & _guard2646;
wire _guard2648 = cond_wire854_out;
wire _guard2649 = early_reset_static_par0_go_out;
wire _guard2650 = _guard2648 & _guard2649;
wire _guard2651 = cond_wire859_out;
wire _guard2652 = early_reset_static_par0_go_out;
wire _guard2653 = _guard2651 & _guard2652;
wire _guard2654 = cond_wire412_out;
wire _guard2655 = early_reset_static_par0_go_out;
wire _guard2656 = _guard2654 & _guard2655;
wire _guard2657 = cond_wire468_out;
wire _guard2658 = early_reset_static_par0_go_out;
wire _guard2659 = _guard2657 & _guard2658;
wire _guard2660 = cond_wire408_out;
wire _guard2661 = early_reset_static_par0_go_out;
wire _guard2662 = _guard2660 & _guard2661;
wire _guard2663 = cond_wire420_out;
wire _guard2664 = early_reset_static_par0_go_out;
wire _guard2665 = _guard2663 & _guard2664;
wire _guard2666 = cond_wire460_out;
wire _guard2667 = early_reset_static_par0_go_out;
wire _guard2668 = _guard2666 & _guard2667;
wire _guard2669 = cond_wire464_out;
wire _guard2670 = early_reset_static_par0_go_out;
wire _guard2671 = _guard2669 & _guard2670;
wire _guard2672 = cond_wire428_out;
wire _guard2673 = early_reset_static_par0_go_out;
wire _guard2674 = _guard2672 & _guard2673;
wire _guard2675 = cond_wire456_out;
wire _guard2676 = early_reset_static_par0_go_out;
wire _guard2677 = _guard2675 & _guard2676;
wire _guard2678 = cond_wire416_out;
wire _guard2679 = early_reset_static_par0_go_out;
wire _guard2680 = _guard2678 & _guard2679;
wire _guard2681 = cond_wire440_out;
wire _guard2682 = early_reset_static_par0_go_out;
wire _guard2683 = _guard2681 & _guard2682;
wire _guard2684 = cond_wire448_out;
wire _guard2685 = early_reset_static_par0_go_out;
wire _guard2686 = _guard2684 & _guard2685;
wire _guard2687 = cond_wire436_out;
wire _guard2688 = early_reset_static_par0_go_out;
wire _guard2689 = _guard2687 & _guard2688;
wire _guard2690 = cond_wire452_out;
wire _guard2691 = early_reset_static_par0_go_out;
wire _guard2692 = _guard2690 & _guard2691;
wire _guard2693 = cond_wire424_out;
wire _guard2694 = early_reset_static_par0_go_out;
wire _guard2695 = _guard2693 & _guard2694;
wire _guard2696 = cond_wire432_out;
wire _guard2697 = early_reset_static_par0_go_out;
wire _guard2698 = _guard2696 & _guard2697;
wire _guard2699 = cond_wire444_out;
wire _guard2700 = early_reset_static_par0_go_out;
wire _guard2701 = _guard2699 & _guard2700;
wire _guard2702 = cond_wire729_out;
wire _guard2703 = early_reset_static_par0_go_out;
wire _guard2704 = _guard2702 & _guard2703;
wire _guard2705 = cond_wire924_out;
wire _guard2706 = early_reset_static_par0_go_out;
wire _guard2707 = _guard2705 & _guard2706;
wire _guard2708 = cond_wire245_out;
wire _guard2709 = early_reset_static_par0_go_out;
wire _guard2710 = _guard2708 & _guard2709;
wire _guard2711 = cond_wire229_out;
wire _guard2712 = early_reset_static_par0_go_out;
wire _guard2713 = _guard2711 & _guard2712;
wire _guard2714 = cond_wire241_out;
wire _guard2715 = early_reset_static_par0_go_out;
wire _guard2716 = _guard2714 & _guard2715;
wire _guard2717 = cond_wire273_out;
wire _guard2718 = early_reset_static_par0_go_out;
wire _guard2719 = _guard2717 & _guard2718;
wire _guard2720 = cond_wire221_out;
wire _guard2721 = early_reset_static_par0_go_out;
wire _guard2722 = _guard2720 & _guard2721;
wire _guard2723 = cond_wire233_out;
wire _guard2724 = early_reset_static_par0_go_out;
wire _guard2725 = _guard2723 & _guard2724;
wire _guard2726 = cond_wire237_out;
wire _guard2727 = early_reset_static_par0_go_out;
wire _guard2728 = _guard2726 & _guard2727;
wire _guard2729 = cond_wire213_out;
wire _guard2730 = early_reset_static_par0_go_out;
wire _guard2731 = _guard2729 & _guard2730;
wire _guard2732 = cond_wire265_out;
wire _guard2733 = early_reset_static_par0_go_out;
wire _guard2734 = _guard2732 & _guard2733;
wire _guard2735 = cond_wire269_out;
wire _guard2736 = early_reset_static_par0_go_out;
wire _guard2737 = _guard2735 & _guard2736;
wire _guard2738 = cond_wire217_out;
wire _guard2739 = early_reset_static_par0_go_out;
wire _guard2740 = _guard2738 & _guard2739;
wire _guard2741 = cond_wire253_out;
wire _guard2742 = early_reset_static_par0_go_out;
wire _guard2743 = _guard2741 & _guard2742;
wire _guard2744 = cond_wire249_out;
wire _guard2745 = early_reset_static_par0_go_out;
wire _guard2746 = _guard2744 & _guard2745;
wire _guard2747 = cond_wire257_out;
wire _guard2748 = early_reset_static_par0_go_out;
wire _guard2749 = _guard2747 & _guard2748;
wire _guard2750 = cond_wire261_out;
wire _guard2751 = early_reset_static_par0_go_out;
wire _guard2752 = _guard2750 & _guard2751;
wire _guard2753 = cond_wire225_out;
wire _guard2754 = early_reset_static_par0_go_out;
wire _guard2755 = _guard2753 & _guard2754;
wire _guard2756 = fsm_out == 1'd0;
wire _guard2757 = cond_wire603_out;
wire _guard2758 = _guard2756 & _guard2757;
wire _guard2759 = fsm_out == 1'd0;
wire _guard2760 = _guard2758 & _guard2759;
wire _guard2761 = fsm_out == 1'd0;
wire _guard2762 = cond_wire607_out;
wire _guard2763 = _guard2761 & _guard2762;
wire _guard2764 = fsm_out == 1'd0;
wire _guard2765 = _guard2763 & _guard2764;
wire _guard2766 = _guard2760 | _guard2765;
wire _guard2767 = fsm_out == 1'd0;
wire _guard2768 = cond_wire611_out;
wire _guard2769 = _guard2767 & _guard2768;
wire _guard2770 = fsm_out == 1'd0;
wire _guard2771 = _guard2769 & _guard2770;
wire _guard2772 = _guard2766 | _guard2771;
wire _guard2773 = fsm_out == 1'd0;
wire _guard2774 = cond_wire615_out;
wire _guard2775 = _guard2773 & _guard2774;
wire _guard2776 = fsm_out == 1'd0;
wire _guard2777 = _guard2775 & _guard2776;
wire _guard2778 = _guard2772 | _guard2777;
wire _guard2779 = fsm_out == 1'd0;
wire _guard2780 = cond_wire619_out;
wire _guard2781 = _guard2779 & _guard2780;
wire _guard2782 = fsm_out == 1'd0;
wire _guard2783 = _guard2781 & _guard2782;
wire _guard2784 = _guard2778 | _guard2783;
wire _guard2785 = fsm_out == 1'd0;
wire _guard2786 = cond_wire623_out;
wire _guard2787 = _guard2785 & _guard2786;
wire _guard2788 = fsm_out == 1'd0;
wire _guard2789 = _guard2787 & _guard2788;
wire _guard2790 = _guard2784 | _guard2789;
wire _guard2791 = fsm_out == 1'd0;
wire _guard2792 = cond_wire627_out;
wire _guard2793 = _guard2791 & _guard2792;
wire _guard2794 = fsm_out == 1'd0;
wire _guard2795 = _guard2793 & _guard2794;
wire _guard2796 = _guard2790 | _guard2795;
wire _guard2797 = fsm_out == 1'd0;
wire _guard2798 = cond_wire631_out;
wire _guard2799 = _guard2797 & _guard2798;
wire _guard2800 = fsm_out == 1'd0;
wire _guard2801 = _guard2799 & _guard2800;
wire _guard2802 = _guard2796 | _guard2801;
wire _guard2803 = fsm_out == 1'd0;
wire _guard2804 = cond_wire635_out;
wire _guard2805 = _guard2803 & _guard2804;
wire _guard2806 = fsm_out == 1'd0;
wire _guard2807 = _guard2805 & _guard2806;
wire _guard2808 = _guard2802 | _guard2807;
wire _guard2809 = fsm_out == 1'd0;
wire _guard2810 = cond_wire639_out;
wire _guard2811 = _guard2809 & _guard2810;
wire _guard2812 = fsm_out == 1'd0;
wire _guard2813 = _guard2811 & _guard2812;
wire _guard2814 = _guard2808 | _guard2813;
wire _guard2815 = fsm_out == 1'd0;
wire _guard2816 = cond_wire643_out;
wire _guard2817 = _guard2815 & _guard2816;
wire _guard2818 = fsm_out == 1'd0;
wire _guard2819 = _guard2817 & _guard2818;
wire _guard2820 = _guard2814 | _guard2819;
wire _guard2821 = fsm_out == 1'd0;
wire _guard2822 = cond_wire647_out;
wire _guard2823 = _guard2821 & _guard2822;
wire _guard2824 = fsm_out == 1'd0;
wire _guard2825 = _guard2823 & _guard2824;
wire _guard2826 = _guard2820 | _guard2825;
wire _guard2827 = fsm_out == 1'd0;
wire _guard2828 = cond_wire651_out;
wire _guard2829 = _guard2827 & _guard2828;
wire _guard2830 = fsm_out == 1'd0;
wire _guard2831 = _guard2829 & _guard2830;
wire _guard2832 = _guard2826 | _guard2831;
wire _guard2833 = fsm_out == 1'd0;
wire _guard2834 = cond_wire655_out;
wire _guard2835 = _guard2833 & _guard2834;
wire _guard2836 = fsm_out == 1'd0;
wire _guard2837 = _guard2835 & _guard2836;
wire _guard2838 = _guard2832 | _guard2837;
wire _guard2839 = fsm_out == 1'd0;
wire _guard2840 = cond_wire659_out;
wire _guard2841 = _guard2839 & _guard2840;
wire _guard2842 = fsm_out == 1'd0;
wire _guard2843 = _guard2841 & _guard2842;
wire _guard2844 = _guard2838 | _guard2843;
wire _guard2845 = fsm_out == 1'd0;
wire _guard2846 = cond_wire663_out;
wire _guard2847 = _guard2845 & _guard2846;
wire _guard2848 = fsm_out == 1'd0;
wire _guard2849 = _guard2847 & _guard2848;
wire _guard2850 = _guard2844 | _guard2849;
wire _guard2851 = early_reset_static_par0_go_out;
wire _guard2852 = _guard2850 & _guard2851;
wire _guard2853 = cond_wire688_out;
wire _guard2854 = early_reset_static_par0_go_out;
wire _guard2855 = _guard2853 & _guard2854;
wire _guard2856 = cond_wire696_out;
wire _guard2857 = early_reset_static_par0_go_out;
wire _guard2858 = _guard2856 & _guard2857;
wire _guard2859 = cond_wire704_out;
wire _guard2860 = early_reset_static_par0_go_out;
wire _guard2861 = _guard2859 & _guard2860;
wire _guard2862 = cond_wire700_out;
wire _guard2863 = early_reset_static_par0_go_out;
wire _guard2864 = _guard2862 & _guard2863;
wire _guard2865 = cond_wire720_out;
wire _guard2866 = early_reset_static_par0_go_out;
wire _guard2867 = _guard2865 & _guard2866;
wire _guard2868 = cond_wire716_out;
wire _guard2869 = early_reset_static_par0_go_out;
wire _guard2870 = _guard2868 & _guard2869;
wire _guard2871 = cond_wire668_out;
wire _guard2872 = early_reset_static_par0_go_out;
wire _guard2873 = _guard2871 & _guard2872;
wire _guard2874 = cond_wire724_out;
wire _guard2875 = early_reset_static_par0_go_out;
wire _guard2876 = _guard2874 & _guard2875;
wire _guard2877 = cond_wire708_out;
wire _guard2878 = early_reset_static_par0_go_out;
wire _guard2879 = _guard2877 & _guard2878;
wire _guard2880 = cond_wire676_out;
wire _guard2881 = early_reset_static_par0_go_out;
wire _guard2882 = _guard2880 & _guard2881;
wire _guard2883 = cond_wire680_out;
wire _guard2884 = early_reset_static_par0_go_out;
wire _guard2885 = _guard2883 & _guard2884;
wire _guard2886 = cond_wire684_out;
wire _guard2887 = early_reset_static_par0_go_out;
wire _guard2888 = _guard2886 & _guard2887;
wire _guard2889 = cond_wire728_out;
wire _guard2890 = early_reset_static_par0_go_out;
wire _guard2891 = _guard2889 & _guard2890;
wire _guard2892 = cond_wire712_out;
wire _guard2893 = early_reset_static_par0_go_out;
wire _guard2894 = _guard2892 & _guard2893;
wire _guard2895 = cond_wire672_out;
wire _guard2896 = early_reset_static_par0_go_out;
wire _guard2897 = _guard2895 & _guard2896;
wire _guard2898 = cond_wire692_out;
wire _guard2899 = early_reset_static_par0_go_out;
wire _guard2900 = _guard2898 & _guard2899;
wire _guard2901 = fsm_out == 1'd0;
wire _guard2902 = cond_wire798_out;
wire _guard2903 = _guard2901 & _guard2902;
wire _guard2904 = fsm_out == 1'd0;
wire _guard2905 = _guard2903 & _guard2904;
wire _guard2906 = fsm_out == 1'd0;
wire _guard2907 = cond_wire802_out;
wire _guard2908 = _guard2906 & _guard2907;
wire _guard2909 = fsm_out == 1'd0;
wire _guard2910 = _guard2908 & _guard2909;
wire _guard2911 = _guard2905 | _guard2910;
wire _guard2912 = fsm_out == 1'd0;
wire _guard2913 = cond_wire806_out;
wire _guard2914 = _guard2912 & _guard2913;
wire _guard2915 = fsm_out == 1'd0;
wire _guard2916 = _guard2914 & _guard2915;
wire _guard2917 = _guard2911 | _guard2916;
wire _guard2918 = fsm_out == 1'd0;
wire _guard2919 = cond_wire810_out;
wire _guard2920 = _guard2918 & _guard2919;
wire _guard2921 = fsm_out == 1'd0;
wire _guard2922 = _guard2920 & _guard2921;
wire _guard2923 = _guard2917 | _guard2922;
wire _guard2924 = fsm_out == 1'd0;
wire _guard2925 = cond_wire814_out;
wire _guard2926 = _guard2924 & _guard2925;
wire _guard2927 = fsm_out == 1'd0;
wire _guard2928 = _guard2926 & _guard2927;
wire _guard2929 = _guard2923 | _guard2928;
wire _guard2930 = fsm_out == 1'd0;
wire _guard2931 = cond_wire818_out;
wire _guard2932 = _guard2930 & _guard2931;
wire _guard2933 = fsm_out == 1'd0;
wire _guard2934 = _guard2932 & _guard2933;
wire _guard2935 = _guard2929 | _guard2934;
wire _guard2936 = fsm_out == 1'd0;
wire _guard2937 = cond_wire822_out;
wire _guard2938 = _guard2936 & _guard2937;
wire _guard2939 = fsm_out == 1'd0;
wire _guard2940 = _guard2938 & _guard2939;
wire _guard2941 = _guard2935 | _guard2940;
wire _guard2942 = fsm_out == 1'd0;
wire _guard2943 = cond_wire826_out;
wire _guard2944 = _guard2942 & _guard2943;
wire _guard2945 = fsm_out == 1'd0;
wire _guard2946 = _guard2944 & _guard2945;
wire _guard2947 = _guard2941 | _guard2946;
wire _guard2948 = fsm_out == 1'd0;
wire _guard2949 = cond_wire830_out;
wire _guard2950 = _guard2948 & _guard2949;
wire _guard2951 = fsm_out == 1'd0;
wire _guard2952 = _guard2950 & _guard2951;
wire _guard2953 = _guard2947 | _guard2952;
wire _guard2954 = fsm_out == 1'd0;
wire _guard2955 = cond_wire834_out;
wire _guard2956 = _guard2954 & _guard2955;
wire _guard2957 = fsm_out == 1'd0;
wire _guard2958 = _guard2956 & _guard2957;
wire _guard2959 = _guard2953 | _guard2958;
wire _guard2960 = fsm_out == 1'd0;
wire _guard2961 = cond_wire838_out;
wire _guard2962 = _guard2960 & _guard2961;
wire _guard2963 = fsm_out == 1'd0;
wire _guard2964 = _guard2962 & _guard2963;
wire _guard2965 = _guard2959 | _guard2964;
wire _guard2966 = fsm_out == 1'd0;
wire _guard2967 = cond_wire842_out;
wire _guard2968 = _guard2966 & _guard2967;
wire _guard2969 = fsm_out == 1'd0;
wire _guard2970 = _guard2968 & _guard2969;
wire _guard2971 = _guard2965 | _guard2970;
wire _guard2972 = fsm_out == 1'd0;
wire _guard2973 = cond_wire846_out;
wire _guard2974 = _guard2972 & _guard2973;
wire _guard2975 = fsm_out == 1'd0;
wire _guard2976 = _guard2974 & _guard2975;
wire _guard2977 = _guard2971 | _guard2976;
wire _guard2978 = fsm_out == 1'd0;
wire _guard2979 = cond_wire850_out;
wire _guard2980 = _guard2978 & _guard2979;
wire _guard2981 = fsm_out == 1'd0;
wire _guard2982 = _guard2980 & _guard2981;
wire _guard2983 = _guard2977 | _guard2982;
wire _guard2984 = fsm_out == 1'd0;
wire _guard2985 = cond_wire854_out;
wire _guard2986 = _guard2984 & _guard2985;
wire _guard2987 = fsm_out == 1'd0;
wire _guard2988 = _guard2986 & _guard2987;
wire _guard2989 = _guard2983 | _guard2988;
wire _guard2990 = fsm_out == 1'd0;
wire _guard2991 = cond_wire858_out;
wire _guard2992 = _guard2990 & _guard2991;
wire _guard2993 = fsm_out == 1'd0;
wire _guard2994 = _guard2992 & _guard2993;
wire _guard2995 = _guard2989 | _guard2994;
wire _guard2996 = early_reset_static_par0_go_out;
wire _guard2997 = _guard2995 & _guard2996;
wire _guard2998 = cond_wire24_out;
wire _guard2999 = early_reset_static_par0_go_out;
wire _guard3000 = _guard2998 & _guard2999;
wire _guard3001 = cond_wire74_out;
wire _guard3002 = early_reset_static_par0_go_out;
wire _guard3003 = _guard3001 & _guard3002;
wire _guard3004 = cond_wire79_out;
wire _guard3005 = early_reset_static_par0_go_out;
wire _guard3006 = _guard3004 & _guard3005;
wire _guard3007 = fsm_out == 1'd0;
wire _guard3008 = cond_wire343_out;
wire _guard3009 = _guard3007 & _guard3008;
wire _guard3010 = fsm_out == 1'd0;
wire _guard3011 = _guard3009 & _guard3010;
wire _guard3012 = fsm_out == 1'd0;
wire _guard3013 = cond_wire347_out;
wire _guard3014 = _guard3012 & _guard3013;
wire _guard3015 = fsm_out == 1'd0;
wire _guard3016 = _guard3014 & _guard3015;
wire _guard3017 = _guard3011 | _guard3016;
wire _guard3018 = fsm_out == 1'd0;
wire _guard3019 = cond_wire351_out;
wire _guard3020 = _guard3018 & _guard3019;
wire _guard3021 = fsm_out == 1'd0;
wire _guard3022 = _guard3020 & _guard3021;
wire _guard3023 = _guard3017 | _guard3022;
wire _guard3024 = fsm_out == 1'd0;
wire _guard3025 = cond_wire355_out;
wire _guard3026 = _guard3024 & _guard3025;
wire _guard3027 = fsm_out == 1'd0;
wire _guard3028 = _guard3026 & _guard3027;
wire _guard3029 = _guard3023 | _guard3028;
wire _guard3030 = fsm_out == 1'd0;
wire _guard3031 = cond_wire359_out;
wire _guard3032 = _guard3030 & _guard3031;
wire _guard3033 = fsm_out == 1'd0;
wire _guard3034 = _guard3032 & _guard3033;
wire _guard3035 = _guard3029 | _guard3034;
wire _guard3036 = fsm_out == 1'd0;
wire _guard3037 = cond_wire363_out;
wire _guard3038 = _guard3036 & _guard3037;
wire _guard3039 = fsm_out == 1'd0;
wire _guard3040 = _guard3038 & _guard3039;
wire _guard3041 = _guard3035 | _guard3040;
wire _guard3042 = fsm_out == 1'd0;
wire _guard3043 = cond_wire367_out;
wire _guard3044 = _guard3042 & _guard3043;
wire _guard3045 = fsm_out == 1'd0;
wire _guard3046 = _guard3044 & _guard3045;
wire _guard3047 = _guard3041 | _guard3046;
wire _guard3048 = fsm_out == 1'd0;
wire _guard3049 = cond_wire371_out;
wire _guard3050 = _guard3048 & _guard3049;
wire _guard3051 = fsm_out == 1'd0;
wire _guard3052 = _guard3050 & _guard3051;
wire _guard3053 = _guard3047 | _guard3052;
wire _guard3054 = fsm_out == 1'd0;
wire _guard3055 = cond_wire375_out;
wire _guard3056 = _guard3054 & _guard3055;
wire _guard3057 = fsm_out == 1'd0;
wire _guard3058 = _guard3056 & _guard3057;
wire _guard3059 = _guard3053 | _guard3058;
wire _guard3060 = fsm_out == 1'd0;
wire _guard3061 = cond_wire379_out;
wire _guard3062 = _guard3060 & _guard3061;
wire _guard3063 = fsm_out == 1'd0;
wire _guard3064 = _guard3062 & _guard3063;
wire _guard3065 = _guard3059 | _guard3064;
wire _guard3066 = fsm_out == 1'd0;
wire _guard3067 = cond_wire383_out;
wire _guard3068 = _guard3066 & _guard3067;
wire _guard3069 = fsm_out == 1'd0;
wire _guard3070 = _guard3068 & _guard3069;
wire _guard3071 = _guard3065 | _guard3070;
wire _guard3072 = fsm_out == 1'd0;
wire _guard3073 = cond_wire387_out;
wire _guard3074 = _guard3072 & _guard3073;
wire _guard3075 = fsm_out == 1'd0;
wire _guard3076 = _guard3074 & _guard3075;
wire _guard3077 = _guard3071 | _guard3076;
wire _guard3078 = fsm_out == 1'd0;
wire _guard3079 = cond_wire391_out;
wire _guard3080 = _guard3078 & _guard3079;
wire _guard3081 = fsm_out == 1'd0;
wire _guard3082 = _guard3080 & _guard3081;
wire _guard3083 = _guard3077 | _guard3082;
wire _guard3084 = fsm_out == 1'd0;
wire _guard3085 = cond_wire395_out;
wire _guard3086 = _guard3084 & _guard3085;
wire _guard3087 = fsm_out == 1'd0;
wire _guard3088 = _guard3086 & _guard3087;
wire _guard3089 = _guard3083 | _guard3088;
wire _guard3090 = fsm_out == 1'd0;
wire _guard3091 = cond_wire399_out;
wire _guard3092 = _guard3090 & _guard3091;
wire _guard3093 = fsm_out == 1'd0;
wire _guard3094 = _guard3092 & _guard3093;
wire _guard3095 = _guard3089 | _guard3094;
wire _guard3096 = fsm_out == 1'd0;
wire _guard3097 = cond_wire403_out;
wire _guard3098 = _guard3096 & _guard3097;
wire _guard3099 = fsm_out == 1'd0;
wire _guard3100 = _guard3098 & _guard3099;
wire _guard3101 = _guard3095 | _guard3100;
wire _guard3102 = early_reset_static_par0_go_out;
wire _guard3103 = _guard3101 & _guard3102;
wire _guard3104 = cond_wire477_out;
wire _guard3105 = early_reset_static_par0_go_out;
wire _guard3106 = _guard3104 & _guard3105;
wire _guard3107 = cond_wire533_out;
wire _guard3108 = early_reset_static_par0_go_out;
wire _guard3109 = _guard3107 & _guard3108;
wire _guard3110 = cond_wire473_out;
wire _guard3111 = early_reset_static_par0_go_out;
wire _guard3112 = _guard3110 & _guard3111;
wire _guard3113 = cond_wire485_out;
wire _guard3114 = early_reset_static_par0_go_out;
wire _guard3115 = _guard3113 & _guard3114;
wire _guard3116 = cond_wire525_out;
wire _guard3117 = early_reset_static_par0_go_out;
wire _guard3118 = _guard3116 & _guard3117;
wire _guard3119 = cond_wire529_out;
wire _guard3120 = early_reset_static_par0_go_out;
wire _guard3121 = _guard3119 & _guard3120;
wire _guard3122 = cond_wire493_out;
wire _guard3123 = early_reset_static_par0_go_out;
wire _guard3124 = _guard3122 & _guard3123;
wire _guard3125 = cond_wire521_out;
wire _guard3126 = early_reset_static_par0_go_out;
wire _guard3127 = _guard3125 & _guard3126;
wire _guard3128 = cond_wire481_out;
wire _guard3129 = early_reset_static_par0_go_out;
wire _guard3130 = _guard3128 & _guard3129;
wire _guard3131 = cond_wire505_out;
wire _guard3132 = early_reset_static_par0_go_out;
wire _guard3133 = _guard3131 & _guard3132;
wire _guard3134 = cond_wire513_out;
wire _guard3135 = early_reset_static_par0_go_out;
wire _guard3136 = _guard3134 & _guard3135;
wire _guard3137 = cond_wire501_out;
wire _guard3138 = early_reset_static_par0_go_out;
wire _guard3139 = _guard3137 & _guard3138;
wire _guard3140 = cond_wire517_out;
wire _guard3141 = early_reset_static_par0_go_out;
wire _guard3142 = _guard3140 & _guard3141;
wire _guard3143 = cond_wire489_out;
wire _guard3144 = early_reset_static_par0_go_out;
wire _guard3145 = _guard3143 & _guard3144;
wire _guard3146 = cond_wire497_out;
wire _guard3147 = early_reset_static_par0_go_out;
wire _guard3148 = _guard3146 & _guard3147;
wire _guard3149 = cond_wire509_out;
wire _guard3150 = early_reset_static_par0_go_out;
wire _guard3151 = _guard3149 & _guard3150;
wire _guard3152 = cond_wire607_out;
wire _guard3153 = early_reset_static_par0_go_out;
wire _guard3154 = _guard3152 & _guard3153;
wire _guard3155 = cond_wire663_out;
wire _guard3156 = early_reset_static_par0_go_out;
wire _guard3157 = _guard3155 & _guard3156;
wire _guard3158 = cond_wire603_out;
wire _guard3159 = early_reset_static_par0_go_out;
wire _guard3160 = _guard3158 & _guard3159;
wire _guard3161 = cond_wire615_out;
wire _guard3162 = early_reset_static_par0_go_out;
wire _guard3163 = _guard3161 & _guard3162;
wire _guard3164 = cond_wire655_out;
wire _guard3165 = early_reset_static_par0_go_out;
wire _guard3166 = _guard3164 & _guard3165;
wire _guard3167 = cond_wire659_out;
wire _guard3168 = early_reset_static_par0_go_out;
wire _guard3169 = _guard3167 & _guard3168;
wire _guard3170 = cond_wire623_out;
wire _guard3171 = early_reset_static_par0_go_out;
wire _guard3172 = _guard3170 & _guard3171;
wire _guard3173 = cond_wire651_out;
wire _guard3174 = early_reset_static_par0_go_out;
wire _guard3175 = _guard3173 & _guard3174;
wire _guard3176 = cond_wire611_out;
wire _guard3177 = early_reset_static_par0_go_out;
wire _guard3178 = _guard3176 & _guard3177;
wire _guard3179 = cond_wire635_out;
wire _guard3180 = early_reset_static_par0_go_out;
wire _guard3181 = _guard3179 & _guard3180;
wire _guard3182 = cond_wire643_out;
wire _guard3183 = early_reset_static_par0_go_out;
wire _guard3184 = _guard3182 & _guard3183;
wire _guard3185 = cond_wire631_out;
wire _guard3186 = early_reset_static_par0_go_out;
wire _guard3187 = _guard3185 & _guard3186;
wire _guard3188 = cond_wire647_out;
wire _guard3189 = early_reset_static_par0_go_out;
wire _guard3190 = _guard3188 & _guard3189;
wire _guard3191 = cond_wire619_out;
wire _guard3192 = early_reset_static_par0_go_out;
wire _guard3193 = _guard3191 & _guard3192;
wire _guard3194 = cond_wire627_out;
wire _guard3195 = early_reset_static_par0_go_out;
wire _guard3196 = _guard3194 & _guard3195;
wire _guard3197 = cond_wire639_out;
wire _guard3198 = early_reset_static_par0_go_out;
wire _guard3199 = _guard3197 & _guard3198;
wire _guard3200 = fsm_out == 1'd0;
wire _guard3201 = cond_wire863_out;
wire _guard3202 = _guard3200 & _guard3201;
wire _guard3203 = fsm_out == 1'd0;
wire _guard3204 = _guard3202 & _guard3203;
wire _guard3205 = fsm_out == 1'd0;
wire _guard3206 = cond_wire867_out;
wire _guard3207 = _guard3205 & _guard3206;
wire _guard3208 = fsm_out == 1'd0;
wire _guard3209 = _guard3207 & _guard3208;
wire _guard3210 = _guard3204 | _guard3209;
wire _guard3211 = fsm_out == 1'd0;
wire _guard3212 = cond_wire871_out;
wire _guard3213 = _guard3211 & _guard3212;
wire _guard3214 = fsm_out == 1'd0;
wire _guard3215 = _guard3213 & _guard3214;
wire _guard3216 = _guard3210 | _guard3215;
wire _guard3217 = fsm_out == 1'd0;
wire _guard3218 = cond_wire875_out;
wire _guard3219 = _guard3217 & _guard3218;
wire _guard3220 = fsm_out == 1'd0;
wire _guard3221 = _guard3219 & _guard3220;
wire _guard3222 = _guard3216 | _guard3221;
wire _guard3223 = fsm_out == 1'd0;
wire _guard3224 = cond_wire879_out;
wire _guard3225 = _guard3223 & _guard3224;
wire _guard3226 = fsm_out == 1'd0;
wire _guard3227 = _guard3225 & _guard3226;
wire _guard3228 = _guard3222 | _guard3227;
wire _guard3229 = fsm_out == 1'd0;
wire _guard3230 = cond_wire883_out;
wire _guard3231 = _guard3229 & _guard3230;
wire _guard3232 = fsm_out == 1'd0;
wire _guard3233 = _guard3231 & _guard3232;
wire _guard3234 = _guard3228 | _guard3233;
wire _guard3235 = fsm_out == 1'd0;
wire _guard3236 = cond_wire887_out;
wire _guard3237 = _guard3235 & _guard3236;
wire _guard3238 = fsm_out == 1'd0;
wire _guard3239 = _guard3237 & _guard3238;
wire _guard3240 = _guard3234 | _guard3239;
wire _guard3241 = fsm_out == 1'd0;
wire _guard3242 = cond_wire891_out;
wire _guard3243 = _guard3241 & _guard3242;
wire _guard3244 = fsm_out == 1'd0;
wire _guard3245 = _guard3243 & _guard3244;
wire _guard3246 = _guard3240 | _guard3245;
wire _guard3247 = fsm_out == 1'd0;
wire _guard3248 = cond_wire895_out;
wire _guard3249 = _guard3247 & _guard3248;
wire _guard3250 = fsm_out == 1'd0;
wire _guard3251 = _guard3249 & _guard3250;
wire _guard3252 = _guard3246 | _guard3251;
wire _guard3253 = fsm_out == 1'd0;
wire _guard3254 = cond_wire899_out;
wire _guard3255 = _guard3253 & _guard3254;
wire _guard3256 = fsm_out == 1'd0;
wire _guard3257 = _guard3255 & _guard3256;
wire _guard3258 = _guard3252 | _guard3257;
wire _guard3259 = fsm_out == 1'd0;
wire _guard3260 = cond_wire903_out;
wire _guard3261 = _guard3259 & _guard3260;
wire _guard3262 = fsm_out == 1'd0;
wire _guard3263 = _guard3261 & _guard3262;
wire _guard3264 = _guard3258 | _guard3263;
wire _guard3265 = fsm_out == 1'd0;
wire _guard3266 = cond_wire907_out;
wire _guard3267 = _guard3265 & _guard3266;
wire _guard3268 = fsm_out == 1'd0;
wire _guard3269 = _guard3267 & _guard3268;
wire _guard3270 = _guard3264 | _guard3269;
wire _guard3271 = fsm_out == 1'd0;
wire _guard3272 = cond_wire911_out;
wire _guard3273 = _guard3271 & _guard3272;
wire _guard3274 = fsm_out == 1'd0;
wire _guard3275 = _guard3273 & _guard3274;
wire _guard3276 = _guard3270 | _guard3275;
wire _guard3277 = fsm_out == 1'd0;
wire _guard3278 = cond_wire915_out;
wire _guard3279 = _guard3277 & _guard3278;
wire _guard3280 = fsm_out == 1'd0;
wire _guard3281 = _guard3279 & _guard3280;
wire _guard3282 = _guard3276 | _guard3281;
wire _guard3283 = fsm_out == 1'd0;
wire _guard3284 = cond_wire919_out;
wire _guard3285 = _guard3283 & _guard3284;
wire _guard3286 = fsm_out == 1'd0;
wire _guard3287 = _guard3285 & _guard3286;
wire _guard3288 = _guard3282 | _guard3287;
wire _guard3289 = fsm_out == 1'd0;
wire _guard3290 = cond_wire923_out;
wire _guard3291 = _guard3289 & _guard3290;
wire _guard3292 = fsm_out == 1'd0;
wire _guard3293 = _guard3291 & _guard3292;
wire _guard3294 = _guard3288 | _guard3293;
wire _guard3295 = early_reset_static_par0_go_out;
wire _guard3296 = _guard3294 & _guard3295;
wire _guard3297 = cond_wire69_out;
wire _guard3298 = early_reset_static_par0_go_out;
wire _guard3299 = _guard3297 & _guard3298;
wire _guard3300 = cond_wire672_out;
wire _guard3301 = early_reset_static_par0_go_out;
wire _guard3302 = _guard3300 & _guard3301;
wire _guard3303 = cond_wire728_out;
wire _guard3304 = early_reset_static_par0_go_out;
wire _guard3305 = _guard3303 & _guard3304;
wire _guard3306 = cond_wire668_out;
wire _guard3307 = early_reset_static_par0_go_out;
wire _guard3308 = _guard3306 & _guard3307;
wire _guard3309 = cond_wire680_out;
wire _guard3310 = early_reset_static_par0_go_out;
wire _guard3311 = _guard3309 & _guard3310;
wire _guard3312 = cond_wire720_out;
wire _guard3313 = early_reset_static_par0_go_out;
wire _guard3314 = _guard3312 & _guard3313;
wire _guard3315 = cond_wire724_out;
wire _guard3316 = early_reset_static_par0_go_out;
wire _guard3317 = _guard3315 & _guard3316;
wire _guard3318 = cond_wire688_out;
wire _guard3319 = early_reset_static_par0_go_out;
wire _guard3320 = _guard3318 & _guard3319;
wire _guard3321 = cond_wire716_out;
wire _guard3322 = early_reset_static_par0_go_out;
wire _guard3323 = _guard3321 & _guard3322;
wire _guard3324 = cond_wire676_out;
wire _guard3325 = early_reset_static_par0_go_out;
wire _guard3326 = _guard3324 & _guard3325;
wire _guard3327 = cond_wire700_out;
wire _guard3328 = early_reset_static_par0_go_out;
wire _guard3329 = _guard3327 & _guard3328;
wire _guard3330 = cond_wire708_out;
wire _guard3331 = early_reset_static_par0_go_out;
wire _guard3332 = _guard3330 & _guard3331;
wire _guard3333 = cond_wire696_out;
wire _guard3334 = early_reset_static_par0_go_out;
wire _guard3335 = _guard3333 & _guard3334;
wire _guard3336 = cond_wire712_out;
wire _guard3337 = early_reset_static_par0_go_out;
wire _guard3338 = _guard3336 & _guard3337;
wire _guard3339 = cond_wire684_out;
wire _guard3340 = early_reset_static_par0_go_out;
wire _guard3341 = _guard3339 & _guard3340;
wire _guard3342 = cond_wire692_out;
wire _guard3343 = early_reset_static_par0_go_out;
wire _guard3344 = _guard3342 & _guard3343;
wire _guard3345 = cond_wire704_out;
wire _guard3346 = early_reset_static_par0_go_out;
wire _guard3347 = _guard3345 & _guard3346;
wire _guard3348 = cond_wire19_out;
wire _guard3349 = early_reset_static_par0_go_out;
wire _guard3350 = _guard3348 & _guard3349;
wire _guard3351 = cond_wire29_out;
wire _guard3352 = early_reset_static_par0_go_out;
wire _guard3353 = _guard3351 & _guard3352;
wire _guard3354 = cond_wire59_out;
wire _guard3355 = early_reset_static_par0_go_out;
wire _guard3356 = _guard3354 & _guard3355;
wire _guard3357 = fsm_out == 1'd0;
wire _guard3358 = cond_wire473_out;
wire _guard3359 = _guard3357 & _guard3358;
wire _guard3360 = fsm_out == 1'd0;
wire _guard3361 = _guard3359 & _guard3360;
wire _guard3362 = fsm_out == 1'd0;
wire _guard3363 = cond_wire477_out;
wire _guard3364 = _guard3362 & _guard3363;
wire _guard3365 = fsm_out == 1'd0;
wire _guard3366 = _guard3364 & _guard3365;
wire _guard3367 = _guard3361 | _guard3366;
wire _guard3368 = fsm_out == 1'd0;
wire _guard3369 = cond_wire481_out;
wire _guard3370 = _guard3368 & _guard3369;
wire _guard3371 = fsm_out == 1'd0;
wire _guard3372 = _guard3370 & _guard3371;
wire _guard3373 = _guard3367 | _guard3372;
wire _guard3374 = fsm_out == 1'd0;
wire _guard3375 = cond_wire485_out;
wire _guard3376 = _guard3374 & _guard3375;
wire _guard3377 = fsm_out == 1'd0;
wire _guard3378 = _guard3376 & _guard3377;
wire _guard3379 = _guard3373 | _guard3378;
wire _guard3380 = fsm_out == 1'd0;
wire _guard3381 = cond_wire489_out;
wire _guard3382 = _guard3380 & _guard3381;
wire _guard3383 = fsm_out == 1'd0;
wire _guard3384 = _guard3382 & _guard3383;
wire _guard3385 = _guard3379 | _guard3384;
wire _guard3386 = fsm_out == 1'd0;
wire _guard3387 = cond_wire493_out;
wire _guard3388 = _guard3386 & _guard3387;
wire _guard3389 = fsm_out == 1'd0;
wire _guard3390 = _guard3388 & _guard3389;
wire _guard3391 = _guard3385 | _guard3390;
wire _guard3392 = fsm_out == 1'd0;
wire _guard3393 = cond_wire497_out;
wire _guard3394 = _guard3392 & _guard3393;
wire _guard3395 = fsm_out == 1'd0;
wire _guard3396 = _guard3394 & _guard3395;
wire _guard3397 = _guard3391 | _guard3396;
wire _guard3398 = fsm_out == 1'd0;
wire _guard3399 = cond_wire501_out;
wire _guard3400 = _guard3398 & _guard3399;
wire _guard3401 = fsm_out == 1'd0;
wire _guard3402 = _guard3400 & _guard3401;
wire _guard3403 = _guard3397 | _guard3402;
wire _guard3404 = fsm_out == 1'd0;
wire _guard3405 = cond_wire505_out;
wire _guard3406 = _guard3404 & _guard3405;
wire _guard3407 = fsm_out == 1'd0;
wire _guard3408 = _guard3406 & _guard3407;
wire _guard3409 = _guard3403 | _guard3408;
wire _guard3410 = fsm_out == 1'd0;
wire _guard3411 = cond_wire509_out;
wire _guard3412 = _guard3410 & _guard3411;
wire _guard3413 = fsm_out == 1'd0;
wire _guard3414 = _guard3412 & _guard3413;
wire _guard3415 = _guard3409 | _guard3414;
wire _guard3416 = fsm_out == 1'd0;
wire _guard3417 = cond_wire513_out;
wire _guard3418 = _guard3416 & _guard3417;
wire _guard3419 = fsm_out == 1'd0;
wire _guard3420 = _guard3418 & _guard3419;
wire _guard3421 = _guard3415 | _guard3420;
wire _guard3422 = fsm_out == 1'd0;
wire _guard3423 = cond_wire517_out;
wire _guard3424 = _guard3422 & _guard3423;
wire _guard3425 = fsm_out == 1'd0;
wire _guard3426 = _guard3424 & _guard3425;
wire _guard3427 = _guard3421 | _guard3426;
wire _guard3428 = fsm_out == 1'd0;
wire _guard3429 = cond_wire521_out;
wire _guard3430 = _guard3428 & _guard3429;
wire _guard3431 = fsm_out == 1'd0;
wire _guard3432 = _guard3430 & _guard3431;
wire _guard3433 = _guard3427 | _guard3432;
wire _guard3434 = fsm_out == 1'd0;
wire _guard3435 = cond_wire525_out;
wire _guard3436 = _guard3434 & _guard3435;
wire _guard3437 = fsm_out == 1'd0;
wire _guard3438 = _guard3436 & _guard3437;
wire _guard3439 = _guard3433 | _guard3438;
wire _guard3440 = fsm_out == 1'd0;
wire _guard3441 = cond_wire529_out;
wire _guard3442 = _guard3440 & _guard3441;
wire _guard3443 = fsm_out == 1'd0;
wire _guard3444 = _guard3442 & _guard3443;
wire _guard3445 = _guard3439 | _guard3444;
wire _guard3446 = fsm_out == 1'd0;
wire _guard3447 = cond_wire533_out;
wire _guard3448 = _guard3446 & _guard3447;
wire _guard3449 = fsm_out == 1'd0;
wire _guard3450 = _guard3448 & _guard3449;
wire _guard3451 = _guard3445 | _guard3450;
wire _guard3452 = early_reset_static_par0_go_out;
wire _guard3453 = _guard3451 & _guard3452;
wire _guard3454 = cond_wire39_out;
wire _guard3455 = early_reset_static_par0_go_out;
wire _guard3456 = _guard3454 & _guard3455;
wire _guard3457 = cond_wire282_out;
wire _guard3458 = early_reset_static_par0_go_out;
wire _guard3459 = _guard3457 & _guard3458;
wire _guard3460 = cond_wire338_out;
wire _guard3461 = early_reset_static_par0_go_out;
wire _guard3462 = _guard3460 & _guard3461;
wire _guard3463 = cond_wire278_out;
wire _guard3464 = early_reset_static_par0_go_out;
wire _guard3465 = _guard3463 & _guard3464;
wire _guard3466 = cond_wire290_out;
wire _guard3467 = early_reset_static_par0_go_out;
wire _guard3468 = _guard3466 & _guard3467;
wire _guard3469 = cond_wire330_out;
wire _guard3470 = early_reset_static_par0_go_out;
wire _guard3471 = _guard3469 & _guard3470;
wire _guard3472 = cond_wire334_out;
wire _guard3473 = early_reset_static_par0_go_out;
wire _guard3474 = _guard3472 & _guard3473;
wire _guard3475 = cond_wire298_out;
wire _guard3476 = early_reset_static_par0_go_out;
wire _guard3477 = _guard3475 & _guard3476;
wire _guard3478 = cond_wire326_out;
wire _guard3479 = early_reset_static_par0_go_out;
wire _guard3480 = _guard3478 & _guard3479;
wire _guard3481 = cond_wire286_out;
wire _guard3482 = early_reset_static_par0_go_out;
wire _guard3483 = _guard3481 & _guard3482;
wire _guard3484 = cond_wire310_out;
wire _guard3485 = early_reset_static_par0_go_out;
wire _guard3486 = _guard3484 & _guard3485;
wire _guard3487 = cond_wire318_out;
wire _guard3488 = early_reset_static_par0_go_out;
wire _guard3489 = _guard3487 & _guard3488;
wire _guard3490 = cond_wire306_out;
wire _guard3491 = early_reset_static_par0_go_out;
wire _guard3492 = _guard3490 & _guard3491;
wire _guard3493 = cond_wire322_out;
wire _guard3494 = early_reset_static_par0_go_out;
wire _guard3495 = _guard3493 & _guard3494;
wire _guard3496 = cond_wire294_out;
wire _guard3497 = early_reset_static_par0_go_out;
wire _guard3498 = _guard3496 & _guard3497;
wire _guard3499 = cond_wire302_out;
wire _guard3500 = early_reset_static_par0_go_out;
wire _guard3501 = _guard3499 & _guard3500;
wire _guard3502 = cond_wire314_out;
wire _guard3503 = early_reset_static_par0_go_out;
wire _guard3504 = _guard3502 & _guard3503;
wire _guard3505 = fsm_out == 1'd0;
wire _guard3506 = cond_wire733_out;
wire _guard3507 = _guard3505 & _guard3506;
wire _guard3508 = fsm_out == 1'd0;
wire _guard3509 = _guard3507 & _guard3508;
wire _guard3510 = fsm_out == 1'd0;
wire _guard3511 = cond_wire737_out;
wire _guard3512 = _guard3510 & _guard3511;
wire _guard3513 = fsm_out == 1'd0;
wire _guard3514 = _guard3512 & _guard3513;
wire _guard3515 = _guard3509 | _guard3514;
wire _guard3516 = fsm_out == 1'd0;
wire _guard3517 = cond_wire741_out;
wire _guard3518 = _guard3516 & _guard3517;
wire _guard3519 = fsm_out == 1'd0;
wire _guard3520 = _guard3518 & _guard3519;
wire _guard3521 = _guard3515 | _guard3520;
wire _guard3522 = fsm_out == 1'd0;
wire _guard3523 = cond_wire745_out;
wire _guard3524 = _guard3522 & _guard3523;
wire _guard3525 = fsm_out == 1'd0;
wire _guard3526 = _guard3524 & _guard3525;
wire _guard3527 = _guard3521 | _guard3526;
wire _guard3528 = fsm_out == 1'd0;
wire _guard3529 = cond_wire749_out;
wire _guard3530 = _guard3528 & _guard3529;
wire _guard3531 = fsm_out == 1'd0;
wire _guard3532 = _guard3530 & _guard3531;
wire _guard3533 = _guard3527 | _guard3532;
wire _guard3534 = fsm_out == 1'd0;
wire _guard3535 = cond_wire753_out;
wire _guard3536 = _guard3534 & _guard3535;
wire _guard3537 = fsm_out == 1'd0;
wire _guard3538 = _guard3536 & _guard3537;
wire _guard3539 = _guard3533 | _guard3538;
wire _guard3540 = fsm_out == 1'd0;
wire _guard3541 = cond_wire757_out;
wire _guard3542 = _guard3540 & _guard3541;
wire _guard3543 = fsm_out == 1'd0;
wire _guard3544 = _guard3542 & _guard3543;
wire _guard3545 = _guard3539 | _guard3544;
wire _guard3546 = fsm_out == 1'd0;
wire _guard3547 = cond_wire761_out;
wire _guard3548 = _guard3546 & _guard3547;
wire _guard3549 = fsm_out == 1'd0;
wire _guard3550 = _guard3548 & _guard3549;
wire _guard3551 = _guard3545 | _guard3550;
wire _guard3552 = fsm_out == 1'd0;
wire _guard3553 = cond_wire765_out;
wire _guard3554 = _guard3552 & _guard3553;
wire _guard3555 = fsm_out == 1'd0;
wire _guard3556 = _guard3554 & _guard3555;
wire _guard3557 = _guard3551 | _guard3556;
wire _guard3558 = fsm_out == 1'd0;
wire _guard3559 = cond_wire769_out;
wire _guard3560 = _guard3558 & _guard3559;
wire _guard3561 = fsm_out == 1'd0;
wire _guard3562 = _guard3560 & _guard3561;
wire _guard3563 = _guard3557 | _guard3562;
wire _guard3564 = fsm_out == 1'd0;
wire _guard3565 = cond_wire773_out;
wire _guard3566 = _guard3564 & _guard3565;
wire _guard3567 = fsm_out == 1'd0;
wire _guard3568 = _guard3566 & _guard3567;
wire _guard3569 = _guard3563 | _guard3568;
wire _guard3570 = fsm_out == 1'd0;
wire _guard3571 = cond_wire777_out;
wire _guard3572 = _guard3570 & _guard3571;
wire _guard3573 = fsm_out == 1'd0;
wire _guard3574 = _guard3572 & _guard3573;
wire _guard3575 = _guard3569 | _guard3574;
wire _guard3576 = fsm_out == 1'd0;
wire _guard3577 = cond_wire781_out;
wire _guard3578 = _guard3576 & _guard3577;
wire _guard3579 = fsm_out == 1'd0;
wire _guard3580 = _guard3578 & _guard3579;
wire _guard3581 = _guard3575 | _guard3580;
wire _guard3582 = fsm_out == 1'd0;
wire _guard3583 = cond_wire785_out;
wire _guard3584 = _guard3582 & _guard3583;
wire _guard3585 = fsm_out == 1'd0;
wire _guard3586 = _guard3584 & _guard3585;
wire _guard3587 = _guard3581 | _guard3586;
wire _guard3588 = fsm_out == 1'd0;
wire _guard3589 = cond_wire789_out;
wire _guard3590 = _guard3588 & _guard3589;
wire _guard3591 = fsm_out == 1'd0;
wire _guard3592 = _guard3590 & _guard3591;
wire _guard3593 = _guard3587 | _guard3592;
wire _guard3594 = fsm_out == 1'd0;
wire _guard3595 = cond_wire793_out;
wire _guard3596 = _guard3594 & _guard3595;
wire _guard3597 = fsm_out == 1'd0;
wire _guard3598 = _guard3596 & _guard3597;
wire _guard3599 = _guard3593 | _guard3598;
wire _guard3600 = early_reset_static_par0_go_out;
wire _guard3601 = _guard3599 & _guard3600;
wire _guard3602 = cond_wire44_out;
wire _guard3603 = early_reset_static_par0_go_out;
wire _guard3604 = _guard3602 & _guard3603;
wire _guard3605 = cond_wire209_out;
wire _guard3606 = early_reset_static_par0_go_out;
wire _guard3607 = _guard3605 & _guard3606;
wire _guard3608 = cond_wire664_out;
wire _guard3609 = early_reset_static_par0_go_out;
wire _guard3610 = _guard3608 & _guard3609;
wire _guard3611 = cond_wire196_out;
wire _guard3612 = early_reset_static_par0_go_out;
wire _guard3613 = _guard3611 & _guard3612;
wire _guard3614 = cond_wire192_out;
wire _guard3615 = early_reset_static_par0_go_out;
wire _guard3616 = _guard3614 & _guard3615;
wire _guard3617 = cond_wire204_out;
wire _guard3618 = early_reset_static_par0_go_out;
wire _guard3619 = _guard3617 & _guard3618;
wire _guard3620 = cond_wire176_out;
wire _guard3621 = early_reset_static_par0_go_out;
wire _guard3622 = _guard3620 & _guard3621;
wire _guard3623 = cond_wire200_out;
wire _guard3624 = early_reset_static_par0_go_out;
wire _guard3625 = _guard3623 & _guard3624;
wire _guard3626 = cond_wire164_out;
wire _guard3627 = early_reset_static_par0_go_out;
wire _guard3628 = _guard3626 & _guard3627;
wire _guard3629 = cond_wire208_out;
wire _guard3630 = early_reset_static_par0_go_out;
wire _guard3631 = _guard3629 & _guard3630;
wire _guard3632 = cond_wire152_out;
wire _guard3633 = early_reset_static_par0_go_out;
wire _guard3634 = _guard3632 & _guard3633;
wire _guard3635 = cond_wire160_out;
wire _guard3636 = early_reset_static_par0_go_out;
wire _guard3637 = _guard3635 & _guard3636;
wire _guard3638 = cond_wire168_out;
wire _guard3639 = early_reset_static_par0_go_out;
wire _guard3640 = _guard3638 & _guard3639;
wire _guard3641 = cond_wire172_out;
wire _guard3642 = early_reset_static_par0_go_out;
wire _guard3643 = _guard3641 & _guard3642;
wire _guard3644 = cond_wire180_out;
wire _guard3645 = early_reset_static_par0_go_out;
wire _guard3646 = _guard3644 & _guard3645;
wire _guard3647 = cond_wire148_out;
wire _guard3648 = early_reset_static_par0_go_out;
wire _guard3649 = _guard3647 & _guard3648;
wire _guard3650 = cond_wire156_out;
wire _guard3651 = early_reset_static_par0_go_out;
wire _guard3652 = _guard3650 & _guard3651;
wire _guard3653 = cond_wire184_out;
wire _guard3654 = early_reset_static_par0_go_out;
wire _guard3655 = _guard3653 & _guard3654;
wire _guard3656 = cond_wire188_out;
wire _guard3657 = early_reset_static_par0_go_out;
wire _guard3658 = _guard3656 & _guard3657;
wire _guard3659 = cond_wire274_out;
wire _guard3660 = early_reset_static_par0_go_out;
wire _guard3661 = _guard3659 & _guard3660;
wire _guard3662 = cond_wire469_out;
wire _guard3663 = early_reset_static_par0_go_out;
wire _guard3664 = _guard3662 & _guard3663;
wire _guard3665 = cond_wire99_out;
wire _guard3666 = early_reset_static_par0_go_out;
wire _guard3667 = _guard3665 & _guard3666;
wire _guard3668 = cond_wire111_out;
wire _guard3669 = early_reset_static_par0_go_out;
wire _guard3670 = _guard3668 & _guard3669;
wire _guard3671 = cond_wire91_out;
wire _guard3672 = early_reset_static_par0_go_out;
wire _guard3673 = _guard3671 & _guard3672;
wire _guard3674 = cond_wire95_out;
wire _guard3675 = early_reset_static_par0_go_out;
wire _guard3676 = _guard3674 & _guard3675;
wire _guard3677 = cond_wire115_out;
wire _guard3678 = early_reset_static_par0_go_out;
wire _guard3679 = _guard3677 & _guard3678;
wire _guard3680 = cond_wire143_out;
wire _guard3681 = early_reset_static_par0_go_out;
wire _guard3682 = _guard3680 & _guard3681;
wire _guard3683 = cond_wire83_out;
wire _guard3684 = early_reset_static_par0_go_out;
wire _guard3685 = _guard3683 & _guard3684;
wire _guard3686 = cond_wire107_out;
wire _guard3687 = early_reset_static_par0_go_out;
wire _guard3688 = _guard3686 & _guard3687;
wire _guard3689 = cond_wire131_out;
wire _guard3690 = early_reset_static_par0_go_out;
wire _guard3691 = _guard3689 & _guard3690;
wire _guard3692 = cond_wire103_out;
wire _guard3693 = early_reset_static_par0_go_out;
wire _guard3694 = _guard3692 & _guard3693;
wire _guard3695 = cond_wire119_out;
wire _guard3696 = early_reset_static_par0_go_out;
wire _guard3697 = _guard3695 & _guard3696;
wire _guard3698 = cond_wire127_out;
wire _guard3699 = early_reset_static_par0_go_out;
wire _guard3700 = _guard3698 & _guard3699;
wire _guard3701 = cond_wire87_out;
wire _guard3702 = early_reset_static_par0_go_out;
wire _guard3703 = _guard3701 & _guard3702;
wire _guard3704 = cond_wire135_out;
wire _guard3705 = early_reset_static_par0_go_out;
wire _guard3706 = _guard3704 & _guard3705;
wire _guard3707 = cond_wire123_out;
wire _guard3708 = early_reset_static_par0_go_out;
wire _guard3709 = _guard3707 & _guard3708;
wire _guard3710 = cond_wire139_out;
wire _guard3711 = early_reset_static_par0_go_out;
wire _guard3712 = _guard3710 & _guard3711;
wire _guard3713 = fsm_out == 1'd0;
wire _guard3714 = cond_wire83_out;
wire _guard3715 = _guard3713 & _guard3714;
wire _guard3716 = fsm_out == 1'd0;
wire _guard3717 = _guard3715 & _guard3716;
wire _guard3718 = fsm_out == 1'd0;
wire _guard3719 = cond_wire87_out;
wire _guard3720 = _guard3718 & _guard3719;
wire _guard3721 = fsm_out == 1'd0;
wire _guard3722 = _guard3720 & _guard3721;
wire _guard3723 = _guard3717 | _guard3722;
wire _guard3724 = fsm_out == 1'd0;
wire _guard3725 = cond_wire91_out;
wire _guard3726 = _guard3724 & _guard3725;
wire _guard3727 = fsm_out == 1'd0;
wire _guard3728 = _guard3726 & _guard3727;
wire _guard3729 = _guard3723 | _guard3728;
wire _guard3730 = fsm_out == 1'd0;
wire _guard3731 = cond_wire95_out;
wire _guard3732 = _guard3730 & _guard3731;
wire _guard3733 = fsm_out == 1'd0;
wire _guard3734 = _guard3732 & _guard3733;
wire _guard3735 = _guard3729 | _guard3734;
wire _guard3736 = fsm_out == 1'd0;
wire _guard3737 = cond_wire99_out;
wire _guard3738 = _guard3736 & _guard3737;
wire _guard3739 = fsm_out == 1'd0;
wire _guard3740 = _guard3738 & _guard3739;
wire _guard3741 = _guard3735 | _guard3740;
wire _guard3742 = fsm_out == 1'd0;
wire _guard3743 = cond_wire103_out;
wire _guard3744 = _guard3742 & _guard3743;
wire _guard3745 = fsm_out == 1'd0;
wire _guard3746 = _guard3744 & _guard3745;
wire _guard3747 = _guard3741 | _guard3746;
wire _guard3748 = fsm_out == 1'd0;
wire _guard3749 = cond_wire107_out;
wire _guard3750 = _guard3748 & _guard3749;
wire _guard3751 = fsm_out == 1'd0;
wire _guard3752 = _guard3750 & _guard3751;
wire _guard3753 = _guard3747 | _guard3752;
wire _guard3754 = fsm_out == 1'd0;
wire _guard3755 = cond_wire111_out;
wire _guard3756 = _guard3754 & _guard3755;
wire _guard3757 = fsm_out == 1'd0;
wire _guard3758 = _guard3756 & _guard3757;
wire _guard3759 = _guard3753 | _guard3758;
wire _guard3760 = fsm_out == 1'd0;
wire _guard3761 = cond_wire115_out;
wire _guard3762 = _guard3760 & _guard3761;
wire _guard3763 = fsm_out == 1'd0;
wire _guard3764 = _guard3762 & _guard3763;
wire _guard3765 = _guard3759 | _guard3764;
wire _guard3766 = fsm_out == 1'd0;
wire _guard3767 = cond_wire119_out;
wire _guard3768 = _guard3766 & _guard3767;
wire _guard3769 = fsm_out == 1'd0;
wire _guard3770 = _guard3768 & _guard3769;
wire _guard3771 = _guard3765 | _guard3770;
wire _guard3772 = fsm_out == 1'd0;
wire _guard3773 = cond_wire123_out;
wire _guard3774 = _guard3772 & _guard3773;
wire _guard3775 = fsm_out == 1'd0;
wire _guard3776 = _guard3774 & _guard3775;
wire _guard3777 = _guard3771 | _guard3776;
wire _guard3778 = fsm_out == 1'd0;
wire _guard3779 = cond_wire127_out;
wire _guard3780 = _guard3778 & _guard3779;
wire _guard3781 = fsm_out == 1'd0;
wire _guard3782 = _guard3780 & _guard3781;
wire _guard3783 = _guard3777 | _guard3782;
wire _guard3784 = fsm_out == 1'd0;
wire _guard3785 = cond_wire131_out;
wire _guard3786 = _guard3784 & _guard3785;
wire _guard3787 = fsm_out == 1'd0;
wire _guard3788 = _guard3786 & _guard3787;
wire _guard3789 = _guard3783 | _guard3788;
wire _guard3790 = fsm_out == 1'd0;
wire _guard3791 = cond_wire135_out;
wire _guard3792 = _guard3790 & _guard3791;
wire _guard3793 = fsm_out == 1'd0;
wire _guard3794 = _guard3792 & _guard3793;
wire _guard3795 = _guard3789 | _guard3794;
wire _guard3796 = fsm_out == 1'd0;
wire _guard3797 = cond_wire139_out;
wire _guard3798 = _guard3796 & _guard3797;
wire _guard3799 = fsm_out == 1'd0;
wire _guard3800 = _guard3798 & _guard3799;
wire _guard3801 = _guard3795 | _guard3800;
wire _guard3802 = fsm_out == 1'd0;
wire _guard3803 = cond_wire143_out;
wire _guard3804 = _guard3802 & _guard3803;
wire _guard3805 = fsm_out == 1'd0;
wire _guard3806 = _guard3804 & _guard3805;
wire _guard3807 = _guard3801 | _guard3806;
wire _guard3808 = early_reset_static_par0_go_out;
wire _guard3809 = _guard3807 & _guard3808;
wire _guard3810 = fsm_out == 1'd0;
wire _guard3811 = cond_wire278_out;
wire _guard3812 = _guard3810 & _guard3811;
wire _guard3813 = fsm_out == 1'd0;
wire _guard3814 = _guard3812 & _guard3813;
wire _guard3815 = fsm_out == 1'd0;
wire _guard3816 = cond_wire282_out;
wire _guard3817 = _guard3815 & _guard3816;
wire _guard3818 = fsm_out == 1'd0;
wire _guard3819 = _guard3817 & _guard3818;
wire _guard3820 = _guard3814 | _guard3819;
wire _guard3821 = fsm_out == 1'd0;
wire _guard3822 = cond_wire286_out;
wire _guard3823 = _guard3821 & _guard3822;
wire _guard3824 = fsm_out == 1'd0;
wire _guard3825 = _guard3823 & _guard3824;
wire _guard3826 = _guard3820 | _guard3825;
wire _guard3827 = fsm_out == 1'd0;
wire _guard3828 = cond_wire290_out;
wire _guard3829 = _guard3827 & _guard3828;
wire _guard3830 = fsm_out == 1'd0;
wire _guard3831 = _guard3829 & _guard3830;
wire _guard3832 = _guard3826 | _guard3831;
wire _guard3833 = fsm_out == 1'd0;
wire _guard3834 = cond_wire294_out;
wire _guard3835 = _guard3833 & _guard3834;
wire _guard3836 = fsm_out == 1'd0;
wire _guard3837 = _guard3835 & _guard3836;
wire _guard3838 = _guard3832 | _guard3837;
wire _guard3839 = fsm_out == 1'd0;
wire _guard3840 = cond_wire298_out;
wire _guard3841 = _guard3839 & _guard3840;
wire _guard3842 = fsm_out == 1'd0;
wire _guard3843 = _guard3841 & _guard3842;
wire _guard3844 = _guard3838 | _guard3843;
wire _guard3845 = fsm_out == 1'd0;
wire _guard3846 = cond_wire302_out;
wire _guard3847 = _guard3845 & _guard3846;
wire _guard3848 = fsm_out == 1'd0;
wire _guard3849 = _guard3847 & _guard3848;
wire _guard3850 = _guard3844 | _guard3849;
wire _guard3851 = fsm_out == 1'd0;
wire _guard3852 = cond_wire306_out;
wire _guard3853 = _guard3851 & _guard3852;
wire _guard3854 = fsm_out == 1'd0;
wire _guard3855 = _guard3853 & _guard3854;
wire _guard3856 = _guard3850 | _guard3855;
wire _guard3857 = fsm_out == 1'd0;
wire _guard3858 = cond_wire310_out;
wire _guard3859 = _guard3857 & _guard3858;
wire _guard3860 = fsm_out == 1'd0;
wire _guard3861 = _guard3859 & _guard3860;
wire _guard3862 = _guard3856 | _guard3861;
wire _guard3863 = fsm_out == 1'd0;
wire _guard3864 = cond_wire314_out;
wire _guard3865 = _guard3863 & _guard3864;
wire _guard3866 = fsm_out == 1'd0;
wire _guard3867 = _guard3865 & _guard3866;
wire _guard3868 = _guard3862 | _guard3867;
wire _guard3869 = fsm_out == 1'd0;
wire _guard3870 = cond_wire318_out;
wire _guard3871 = _guard3869 & _guard3870;
wire _guard3872 = fsm_out == 1'd0;
wire _guard3873 = _guard3871 & _guard3872;
wire _guard3874 = _guard3868 | _guard3873;
wire _guard3875 = fsm_out == 1'd0;
wire _guard3876 = cond_wire322_out;
wire _guard3877 = _guard3875 & _guard3876;
wire _guard3878 = fsm_out == 1'd0;
wire _guard3879 = _guard3877 & _guard3878;
wire _guard3880 = _guard3874 | _guard3879;
wire _guard3881 = fsm_out == 1'd0;
wire _guard3882 = cond_wire326_out;
wire _guard3883 = _guard3881 & _guard3882;
wire _guard3884 = fsm_out == 1'd0;
wire _guard3885 = _guard3883 & _guard3884;
wire _guard3886 = _guard3880 | _guard3885;
wire _guard3887 = fsm_out == 1'd0;
wire _guard3888 = cond_wire330_out;
wire _guard3889 = _guard3887 & _guard3888;
wire _guard3890 = fsm_out == 1'd0;
wire _guard3891 = _guard3889 & _guard3890;
wire _guard3892 = _guard3886 | _guard3891;
wire _guard3893 = fsm_out == 1'd0;
wire _guard3894 = cond_wire334_out;
wire _guard3895 = _guard3893 & _guard3894;
wire _guard3896 = fsm_out == 1'd0;
wire _guard3897 = _guard3895 & _guard3896;
wire _guard3898 = _guard3892 | _guard3897;
wire _guard3899 = fsm_out == 1'd0;
wire _guard3900 = cond_wire338_out;
wire _guard3901 = _guard3899 & _guard3900;
wire _guard3902 = fsm_out == 1'd0;
wire _guard3903 = _guard3901 & _guard3902;
wire _guard3904 = _guard3898 | _guard3903;
wire _guard3905 = early_reset_static_par0_go_out;
wire _guard3906 = _guard3904 & _guard3905;
wire _guard3907 = cond_wire_out;
wire _guard3908 = early_reset_static_par0_go_out;
wire _guard3909 = _guard3907 & _guard3908;
wire _guard3910 = cond_wire4_out;
wire _guard3911 = early_reset_static_par0_go_out;
wire _guard3912 = _guard3910 & _guard3911;
wire _guard3913 = cond_wire54_out;
wire _guard3914 = early_reset_static_par0_go_out;
wire _guard3915 = _guard3913 & _guard3914;
wire _guard3916 = fsm_out == 1'd0;
wire _guard3917 = cond_wire3_out;
wire _guard3918 = _guard3916 & _guard3917;
wire _guard3919 = fsm_out == 1'd0;
wire _guard3920 = _guard3918 & _guard3919;
wire _guard3921 = fsm_out == 1'd0;
wire _guard3922 = cond_wire8_out;
wire _guard3923 = _guard3921 & _guard3922;
wire _guard3924 = fsm_out == 1'd0;
wire _guard3925 = _guard3923 & _guard3924;
wire _guard3926 = _guard3920 | _guard3925;
wire _guard3927 = fsm_out == 1'd0;
wire _guard3928 = cond_wire13_out;
wire _guard3929 = _guard3927 & _guard3928;
wire _guard3930 = fsm_out == 1'd0;
wire _guard3931 = _guard3929 & _guard3930;
wire _guard3932 = _guard3926 | _guard3931;
wire _guard3933 = fsm_out == 1'd0;
wire _guard3934 = cond_wire18_out;
wire _guard3935 = _guard3933 & _guard3934;
wire _guard3936 = fsm_out == 1'd0;
wire _guard3937 = _guard3935 & _guard3936;
wire _guard3938 = _guard3932 | _guard3937;
wire _guard3939 = fsm_out == 1'd0;
wire _guard3940 = cond_wire23_out;
wire _guard3941 = _guard3939 & _guard3940;
wire _guard3942 = fsm_out == 1'd0;
wire _guard3943 = _guard3941 & _guard3942;
wire _guard3944 = _guard3938 | _guard3943;
wire _guard3945 = fsm_out == 1'd0;
wire _guard3946 = cond_wire28_out;
wire _guard3947 = _guard3945 & _guard3946;
wire _guard3948 = fsm_out == 1'd0;
wire _guard3949 = _guard3947 & _guard3948;
wire _guard3950 = _guard3944 | _guard3949;
wire _guard3951 = fsm_out == 1'd0;
wire _guard3952 = cond_wire33_out;
wire _guard3953 = _guard3951 & _guard3952;
wire _guard3954 = fsm_out == 1'd0;
wire _guard3955 = _guard3953 & _guard3954;
wire _guard3956 = _guard3950 | _guard3955;
wire _guard3957 = fsm_out == 1'd0;
wire _guard3958 = cond_wire38_out;
wire _guard3959 = _guard3957 & _guard3958;
wire _guard3960 = fsm_out == 1'd0;
wire _guard3961 = _guard3959 & _guard3960;
wire _guard3962 = _guard3956 | _guard3961;
wire _guard3963 = fsm_out == 1'd0;
wire _guard3964 = cond_wire43_out;
wire _guard3965 = _guard3963 & _guard3964;
wire _guard3966 = fsm_out == 1'd0;
wire _guard3967 = _guard3965 & _guard3966;
wire _guard3968 = _guard3962 | _guard3967;
wire _guard3969 = fsm_out == 1'd0;
wire _guard3970 = cond_wire48_out;
wire _guard3971 = _guard3969 & _guard3970;
wire _guard3972 = fsm_out == 1'd0;
wire _guard3973 = _guard3971 & _guard3972;
wire _guard3974 = _guard3968 | _guard3973;
wire _guard3975 = fsm_out == 1'd0;
wire _guard3976 = cond_wire53_out;
wire _guard3977 = _guard3975 & _guard3976;
wire _guard3978 = fsm_out == 1'd0;
wire _guard3979 = _guard3977 & _guard3978;
wire _guard3980 = _guard3974 | _guard3979;
wire _guard3981 = fsm_out == 1'd0;
wire _guard3982 = cond_wire58_out;
wire _guard3983 = _guard3981 & _guard3982;
wire _guard3984 = fsm_out == 1'd0;
wire _guard3985 = _guard3983 & _guard3984;
wire _guard3986 = _guard3980 | _guard3985;
wire _guard3987 = fsm_out == 1'd0;
wire _guard3988 = cond_wire63_out;
wire _guard3989 = _guard3987 & _guard3988;
wire _guard3990 = fsm_out == 1'd0;
wire _guard3991 = _guard3989 & _guard3990;
wire _guard3992 = _guard3986 | _guard3991;
wire _guard3993 = fsm_out == 1'd0;
wire _guard3994 = cond_wire68_out;
wire _guard3995 = _guard3993 & _guard3994;
wire _guard3996 = fsm_out == 1'd0;
wire _guard3997 = _guard3995 & _guard3996;
wire _guard3998 = _guard3992 | _guard3997;
wire _guard3999 = fsm_out == 1'd0;
wire _guard4000 = cond_wire73_out;
wire _guard4001 = _guard3999 & _guard4000;
wire _guard4002 = fsm_out == 1'd0;
wire _guard4003 = _guard4001 & _guard4002;
wire _guard4004 = _guard3998 | _guard4003;
wire _guard4005 = fsm_out == 1'd0;
wire _guard4006 = cond_wire78_out;
wire _guard4007 = _guard4005 & _guard4006;
wire _guard4008 = fsm_out == 1'd0;
wire _guard4009 = _guard4007 & _guard4008;
wire _guard4010 = _guard4004 | _guard4009;
wire _guard4011 = early_reset_static_par0_go_out;
wire _guard4012 = _guard4010 & _guard4011;
wire _guard4013 = fsm_out == 1'd0;
wire _guard4014 = cond_wire148_out;
wire _guard4015 = _guard4013 & _guard4014;
wire _guard4016 = fsm_out == 1'd0;
wire _guard4017 = _guard4015 & _guard4016;
wire _guard4018 = fsm_out == 1'd0;
wire _guard4019 = cond_wire152_out;
wire _guard4020 = _guard4018 & _guard4019;
wire _guard4021 = fsm_out == 1'd0;
wire _guard4022 = _guard4020 & _guard4021;
wire _guard4023 = _guard4017 | _guard4022;
wire _guard4024 = fsm_out == 1'd0;
wire _guard4025 = cond_wire156_out;
wire _guard4026 = _guard4024 & _guard4025;
wire _guard4027 = fsm_out == 1'd0;
wire _guard4028 = _guard4026 & _guard4027;
wire _guard4029 = _guard4023 | _guard4028;
wire _guard4030 = fsm_out == 1'd0;
wire _guard4031 = cond_wire160_out;
wire _guard4032 = _guard4030 & _guard4031;
wire _guard4033 = fsm_out == 1'd0;
wire _guard4034 = _guard4032 & _guard4033;
wire _guard4035 = _guard4029 | _guard4034;
wire _guard4036 = fsm_out == 1'd0;
wire _guard4037 = cond_wire164_out;
wire _guard4038 = _guard4036 & _guard4037;
wire _guard4039 = fsm_out == 1'd0;
wire _guard4040 = _guard4038 & _guard4039;
wire _guard4041 = _guard4035 | _guard4040;
wire _guard4042 = fsm_out == 1'd0;
wire _guard4043 = cond_wire168_out;
wire _guard4044 = _guard4042 & _guard4043;
wire _guard4045 = fsm_out == 1'd0;
wire _guard4046 = _guard4044 & _guard4045;
wire _guard4047 = _guard4041 | _guard4046;
wire _guard4048 = fsm_out == 1'd0;
wire _guard4049 = cond_wire172_out;
wire _guard4050 = _guard4048 & _guard4049;
wire _guard4051 = fsm_out == 1'd0;
wire _guard4052 = _guard4050 & _guard4051;
wire _guard4053 = _guard4047 | _guard4052;
wire _guard4054 = fsm_out == 1'd0;
wire _guard4055 = cond_wire176_out;
wire _guard4056 = _guard4054 & _guard4055;
wire _guard4057 = fsm_out == 1'd0;
wire _guard4058 = _guard4056 & _guard4057;
wire _guard4059 = _guard4053 | _guard4058;
wire _guard4060 = fsm_out == 1'd0;
wire _guard4061 = cond_wire180_out;
wire _guard4062 = _guard4060 & _guard4061;
wire _guard4063 = fsm_out == 1'd0;
wire _guard4064 = _guard4062 & _guard4063;
wire _guard4065 = _guard4059 | _guard4064;
wire _guard4066 = fsm_out == 1'd0;
wire _guard4067 = cond_wire184_out;
wire _guard4068 = _guard4066 & _guard4067;
wire _guard4069 = fsm_out == 1'd0;
wire _guard4070 = _guard4068 & _guard4069;
wire _guard4071 = _guard4065 | _guard4070;
wire _guard4072 = fsm_out == 1'd0;
wire _guard4073 = cond_wire188_out;
wire _guard4074 = _guard4072 & _guard4073;
wire _guard4075 = fsm_out == 1'd0;
wire _guard4076 = _guard4074 & _guard4075;
wire _guard4077 = _guard4071 | _guard4076;
wire _guard4078 = fsm_out == 1'd0;
wire _guard4079 = cond_wire192_out;
wire _guard4080 = _guard4078 & _guard4079;
wire _guard4081 = fsm_out == 1'd0;
wire _guard4082 = _guard4080 & _guard4081;
wire _guard4083 = _guard4077 | _guard4082;
wire _guard4084 = fsm_out == 1'd0;
wire _guard4085 = cond_wire196_out;
wire _guard4086 = _guard4084 & _guard4085;
wire _guard4087 = fsm_out == 1'd0;
wire _guard4088 = _guard4086 & _guard4087;
wire _guard4089 = _guard4083 | _guard4088;
wire _guard4090 = fsm_out == 1'd0;
wire _guard4091 = cond_wire200_out;
wire _guard4092 = _guard4090 & _guard4091;
wire _guard4093 = fsm_out == 1'd0;
wire _guard4094 = _guard4092 & _guard4093;
wire _guard4095 = _guard4089 | _guard4094;
wire _guard4096 = fsm_out == 1'd0;
wire _guard4097 = cond_wire204_out;
wire _guard4098 = _guard4096 & _guard4097;
wire _guard4099 = fsm_out == 1'd0;
wire _guard4100 = _guard4098 & _guard4099;
wire _guard4101 = _guard4095 | _guard4100;
wire _guard4102 = fsm_out == 1'd0;
wire _guard4103 = cond_wire208_out;
wire _guard4104 = _guard4102 & _guard4103;
wire _guard4105 = fsm_out == 1'd0;
wire _guard4106 = _guard4104 & _guard4105;
wire _guard4107 = _guard4101 | _guard4106;
wire _guard4108 = early_reset_static_par0_go_out;
wire _guard4109 = _guard4107 & _guard4108;
wire _guard4110 = cond_wire534_out;
wire _guard4111 = early_reset_static_par0_go_out;
wire _guard4112 = _guard4110 & _guard4111;
wire _guard4113 = fsm_out == 1'd0;
wire _guard4114 = cond_wire213_out;
wire _guard4115 = _guard4113 & _guard4114;
wire _guard4116 = fsm_out == 1'd0;
wire _guard4117 = _guard4115 & _guard4116;
wire _guard4118 = fsm_out == 1'd0;
wire _guard4119 = cond_wire217_out;
wire _guard4120 = _guard4118 & _guard4119;
wire _guard4121 = fsm_out == 1'd0;
wire _guard4122 = _guard4120 & _guard4121;
wire _guard4123 = _guard4117 | _guard4122;
wire _guard4124 = fsm_out == 1'd0;
wire _guard4125 = cond_wire221_out;
wire _guard4126 = _guard4124 & _guard4125;
wire _guard4127 = fsm_out == 1'd0;
wire _guard4128 = _guard4126 & _guard4127;
wire _guard4129 = _guard4123 | _guard4128;
wire _guard4130 = fsm_out == 1'd0;
wire _guard4131 = cond_wire225_out;
wire _guard4132 = _guard4130 & _guard4131;
wire _guard4133 = fsm_out == 1'd0;
wire _guard4134 = _guard4132 & _guard4133;
wire _guard4135 = _guard4129 | _guard4134;
wire _guard4136 = fsm_out == 1'd0;
wire _guard4137 = cond_wire229_out;
wire _guard4138 = _guard4136 & _guard4137;
wire _guard4139 = fsm_out == 1'd0;
wire _guard4140 = _guard4138 & _guard4139;
wire _guard4141 = _guard4135 | _guard4140;
wire _guard4142 = fsm_out == 1'd0;
wire _guard4143 = cond_wire233_out;
wire _guard4144 = _guard4142 & _guard4143;
wire _guard4145 = fsm_out == 1'd0;
wire _guard4146 = _guard4144 & _guard4145;
wire _guard4147 = _guard4141 | _guard4146;
wire _guard4148 = fsm_out == 1'd0;
wire _guard4149 = cond_wire237_out;
wire _guard4150 = _guard4148 & _guard4149;
wire _guard4151 = fsm_out == 1'd0;
wire _guard4152 = _guard4150 & _guard4151;
wire _guard4153 = _guard4147 | _guard4152;
wire _guard4154 = fsm_out == 1'd0;
wire _guard4155 = cond_wire241_out;
wire _guard4156 = _guard4154 & _guard4155;
wire _guard4157 = fsm_out == 1'd0;
wire _guard4158 = _guard4156 & _guard4157;
wire _guard4159 = _guard4153 | _guard4158;
wire _guard4160 = fsm_out == 1'd0;
wire _guard4161 = cond_wire245_out;
wire _guard4162 = _guard4160 & _guard4161;
wire _guard4163 = fsm_out == 1'd0;
wire _guard4164 = _guard4162 & _guard4163;
wire _guard4165 = _guard4159 | _guard4164;
wire _guard4166 = fsm_out == 1'd0;
wire _guard4167 = cond_wire249_out;
wire _guard4168 = _guard4166 & _guard4167;
wire _guard4169 = fsm_out == 1'd0;
wire _guard4170 = _guard4168 & _guard4169;
wire _guard4171 = _guard4165 | _guard4170;
wire _guard4172 = fsm_out == 1'd0;
wire _guard4173 = cond_wire253_out;
wire _guard4174 = _guard4172 & _guard4173;
wire _guard4175 = fsm_out == 1'd0;
wire _guard4176 = _guard4174 & _guard4175;
wire _guard4177 = _guard4171 | _guard4176;
wire _guard4178 = fsm_out == 1'd0;
wire _guard4179 = cond_wire257_out;
wire _guard4180 = _guard4178 & _guard4179;
wire _guard4181 = fsm_out == 1'd0;
wire _guard4182 = _guard4180 & _guard4181;
wire _guard4183 = _guard4177 | _guard4182;
wire _guard4184 = fsm_out == 1'd0;
wire _guard4185 = cond_wire261_out;
wire _guard4186 = _guard4184 & _guard4185;
wire _guard4187 = fsm_out == 1'd0;
wire _guard4188 = _guard4186 & _guard4187;
wire _guard4189 = _guard4183 | _guard4188;
wire _guard4190 = fsm_out == 1'd0;
wire _guard4191 = cond_wire265_out;
wire _guard4192 = _guard4190 & _guard4191;
wire _guard4193 = fsm_out == 1'd0;
wire _guard4194 = _guard4192 & _guard4193;
wire _guard4195 = _guard4189 | _guard4194;
wire _guard4196 = fsm_out == 1'd0;
wire _guard4197 = cond_wire269_out;
wire _guard4198 = _guard4196 & _guard4197;
wire _guard4199 = fsm_out == 1'd0;
wire _guard4200 = _guard4198 & _guard4199;
wire _guard4201 = _guard4195 | _guard4200;
wire _guard4202 = fsm_out == 1'd0;
wire _guard4203 = cond_wire273_out;
wire _guard4204 = _guard4202 & _guard4203;
wire _guard4205 = fsm_out == 1'd0;
wire _guard4206 = _guard4204 & _guard4205;
wire _guard4207 = _guard4201 | _guard4206;
wire _guard4208 = early_reset_static_par0_go_out;
wire _guard4209 = _guard4207 & _guard4208;
wire _guard4210 = cond_wire424_out;
wire _guard4211 = early_reset_static_par0_go_out;
wire _guard4212 = _guard4210 & _guard4211;
wire _guard4213 = cond_wire452_out;
wire _guard4214 = early_reset_static_par0_go_out;
wire _guard4215 = _guard4213 & _guard4214;
wire _guard4216 = cond_wire408_out;
wire _guard4217 = early_reset_static_par0_go_out;
wire _guard4218 = _guard4216 & _guard4217;
wire _guard4219 = cond_wire412_out;
wire _guard4220 = early_reset_static_par0_go_out;
wire _guard4221 = _guard4219 & _guard4220;
wire _guard4222 = cond_wire428_out;
wire _guard4223 = early_reset_static_par0_go_out;
wire _guard4224 = _guard4222 & _guard4223;
wire _guard4225 = cond_wire456_out;
wire _guard4226 = early_reset_static_par0_go_out;
wire _guard4227 = _guard4225 & _guard4226;
wire _guard4228 = cond_wire416_out;
wire _guard4229 = early_reset_static_par0_go_out;
wire _guard4230 = _guard4228 & _guard4229;
wire _guard4231 = cond_wire420_out;
wire _guard4232 = early_reset_static_par0_go_out;
wire _guard4233 = _guard4231 & _guard4232;
wire _guard4234 = cond_wire448_out;
wire _guard4235 = early_reset_static_par0_go_out;
wire _guard4236 = _guard4234 & _guard4235;
wire _guard4237 = cond_wire436_out;
wire _guard4238 = early_reset_static_par0_go_out;
wire _guard4239 = _guard4237 & _guard4238;
wire _guard4240 = cond_wire460_out;
wire _guard4241 = early_reset_static_par0_go_out;
wire _guard4242 = _guard4240 & _guard4241;
wire _guard4243 = cond_wire464_out;
wire _guard4244 = early_reset_static_par0_go_out;
wire _guard4245 = _guard4243 & _guard4244;
wire _guard4246 = cond_wire468_out;
wire _guard4247 = early_reset_static_par0_go_out;
wire _guard4248 = _guard4246 & _guard4247;
wire _guard4249 = cond_wire432_out;
wire _guard4250 = early_reset_static_par0_go_out;
wire _guard4251 = _guard4249 & _guard4250;
wire _guard4252 = cond_wire440_out;
wire _guard4253 = early_reset_static_par0_go_out;
wire _guard4254 = _guard4252 & _guard4253;
wire _guard4255 = cond_wire444_out;
wire _guard4256 = early_reset_static_par0_go_out;
wire _guard4257 = _guard4255 & _guard4256;
wire _guard4258 = fsm_out == 1'd0;
wire _guard4259 = cond_wire408_out;
wire _guard4260 = _guard4258 & _guard4259;
wire _guard4261 = fsm_out == 1'd0;
wire _guard4262 = _guard4260 & _guard4261;
wire _guard4263 = fsm_out == 1'd0;
wire _guard4264 = cond_wire412_out;
wire _guard4265 = _guard4263 & _guard4264;
wire _guard4266 = fsm_out == 1'd0;
wire _guard4267 = _guard4265 & _guard4266;
wire _guard4268 = _guard4262 | _guard4267;
wire _guard4269 = fsm_out == 1'd0;
wire _guard4270 = cond_wire416_out;
wire _guard4271 = _guard4269 & _guard4270;
wire _guard4272 = fsm_out == 1'd0;
wire _guard4273 = _guard4271 & _guard4272;
wire _guard4274 = _guard4268 | _guard4273;
wire _guard4275 = fsm_out == 1'd0;
wire _guard4276 = cond_wire420_out;
wire _guard4277 = _guard4275 & _guard4276;
wire _guard4278 = fsm_out == 1'd0;
wire _guard4279 = _guard4277 & _guard4278;
wire _guard4280 = _guard4274 | _guard4279;
wire _guard4281 = fsm_out == 1'd0;
wire _guard4282 = cond_wire424_out;
wire _guard4283 = _guard4281 & _guard4282;
wire _guard4284 = fsm_out == 1'd0;
wire _guard4285 = _guard4283 & _guard4284;
wire _guard4286 = _guard4280 | _guard4285;
wire _guard4287 = fsm_out == 1'd0;
wire _guard4288 = cond_wire428_out;
wire _guard4289 = _guard4287 & _guard4288;
wire _guard4290 = fsm_out == 1'd0;
wire _guard4291 = _guard4289 & _guard4290;
wire _guard4292 = _guard4286 | _guard4291;
wire _guard4293 = fsm_out == 1'd0;
wire _guard4294 = cond_wire432_out;
wire _guard4295 = _guard4293 & _guard4294;
wire _guard4296 = fsm_out == 1'd0;
wire _guard4297 = _guard4295 & _guard4296;
wire _guard4298 = _guard4292 | _guard4297;
wire _guard4299 = fsm_out == 1'd0;
wire _guard4300 = cond_wire436_out;
wire _guard4301 = _guard4299 & _guard4300;
wire _guard4302 = fsm_out == 1'd0;
wire _guard4303 = _guard4301 & _guard4302;
wire _guard4304 = _guard4298 | _guard4303;
wire _guard4305 = fsm_out == 1'd0;
wire _guard4306 = cond_wire440_out;
wire _guard4307 = _guard4305 & _guard4306;
wire _guard4308 = fsm_out == 1'd0;
wire _guard4309 = _guard4307 & _guard4308;
wire _guard4310 = _guard4304 | _guard4309;
wire _guard4311 = fsm_out == 1'd0;
wire _guard4312 = cond_wire444_out;
wire _guard4313 = _guard4311 & _guard4312;
wire _guard4314 = fsm_out == 1'd0;
wire _guard4315 = _guard4313 & _guard4314;
wire _guard4316 = _guard4310 | _guard4315;
wire _guard4317 = fsm_out == 1'd0;
wire _guard4318 = cond_wire448_out;
wire _guard4319 = _guard4317 & _guard4318;
wire _guard4320 = fsm_out == 1'd0;
wire _guard4321 = _guard4319 & _guard4320;
wire _guard4322 = _guard4316 | _guard4321;
wire _guard4323 = fsm_out == 1'd0;
wire _guard4324 = cond_wire452_out;
wire _guard4325 = _guard4323 & _guard4324;
wire _guard4326 = fsm_out == 1'd0;
wire _guard4327 = _guard4325 & _guard4326;
wire _guard4328 = _guard4322 | _guard4327;
wire _guard4329 = fsm_out == 1'd0;
wire _guard4330 = cond_wire456_out;
wire _guard4331 = _guard4329 & _guard4330;
wire _guard4332 = fsm_out == 1'd0;
wire _guard4333 = _guard4331 & _guard4332;
wire _guard4334 = _guard4328 | _guard4333;
wire _guard4335 = fsm_out == 1'd0;
wire _guard4336 = cond_wire460_out;
wire _guard4337 = _guard4335 & _guard4336;
wire _guard4338 = fsm_out == 1'd0;
wire _guard4339 = _guard4337 & _guard4338;
wire _guard4340 = _guard4334 | _guard4339;
wire _guard4341 = fsm_out == 1'd0;
wire _guard4342 = cond_wire464_out;
wire _guard4343 = _guard4341 & _guard4342;
wire _guard4344 = fsm_out == 1'd0;
wire _guard4345 = _guard4343 & _guard4344;
wire _guard4346 = _guard4340 | _guard4345;
wire _guard4347 = fsm_out == 1'd0;
wire _guard4348 = cond_wire468_out;
wire _guard4349 = _guard4347 & _guard4348;
wire _guard4350 = fsm_out == 1'd0;
wire _guard4351 = _guard4349 & _guard4350;
wire _guard4352 = _guard4346 | _guard4351;
wire _guard4353 = early_reset_static_par0_go_out;
wire _guard4354 = _guard4352 & _guard4353;
wire _guard4355 = cond_wire509_out;
wire _guard4356 = early_reset_static_par0_go_out;
wire _guard4357 = _guard4355 & _guard4356;
wire _guard4358 = cond_wire485_out;
wire _guard4359 = early_reset_static_par0_go_out;
wire _guard4360 = _guard4358 & _guard4359;
wire _guard4361 = cond_wire533_out;
wire _guard4362 = early_reset_static_par0_go_out;
wire _guard4363 = _guard4361 & _guard4362;
wire _guard4364 = cond_wire489_out;
wire _guard4365 = early_reset_static_par0_go_out;
wire _guard4366 = _guard4364 & _guard4365;
wire _guard4367 = cond_wire473_out;
wire _guard4368 = early_reset_static_par0_go_out;
wire _guard4369 = _guard4367 & _guard4368;
wire _guard4370 = cond_wire513_out;
wire _guard4371 = early_reset_static_par0_go_out;
wire _guard4372 = _guard4370 & _guard4371;
wire _guard4373 = cond_wire493_out;
wire _guard4374 = early_reset_static_par0_go_out;
wire _guard4375 = _guard4373 & _guard4374;
wire _guard4376 = cond_wire497_out;
wire _guard4377 = early_reset_static_par0_go_out;
wire _guard4378 = _guard4376 & _guard4377;
wire _guard4379 = cond_wire529_out;
wire _guard4380 = early_reset_static_par0_go_out;
wire _guard4381 = _guard4379 & _guard4380;
wire _guard4382 = cond_wire477_out;
wire _guard4383 = early_reset_static_par0_go_out;
wire _guard4384 = _guard4382 & _guard4383;
wire _guard4385 = cond_wire521_out;
wire _guard4386 = early_reset_static_par0_go_out;
wire _guard4387 = _guard4385 & _guard4386;
wire _guard4388 = cond_wire481_out;
wire _guard4389 = early_reset_static_par0_go_out;
wire _guard4390 = _guard4388 & _guard4389;
wire _guard4391 = cond_wire501_out;
wire _guard4392 = early_reset_static_par0_go_out;
wire _guard4393 = _guard4391 & _guard4392;
wire _guard4394 = cond_wire505_out;
wire _guard4395 = early_reset_static_par0_go_out;
wire _guard4396 = _guard4394 & _guard4395;
wire _guard4397 = cond_wire517_out;
wire _guard4398 = early_reset_static_par0_go_out;
wire _guard4399 = _guard4397 & _guard4398;
wire _guard4400 = cond_wire525_out;
wire _guard4401 = early_reset_static_par0_go_out;
wire _guard4402 = _guard4400 & _guard4401;
wire _guard4403 = fsm_out == 1'd0;
wire _guard4404 = cond_wire668_out;
wire _guard4405 = _guard4403 & _guard4404;
wire _guard4406 = fsm_out == 1'd0;
wire _guard4407 = _guard4405 & _guard4406;
wire _guard4408 = fsm_out == 1'd0;
wire _guard4409 = cond_wire672_out;
wire _guard4410 = _guard4408 & _guard4409;
wire _guard4411 = fsm_out == 1'd0;
wire _guard4412 = _guard4410 & _guard4411;
wire _guard4413 = _guard4407 | _guard4412;
wire _guard4414 = fsm_out == 1'd0;
wire _guard4415 = cond_wire676_out;
wire _guard4416 = _guard4414 & _guard4415;
wire _guard4417 = fsm_out == 1'd0;
wire _guard4418 = _guard4416 & _guard4417;
wire _guard4419 = _guard4413 | _guard4418;
wire _guard4420 = fsm_out == 1'd0;
wire _guard4421 = cond_wire680_out;
wire _guard4422 = _guard4420 & _guard4421;
wire _guard4423 = fsm_out == 1'd0;
wire _guard4424 = _guard4422 & _guard4423;
wire _guard4425 = _guard4419 | _guard4424;
wire _guard4426 = fsm_out == 1'd0;
wire _guard4427 = cond_wire684_out;
wire _guard4428 = _guard4426 & _guard4427;
wire _guard4429 = fsm_out == 1'd0;
wire _guard4430 = _guard4428 & _guard4429;
wire _guard4431 = _guard4425 | _guard4430;
wire _guard4432 = fsm_out == 1'd0;
wire _guard4433 = cond_wire688_out;
wire _guard4434 = _guard4432 & _guard4433;
wire _guard4435 = fsm_out == 1'd0;
wire _guard4436 = _guard4434 & _guard4435;
wire _guard4437 = _guard4431 | _guard4436;
wire _guard4438 = fsm_out == 1'd0;
wire _guard4439 = cond_wire692_out;
wire _guard4440 = _guard4438 & _guard4439;
wire _guard4441 = fsm_out == 1'd0;
wire _guard4442 = _guard4440 & _guard4441;
wire _guard4443 = _guard4437 | _guard4442;
wire _guard4444 = fsm_out == 1'd0;
wire _guard4445 = cond_wire696_out;
wire _guard4446 = _guard4444 & _guard4445;
wire _guard4447 = fsm_out == 1'd0;
wire _guard4448 = _guard4446 & _guard4447;
wire _guard4449 = _guard4443 | _guard4448;
wire _guard4450 = fsm_out == 1'd0;
wire _guard4451 = cond_wire700_out;
wire _guard4452 = _guard4450 & _guard4451;
wire _guard4453 = fsm_out == 1'd0;
wire _guard4454 = _guard4452 & _guard4453;
wire _guard4455 = _guard4449 | _guard4454;
wire _guard4456 = fsm_out == 1'd0;
wire _guard4457 = cond_wire704_out;
wire _guard4458 = _guard4456 & _guard4457;
wire _guard4459 = fsm_out == 1'd0;
wire _guard4460 = _guard4458 & _guard4459;
wire _guard4461 = _guard4455 | _guard4460;
wire _guard4462 = fsm_out == 1'd0;
wire _guard4463 = cond_wire708_out;
wire _guard4464 = _guard4462 & _guard4463;
wire _guard4465 = fsm_out == 1'd0;
wire _guard4466 = _guard4464 & _guard4465;
wire _guard4467 = _guard4461 | _guard4466;
wire _guard4468 = fsm_out == 1'd0;
wire _guard4469 = cond_wire712_out;
wire _guard4470 = _guard4468 & _guard4469;
wire _guard4471 = fsm_out == 1'd0;
wire _guard4472 = _guard4470 & _guard4471;
wire _guard4473 = _guard4467 | _guard4472;
wire _guard4474 = fsm_out == 1'd0;
wire _guard4475 = cond_wire716_out;
wire _guard4476 = _guard4474 & _guard4475;
wire _guard4477 = fsm_out == 1'd0;
wire _guard4478 = _guard4476 & _guard4477;
wire _guard4479 = _guard4473 | _guard4478;
wire _guard4480 = fsm_out == 1'd0;
wire _guard4481 = cond_wire720_out;
wire _guard4482 = _guard4480 & _guard4481;
wire _guard4483 = fsm_out == 1'd0;
wire _guard4484 = _guard4482 & _guard4483;
wire _guard4485 = _guard4479 | _guard4484;
wire _guard4486 = fsm_out == 1'd0;
wire _guard4487 = cond_wire724_out;
wire _guard4488 = _guard4486 & _guard4487;
wire _guard4489 = fsm_out == 1'd0;
wire _guard4490 = _guard4488 & _guard4489;
wire _guard4491 = _guard4485 | _guard4490;
wire _guard4492 = fsm_out == 1'd0;
wire _guard4493 = cond_wire728_out;
wire _guard4494 = _guard4492 & _guard4493;
wire _guard4495 = fsm_out == 1'd0;
wire _guard4496 = _guard4494 & _guard4495;
wire _guard4497 = _guard4491 | _guard4496;
wire _guard4498 = early_reset_static_par0_go_out;
wire _guard4499 = _guard4497 & _guard4498;
wire _guard4500 = fsm_out == 1'd0;
wire _guard4501 = cond_wire928_out;
wire _guard4502 = _guard4500 & _guard4501;
wire _guard4503 = fsm_out == 1'd0;
wire _guard4504 = _guard4502 & _guard4503;
wire _guard4505 = fsm_out == 1'd0;
wire _guard4506 = cond_wire932_out;
wire _guard4507 = _guard4505 & _guard4506;
wire _guard4508 = fsm_out == 1'd0;
wire _guard4509 = _guard4507 & _guard4508;
wire _guard4510 = _guard4504 | _guard4509;
wire _guard4511 = fsm_out == 1'd0;
wire _guard4512 = cond_wire936_out;
wire _guard4513 = _guard4511 & _guard4512;
wire _guard4514 = fsm_out == 1'd0;
wire _guard4515 = _guard4513 & _guard4514;
wire _guard4516 = _guard4510 | _guard4515;
wire _guard4517 = fsm_out == 1'd0;
wire _guard4518 = cond_wire940_out;
wire _guard4519 = _guard4517 & _guard4518;
wire _guard4520 = fsm_out == 1'd0;
wire _guard4521 = _guard4519 & _guard4520;
wire _guard4522 = _guard4516 | _guard4521;
wire _guard4523 = fsm_out == 1'd0;
wire _guard4524 = cond_wire944_out;
wire _guard4525 = _guard4523 & _guard4524;
wire _guard4526 = fsm_out == 1'd0;
wire _guard4527 = _guard4525 & _guard4526;
wire _guard4528 = _guard4522 | _guard4527;
wire _guard4529 = fsm_out == 1'd0;
wire _guard4530 = cond_wire948_out;
wire _guard4531 = _guard4529 & _guard4530;
wire _guard4532 = fsm_out == 1'd0;
wire _guard4533 = _guard4531 & _guard4532;
wire _guard4534 = _guard4528 | _guard4533;
wire _guard4535 = fsm_out == 1'd0;
wire _guard4536 = cond_wire952_out;
wire _guard4537 = _guard4535 & _guard4536;
wire _guard4538 = fsm_out == 1'd0;
wire _guard4539 = _guard4537 & _guard4538;
wire _guard4540 = _guard4534 | _guard4539;
wire _guard4541 = fsm_out == 1'd0;
wire _guard4542 = cond_wire956_out;
wire _guard4543 = _guard4541 & _guard4542;
wire _guard4544 = fsm_out == 1'd0;
wire _guard4545 = _guard4543 & _guard4544;
wire _guard4546 = _guard4540 | _guard4545;
wire _guard4547 = fsm_out == 1'd0;
wire _guard4548 = cond_wire960_out;
wire _guard4549 = _guard4547 & _guard4548;
wire _guard4550 = fsm_out == 1'd0;
wire _guard4551 = _guard4549 & _guard4550;
wire _guard4552 = _guard4546 | _guard4551;
wire _guard4553 = fsm_out == 1'd0;
wire _guard4554 = cond_wire964_out;
wire _guard4555 = _guard4553 & _guard4554;
wire _guard4556 = fsm_out == 1'd0;
wire _guard4557 = _guard4555 & _guard4556;
wire _guard4558 = _guard4552 | _guard4557;
wire _guard4559 = fsm_out == 1'd0;
wire _guard4560 = cond_wire968_out;
wire _guard4561 = _guard4559 & _guard4560;
wire _guard4562 = fsm_out == 1'd0;
wire _guard4563 = _guard4561 & _guard4562;
wire _guard4564 = _guard4558 | _guard4563;
wire _guard4565 = fsm_out == 1'd0;
wire _guard4566 = cond_wire972_out;
wire _guard4567 = _guard4565 & _guard4566;
wire _guard4568 = fsm_out == 1'd0;
wire _guard4569 = _guard4567 & _guard4568;
wire _guard4570 = _guard4564 | _guard4569;
wire _guard4571 = fsm_out == 1'd0;
wire _guard4572 = cond_wire976_out;
wire _guard4573 = _guard4571 & _guard4572;
wire _guard4574 = fsm_out == 1'd0;
wire _guard4575 = _guard4573 & _guard4574;
wire _guard4576 = _guard4570 | _guard4575;
wire _guard4577 = fsm_out == 1'd0;
wire _guard4578 = cond_wire980_out;
wire _guard4579 = _guard4577 & _guard4578;
wire _guard4580 = fsm_out == 1'd0;
wire _guard4581 = _guard4579 & _guard4580;
wire _guard4582 = _guard4576 | _guard4581;
wire _guard4583 = fsm_out == 1'd0;
wire _guard4584 = cond_wire984_out;
wire _guard4585 = _guard4583 & _guard4584;
wire _guard4586 = fsm_out == 1'd0;
wire _guard4587 = _guard4585 & _guard4586;
wire _guard4588 = _guard4582 | _guard4587;
wire _guard4589 = fsm_out == 1'd0;
wire _guard4590 = cond_wire988_out;
wire _guard4591 = _guard4589 & _guard4590;
wire _guard4592 = fsm_out == 1'd0;
wire _guard4593 = _guard4591 & _guard4592;
wire _guard4594 = _guard4588 | _guard4593;
wire _guard4595 = early_reset_static_par0_go_out;
wire _guard4596 = _guard4594 & _guard4595;
wire _guard4597 = cond_wire49_out;
wire _guard4598 = early_reset_static_par0_go_out;
wire _guard4599 = _guard4597 & _guard4598;
wire _guard4600 = cond_wire144_out;
wire _guard4601 = early_reset_static_par0_go_out;
wire _guard4602 = _guard4600 & _guard4601;
wire _guard4603 = cond_wire599_out;
wire _guard4604 = early_reset_static_par0_go_out;
wire _guard4605 = _guard4603 & _guard4604;
wire _guard4606 = cond_wire794_out;
wire _guard4607 = early_reset_static_par0_go_out;
wire _guard4608 = _guard4606 & _guard4607;
wire _guard4609 = cond_wire8_out;
wire _guard4610 = early_reset_static_par0_go_out;
wire _guard4611 = _guard4609 & _guard4610;
wire _guard4612 = cond_wire78_out;
wire _guard4613 = early_reset_static_par0_go_out;
wire _guard4614 = _guard4612 & _guard4613;
wire _guard4615 = cond_wire3_out;
wire _guard4616 = early_reset_static_par0_go_out;
wire _guard4617 = _guard4615 & _guard4616;
wire _guard4618 = cond_wire18_out;
wire _guard4619 = early_reset_static_par0_go_out;
wire _guard4620 = _guard4618 & _guard4619;
wire _guard4621 = cond_wire68_out;
wire _guard4622 = early_reset_static_par0_go_out;
wire _guard4623 = _guard4621 & _guard4622;
wire _guard4624 = cond_wire73_out;
wire _guard4625 = early_reset_static_par0_go_out;
wire _guard4626 = _guard4624 & _guard4625;
wire _guard4627 = cond_wire28_out;
wire _guard4628 = early_reset_static_par0_go_out;
wire _guard4629 = _guard4627 & _guard4628;
wire _guard4630 = cond_wire63_out;
wire _guard4631 = early_reset_static_par0_go_out;
wire _guard4632 = _guard4630 & _guard4631;
wire _guard4633 = cond_wire13_out;
wire _guard4634 = early_reset_static_par0_go_out;
wire _guard4635 = _guard4633 & _guard4634;
wire _guard4636 = cond_wire43_out;
wire _guard4637 = early_reset_static_par0_go_out;
wire _guard4638 = _guard4636 & _guard4637;
wire _guard4639 = cond_wire53_out;
wire _guard4640 = early_reset_static_par0_go_out;
wire _guard4641 = _guard4639 & _guard4640;
wire _guard4642 = cond_wire38_out;
wire _guard4643 = early_reset_static_par0_go_out;
wire _guard4644 = _guard4642 & _guard4643;
wire _guard4645 = cond_wire58_out;
wire _guard4646 = early_reset_static_par0_go_out;
wire _guard4647 = _guard4645 & _guard4646;
wire _guard4648 = cond_wire23_out;
wire _guard4649 = early_reset_static_par0_go_out;
wire _guard4650 = _guard4648 & _guard4649;
wire _guard4651 = cond_wire33_out;
wire _guard4652 = early_reset_static_par0_go_out;
wire _guard4653 = _guard4651 & _guard4652;
wire _guard4654 = cond_wire48_out;
wire _guard4655 = early_reset_static_par0_go_out;
wire _guard4656 = _guard4654 & _guard4655;
wire _guard4657 = cond_wire217_out;
wire _guard4658 = early_reset_static_par0_go_out;
wire _guard4659 = _guard4657 & _guard4658;
wire _guard4660 = cond_wire273_out;
wire _guard4661 = early_reset_static_par0_go_out;
wire _guard4662 = _guard4660 & _guard4661;
wire _guard4663 = cond_wire213_out;
wire _guard4664 = early_reset_static_par0_go_out;
wire _guard4665 = _guard4663 & _guard4664;
wire _guard4666 = cond_wire225_out;
wire _guard4667 = early_reset_static_par0_go_out;
wire _guard4668 = _guard4666 & _guard4667;
wire _guard4669 = cond_wire265_out;
wire _guard4670 = early_reset_static_par0_go_out;
wire _guard4671 = _guard4669 & _guard4670;
wire _guard4672 = cond_wire269_out;
wire _guard4673 = early_reset_static_par0_go_out;
wire _guard4674 = _guard4672 & _guard4673;
wire _guard4675 = cond_wire233_out;
wire _guard4676 = early_reset_static_par0_go_out;
wire _guard4677 = _guard4675 & _guard4676;
wire _guard4678 = cond_wire261_out;
wire _guard4679 = early_reset_static_par0_go_out;
wire _guard4680 = _guard4678 & _guard4679;
wire _guard4681 = cond_wire221_out;
wire _guard4682 = early_reset_static_par0_go_out;
wire _guard4683 = _guard4681 & _guard4682;
wire _guard4684 = cond_wire245_out;
wire _guard4685 = early_reset_static_par0_go_out;
wire _guard4686 = _guard4684 & _guard4685;
wire _guard4687 = cond_wire253_out;
wire _guard4688 = early_reset_static_par0_go_out;
wire _guard4689 = _guard4687 & _guard4688;
wire _guard4690 = cond_wire241_out;
wire _guard4691 = early_reset_static_par0_go_out;
wire _guard4692 = _guard4690 & _guard4691;
wire _guard4693 = cond_wire257_out;
wire _guard4694 = early_reset_static_par0_go_out;
wire _guard4695 = _guard4693 & _guard4694;
wire _guard4696 = cond_wire229_out;
wire _guard4697 = early_reset_static_par0_go_out;
wire _guard4698 = _guard4696 & _guard4697;
wire _guard4699 = cond_wire237_out;
wire _guard4700 = early_reset_static_par0_go_out;
wire _guard4701 = _guard4699 & _guard4700;
wire _guard4702 = cond_wire249_out;
wire _guard4703 = early_reset_static_par0_go_out;
wire _guard4704 = _guard4702 & _guard4703;
wire _guard4705 = cond_wire542_out;
wire _guard4706 = early_reset_static_par0_go_out;
wire _guard4707 = _guard4705 & _guard4706;
wire _guard4708 = cond_wire598_out;
wire _guard4709 = early_reset_static_par0_go_out;
wire _guard4710 = _guard4708 & _guard4709;
wire _guard4711 = cond_wire538_out;
wire _guard4712 = early_reset_static_par0_go_out;
wire _guard4713 = _guard4711 & _guard4712;
wire _guard4714 = cond_wire550_out;
wire _guard4715 = early_reset_static_par0_go_out;
wire _guard4716 = _guard4714 & _guard4715;
wire _guard4717 = cond_wire590_out;
wire _guard4718 = early_reset_static_par0_go_out;
wire _guard4719 = _guard4717 & _guard4718;
wire _guard4720 = cond_wire594_out;
wire _guard4721 = early_reset_static_par0_go_out;
wire _guard4722 = _guard4720 & _guard4721;
wire _guard4723 = cond_wire558_out;
wire _guard4724 = early_reset_static_par0_go_out;
wire _guard4725 = _guard4723 & _guard4724;
wire _guard4726 = cond_wire586_out;
wire _guard4727 = early_reset_static_par0_go_out;
wire _guard4728 = _guard4726 & _guard4727;
wire _guard4729 = cond_wire546_out;
wire _guard4730 = early_reset_static_par0_go_out;
wire _guard4731 = _guard4729 & _guard4730;
wire _guard4732 = cond_wire570_out;
wire _guard4733 = early_reset_static_par0_go_out;
wire _guard4734 = _guard4732 & _guard4733;
wire _guard4735 = cond_wire578_out;
wire _guard4736 = early_reset_static_par0_go_out;
wire _guard4737 = _guard4735 & _guard4736;
wire _guard4738 = cond_wire566_out;
wire _guard4739 = early_reset_static_par0_go_out;
wire _guard4740 = _guard4738 & _guard4739;
wire _guard4741 = cond_wire582_out;
wire _guard4742 = early_reset_static_par0_go_out;
wire _guard4743 = _guard4741 & _guard4742;
wire _guard4744 = cond_wire554_out;
wire _guard4745 = early_reset_static_par0_go_out;
wire _guard4746 = _guard4744 & _guard4745;
wire _guard4747 = cond_wire562_out;
wire _guard4748 = early_reset_static_par0_go_out;
wire _guard4749 = _guard4747 & _guard4748;
wire _guard4750 = cond_wire574_out;
wire _guard4751 = early_reset_static_par0_go_out;
wire _guard4752 = _guard4750 & _guard4751;
wire _guard4753 = cond_wire753_out;
wire _guard4754 = early_reset_static_par0_go_out;
wire _guard4755 = _guard4753 & _guard4754;
wire _guard4756 = cond_wire781_out;
wire _guard4757 = early_reset_static_par0_go_out;
wire _guard4758 = _guard4756 & _guard4757;
wire _guard4759 = cond_wire765_out;
wire _guard4760 = early_reset_static_par0_go_out;
wire _guard4761 = _guard4759 & _guard4760;
wire _guard4762 = cond_wire793_out;
wire _guard4763 = early_reset_static_par0_go_out;
wire _guard4764 = _guard4762 & _guard4763;
wire _guard4765 = cond_wire749_out;
wire _guard4766 = early_reset_static_par0_go_out;
wire _guard4767 = _guard4765 & _guard4766;
wire _guard4768 = cond_wire733_out;
wire _guard4769 = early_reset_static_par0_go_out;
wire _guard4770 = _guard4768 & _guard4769;
wire _guard4771 = cond_wire777_out;
wire _guard4772 = early_reset_static_par0_go_out;
wire _guard4773 = _guard4771 & _guard4772;
wire _guard4774 = cond_wire757_out;
wire _guard4775 = early_reset_static_par0_go_out;
wire _guard4776 = _guard4774 & _guard4775;
wire _guard4777 = cond_wire761_out;
wire _guard4778 = early_reset_static_par0_go_out;
wire _guard4779 = _guard4777 & _guard4778;
wire _guard4780 = cond_wire769_out;
wire _guard4781 = early_reset_static_par0_go_out;
wire _guard4782 = _guard4780 & _guard4781;
wire _guard4783 = cond_wire741_out;
wire _guard4784 = early_reset_static_par0_go_out;
wire _guard4785 = _guard4783 & _guard4784;
wire _guard4786 = cond_wire745_out;
wire _guard4787 = early_reset_static_par0_go_out;
wire _guard4788 = _guard4786 & _guard4787;
wire _guard4789 = cond_wire737_out;
wire _guard4790 = early_reset_static_par0_go_out;
wire _guard4791 = _guard4789 & _guard4790;
wire _guard4792 = cond_wire785_out;
wire _guard4793 = early_reset_static_par0_go_out;
wire _guard4794 = _guard4792 & _guard4793;
wire _guard4795 = cond_wire789_out;
wire _guard4796 = early_reset_static_par0_go_out;
wire _guard4797 = _guard4795 & _guard4796;
wire _guard4798 = cond_wire773_out;
wire _guard4799 = early_reset_static_par0_go_out;
wire _guard4800 = _guard4798 & _guard4799;
wire _guard4801 = cond_wire14_out;
wire _guard4802 = early_reset_static_par0_go_out;
wire _guard4803 = _guard4801 & _guard4802;
wire _guard4804 = cond_wire34_out;
wire _guard4805 = early_reset_static_par0_go_out;
wire _guard4806 = _guard4804 & _guard4805;
wire _guard4807 = cond_wire152_out;
wire _guard4808 = early_reset_static_par0_go_out;
wire _guard4809 = _guard4807 & _guard4808;
wire _guard4810 = cond_wire208_out;
wire _guard4811 = early_reset_static_par0_go_out;
wire _guard4812 = _guard4810 & _guard4811;
wire _guard4813 = cond_wire148_out;
wire _guard4814 = early_reset_static_par0_go_out;
wire _guard4815 = _guard4813 & _guard4814;
wire _guard4816 = cond_wire160_out;
wire _guard4817 = early_reset_static_par0_go_out;
wire _guard4818 = _guard4816 & _guard4817;
wire _guard4819 = cond_wire200_out;
wire _guard4820 = early_reset_static_par0_go_out;
wire _guard4821 = _guard4819 & _guard4820;
wire _guard4822 = cond_wire204_out;
wire _guard4823 = early_reset_static_par0_go_out;
wire _guard4824 = _guard4822 & _guard4823;
wire _guard4825 = cond_wire168_out;
wire _guard4826 = early_reset_static_par0_go_out;
wire _guard4827 = _guard4825 & _guard4826;
wire _guard4828 = cond_wire196_out;
wire _guard4829 = early_reset_static_par0_go_out;
wire _guard4830 = _guard4828 & _guard4829;
wire _guard4831 = cond_wire156_out;
wire _guard4832 = early_reset_static_par0_go_out;
wire _guard4833 = _guard4831 & _guard4832;
wire _guard4834 = cond_wire180_out;
wire _guard4835 = early_reset_static_par0_go_out;
wire _guard4836 = _guard4834 & _guard4835;
wire _guard4837 = cond_wire188_out;
wire _guard4838 = early_reset_static_par0_go_out;
wire _guard4839 = _guard4837 & _guard4838;
wire _guard4840 = cond_wire176_out;
wire _guard4841 = early_reset_static_par0_go_out;
wire _guard4842 = _guard4840 & _guard4841;
wire _guard4843 = cond_wire192_out;
wire _guard4844 = early_reset_static_par0_go_out;
wire _guard4845 = _guard4843 & _guard4844;
wire _guard4846 = cond_wire164_out;
wire _guard4847 = early_reset_static_par0_go_out;
wire _guard4848 = _guard4846 & _guard4847;
wire _guard4849 = cond_wire172_out;
wire _guard4850 = early_reset_static_par0_go_out;
wire _guard4851 = _guard4849 & _guard4850;
wire _guard4852 = cond_wire184_out;
wire _guard4853 = early_reset_static_par0_go_out;
wire _guard4854 = _guard4852 & _guard4853;
wire _guard4855 = cond_wire562_out;
wire _guard4856 = early_reset_static_par0_go_out;
wire _guard4857 = _guard4855 & _guard4856;
wire _guard4858 = cond_wire590_out;
wire _guard4859 = early_reset_static_par0_go_out;
wire _guard4860 = _guard4858 & _guard4859;
wire _guard4861 = cond_wire542_out;
wire _guard4862 = early_reset_static_par0_go_out;
wire _guard4863 = _guard4861 & _guard4862;
wire _guard4864 = cond_wire546_out;
wire _guard4865 = early_reset_static_par0_go_out;
wire _guard4866 = _guard4864 & _guard4865;
wire _guard4867 = cond_wire554_out;
wire _guard4868 = early_reset_static_par0_go_out;
wire _guard4869 = _guard4867 & _guard4868;
wire _guard4870 = cond_wire538_out;
wire _guard4871 = early_reset_static_par0_go_out;
wire _guard4872 = _guard4870 & _guard4871;
wire _guard4873 = cond_wire558_out;
wire _guard4874 = early_reset_static_par0_go_out;
wire _guard4875 = _guard4873 & _guard4874;
wire _guard4876 = cond_wire574_out;
wire _guard4877 = early_reset_static_par0_go_out;
wire _guard4878 = _guard4876 & _guard4877;
wire _guard4879 = cond_wire598_out;
wire _guard4880 = early_reset_static_par0_go_out;
wire _guard4881 = _guard4879 & _guard4880;
wire _guard4882 = cond_wire582_out;
wire _guard4883 = early_reset_static_par0_go_out;
wire _guard4884 = _guard4882 & _guard4883;
wire _guard4885 = cond_wire550_out;
wire _guard4886 = early_reset_static_par0_go_out;
wire _guard4887 = _guard4885 & _guard4886;
wire _guard4888 = cond_wire586_out;
wire _guard4889 = early_reset_static_par0_go_out;
wire _guard4890 = _guard4888 & _guard4889;
wire _guard4891 = cond_wire578_out;
wire _guard4892 = early_reset_static_par0_go_out;
wire _guard4893 = _guard4891 & _guard4892;
wire _guard4894 = cond_wire594_out;
wire _guard4895 = early_reset_static_par0_go_out;
wire _guard4896 = _guard4894 & _guard4895;
wire _guard4897 = cond_wire566_out;
wire _guard4898 = early_reset_static_par0_go_out;
wire _guard4899 = _guard4897 & _guard4898;
wire _guard4900 = cond_wire570_out;
wire _guard4901 = early_reset_static_par0_go_out;
wire _guard4902 = _guard4900 & _guard4901;
wire _guard4903 = fsm_out == 1'd0;
wire _guard4904 = cond_wire538_out;
wire _guard4905 = _guard4903 & _guard4904;
wire _guard4906 = fsm_out == 1'd0;
wire _guard4907 = _guard4905 & _guard4906;
wire _guard4908 = fsm_out == 1'd0;
wire _guard4909 = cond_wire542_out;
wire _guard4910 = _guard4908 & _guard4909;
wire _guard4911 = fsm_out == 1'd0;
wire _guard4912 = _guard4910 & _guard4911;
wire _guard4913 = _guard4907 | _guard4912;
wire _guard4914 = fsm_out == 1'd0;
wire _guard4915 = cond_wire546_out;
wire _guard4916 = _guard4914 & _guard4915;
wire _guard4917 = fsm_out == 1'd0;
wire _guard4918 = _guard4916 & _guard4917;
wire _guard4919 = _guard4913 | _guard4918;
wire _guard4920 = fsm_out == 1'd0;
wire _guard4921 = cond_wire550_out;
wire _guard4922 = _guard4920 & _guard4921;
wire _guard4923 = fsm_out == 1'd0;
wire _guard4924 = _guard4922 & _guard4923;
wire _guard4925 = _guard4919 | _guard4924;
wire _guard4926 = fsm_out == 1'd0;
wire _guard4927 = cond_wire554_out;
wire _guard4928 = _guard4926 & _guard4927;
wire _guard4929 = fsm_out == 1'd0;
wire _guard4930 = _guard4928 & _guard4929;
wire _guard4931 = _guard4925 | _guard4930;
wire _guard4932 = fsm_out == 1'd0;
wire _guard4933 = cond_wire558_out;
wire _guard4934 = _guard4932 & _guard4933;
wire _guard4935 = fsm_out == 1'd0;
wire _guard4936 = _guard4934 & _guard4935;
wire _guard4937 = _guard4931 | _guard4936;
wire _guard4938 = fsm_out == 1'd0;
wire _guard4939 = cond_wire562_out;
wire _guard4940 = _guard4938 & _guard4939;
wire _guard4941 = fsm_out == 1'd0;
wire _guard4942 = _guard4940 & _guard4941;
wire _guard4943 = _guard4937 | _guard4942;
wire _guard4944 = fsm_out == 1'd0;
wire _guard4945 = cond_wire566_out;
wire _guard4946 = _guard4944 & _guard4945;
wire _guard4947 = fsm_out == 1'd0;
wire _guard4948 = _guard4946 & _guard4947;
wire _guard4949 = _guard4943 | _guard4948;
wire _guard4950 = fsm_out == 1'd0;
wire _guard4951 = cond_wire570_out;
wire _guard4952 = _guard4950 & _guard4951;
wire _guard4953 = fsm_out == 1'd0;
wire _guard4954 = _guard4952 & _guard4953;
wire _guard4955 = _guard4949 | _guard4954;
wire _guard4956 = fsm_out == 1'd0;
wire _guard4957 = cond_wire574_out;
wire _guard4958 = _guard4956 & _guard4957;
wire _guard4959 = fsm_out == 1'd0;
wire _guard4960 = _guard4958 & _guard4959;
wire _guard4961 = _guard4955 | _guard4960;
wire _guard4962 = fsm_out == 1'd0;
wire _guard4963 = cond_wire578_out;
wire _guard4964 = _guard4962 & _guard4963;
wire _guard4965 = fsm_out == 1'd0;
wire _guard4966 = _guard4964 & _guard4965;
wire _guard4967 = _guard4961 | _guard4966;
wire _guard4968 = fsm_out == 1'd0;
wire _guard4969 = cond_wire582_out;
wire _guard4970 = _guard4968 & _guard4969;
wire _guard4971 = fsm_out == 1'd0;
wire _guard4972 = _guard4970 & _guard4971;
wire _guard4973 = _guard4967 | _guard4972;
wire _guard4974 = fsm_out == 1'd0;
wire _guard4975 = cond_wire586_out;
wire _guard4976 = _guard4974 & _guard4975;
wire _guard4977 = fsm_out == 1'd0;
wire _guard4978 = _guard4976 & _guard4977;
wire _guard4979 = _guard4973 | _guard4978;
wire _guard4980 = fsm_out == 1'd0;
wire _guard4981 = cond_wire590_out;
wire _guard4982 = _guard4980 & _guard4981;
wire _guard4983 = fsm_out == 1'd0;
wire _guard4984 = _guard4982 & _guard4983;
wire _guard4985 = _guard4979 | _guard4984;
wire _guard4986 = fsm_out == 1'd0;
wire _guard4987 = cond_wire594_out;
wire _guard4988 = _guard4986 & _guard4987;
wire _guard4989 = fsm_out == 1'd0;
wire _guard4990 = _guard4988 & _guard4989;
wire _guard4991 = _guard4985 | _guard4990;
wire _guard4992 = fsm_out == 1'd0;
wire _guard4993 = cond_wire598_out;
wire _guard4994 = _guard4992 & _guard4993;
wire _guard4995 = fsm_out == 1'd0;
wire _guard4996 = _guard4994 & _guard4995;
wire _guard4997 = _guard4991 | _guard4996;
wire _guard4998 = early_reset_static_par0_go_out;
wire _guard4999 = _guard4997 & _guard4998;
wire _guard5000 = cond_wire663_out;
wire _guard5001 = early_reset_static_par0_go_out;
wire _guard5002 = _guard5000 & _guard5001;
wire _guard5003 = cond_wire615_out;
wire _guard5004 = early_reset_static_par0_go_out;
wire _guard5005 = _guard5003 & _guard5004;
wire _guard5006 = cond_wire647_out;
wire _guard5007 = early_reset_static_par0_go_out;
wire _guard5008 = _guard5006 & _guard5007;
wire _guard5009 = cond_wire631_out;
wire _guard5010 = early_reset_static_par0_go_out;
wire _guard5011 = _guard5009 & _guard5010;
wire _guard5012 = cond_wire639_out;
wire _guard5013 = early_reset_static_par0_go_out;
wire _guard5014 = _guard5012 & _guard5013;
wire _guard5015 = cond_wire655_out;
wire _guard5016 = early_reset_static_par0_go_out;
wire _guard5017 = _guard5015 & _guard5016;
wire _guard5018 = cond_wire627_out;
wire _guard5019 = early_reset_static_par0_go_out;
wire _guard5020 = _guard5018 & _guard5019;
wire _guard5021 = cond_wire643_out;
wire _guard5022 = early_reset_static_par0_go_out;
wire _guard5023 = _guard5021 & _guard5022;
wire _guard5024 = cond_wire651_out;
wire _guard5025 = early_reset_static_par0_go_out;
wire _guard5026 = _guard5024 & _guard5025;
wire _guard5027 = cond_wire603_out;
wire _guard5028 = early_reset_static_par0_go_out;
wire _guard5029 = _guard5027 & _guard5028;
wire _guard5030 = cond_wire619_out;
wire _guard5031 = early_reset_static_par0_go_out;
wire _guard5032 = _guard5030 & _guard5031;
wire _guard5033 = cond_wire623_out;
wire _guard5034 = early_reset_static_par0_go_out;
wire _guard5035 = _guard5033 & _guard5034;
wire _guard5036 = cond_wire607_out;
wire _guard5037 = early_reset_static_par0_go_out;
wire _guard5038 = _guard5036 & _guard5037;
wire _guard5039 = cond_wire635_out;
wire _guard5040 = early_reset_static_par0_go_out;
wire _guard5041 = _guard5039 & _guard5040;
wire _guard5042 = cond_wire659_out;
wire _guard5043 = early_reset_static_par0_go_out;
wire _guard5044 = _guard5042 & _guard5043;
wire _guard5045 = cond_wire611_out;
wire _guard5046 = early_reset_static_par0_go_out;
wire _guard5047 = _guard5045 & _guard5046;
wire _guard5048 = cond_wire867_out;
wire _guard5049 = early_reset_static_par0_go_out;
wire _guard5050 = _guard5048 & _guard5049;
wire _guard5051 = cond_wire923_out;
wire _guard5052 = early_reset_static_par0_go_out;
wire _guard5053 = _guard5051 & _guard5052;
wire _guard5054 = cond_wire863_out;
wire _guard5055 = early_reset_static_par0_go_out;
wire _guard5056 = _guard5054 & _guard5055;
wire _guard5057 = cond_wire875_out;
wire _guard5058 = early_reset_static_par0_go_out;
wire _guard5059 = _guard5057 & _guard5058;
wire _guard5060 = cond_wire915_out;
wire _guard5061 = early_reset_static_par0_go_out;
wire _guard5062 = _guard5060 & _guard5061;
wire _guard5063 = cond_wire919_out;
wire _guard5064 = early_reset_static_par0_go_out;
wire _guard5065 = _guard5063 & _guard5064;
wire _guard5066 = cond_wire883_out;
wire _guard5067 = early_reset_static_par0_go_out;
wire _guard5068 = _guard5066 & _guard5067;
wire _guard5069 = cond_wire911_out;
wire _guard5070 = early_reset_static_par0_go_out;
wire _guard5071 = _guard5069 & _guard5070;
wire _guard5072 = cond_wire871_out;
wire _guard5073 = early_reset_static_par0_go_out;
wire _guard5074 = _guard5072 & _guard5073;
wire _guard5075 = cond_wire895_out;
wire _guard5076 = early_reset_static_par0_go_out;
wire _guard5077 = _guard5075 & _guard5076;
wire _guard5078 = cond_wire903_out;
wire _guard5079 = early_reset_static_par0_go_out;
wire _guard5080 = _guard5078 & _guard5079;
wire _guard5081 = cond_wire891_out;
wire _guard5082 = early_reset_static_par0_go_out;
wire _guard5083 = _guard5081 & _guard5082;
wire _guard5084 = cond_wire907_out;
wire _guard5085 = early_reset_static_par0_go_out;
wire _guard5086 = _guard5084 & _guard5085;
wire _guard5087 = cond_wire879_out;
wire _guard5088 = early_reset_static_par0_go_out;
wire _guard5089 = _guard5087 & _guard5088;
wire _guard5090 = cond_wire887_out;
wire _guard5091 = early_reset_static_par0_go_out;
wire _guard5092 = _guard5090 & _guard5091;
wire _guard5093 = cond_wire899_out;
wire _guard5094 = early_reset_static_par0_go_out;
wire _guard5095 = _guard5093 & _guard5094;
wire _guard5096 = cond_wire919_out;
wire _guard5097 = early_reset_static_par0_go_out;
wire _guard5098 = _guard5096 & _guard5097;
wire _guard5099 = cond_wire903_out;
wire _guard5100 = early_reset_static_par0_go_out;
wire _guard5101 = _guard5099 & _guard5100;
wire _guard5102 = cond_wire891_out;
wire _guard5103 = early_reset_static_par0_go_out;
wire _guard5104 = _guard5102 & _guard5103;
wire _guard5105 = cond_wire863_out;
wire _guard5106 = early_reset_static_par0_go_out;
wire _guard5107 = _guard5105 & _guard5106;
wire _guard5108 = cond_wire875_out;
wire _guard5109 = early_reset_static_par0_go_out;
wire _guard5110 = _guard5108 & _guard5109;
wire _guard5111 = cond_wire915_out;
wire _guard5112 = early_reset_static_par0_go_out;
wire _guard5113 = _guard5111 & _guard5112;
wire _guard5114 = cond_wire883_out;
wire _guard5115 = early_reset_static_par0_go_out;
wire _guard5116 = _guard5114 & _guard5115;
wire _guard5117 = cond_wire887_out;
wire _guard5118 = early_reset_static_par0_go_out;
wire _guard5119 = _guard5117 & _guard5118;
wire _guard5120 = cond_wire895_out;
wire _guard5121 = early_reset_static_par0_go_out;
wire _guard5122 = _guard5120 & _guard5121;
wire _guard5123 = cond_wire911_out;
wire _guard5124 = early_reset_static_par0_go_out;
wire _guard5125 = _guard5123 & _guard5124;
wire _guard5126 = cond_wire867_out;
wire _guard5127 = early_reset_static_par0_go_out;
wire _guard5128 = _guard5126 & _guard5127;
wire _guard5129 = cond_wire907_out;
wire _guard5130 = early_reset_static_par0_go_out;
wire _guard5131 = _guard5129 & _guard5130;
wire _guard5132 = cond_wire879_out;
wire _guard5133 = early_reset_static_par0_go_out;
wire _guard5134 = _guard5132 & _guard5133;
wire _guard5135 = cond_wire899_out;
wire _guard5136 = early_reset_static_par0_go_out;
wire _guard5137 = _guard5135 & _guard5136;
wire _guard5138 = cond_wire923_out;
wire _guard5139 = early_reset_static_par0_go_out;
wire _guard5140 = _guard5138 & _guard5139;
wire _guard5141 = cond_wire871_out;
wire _guard5142 = early_reset_static_par0_go_out;
wire _guard5143 = _guard5141 & _guard5142;
wire _guard5144 = cond_wire932_out;
wire _guard5145 = early_reset_static_par0_go_out;
wire _guard5146 = _guard5144 & _guard5145;
wire _guard5147 = cond_wire988_out;
wire _guard5148 = early_reset_static_par0_go_out;
wire _guard5149 = _guard5147 & _guard5148;
wire _guard5150 = cond_wire928_out;
wire _guard5151 = early_reset_static_par0_go_out;
wire _guard5152 = _guard5150 & _guard5151;
wire _guard5153 = cond_wire940_out;
wire _guard5154 = early_reset_static_par0_go_out;
wire _guard5155 = _guard5153 & _guard5154;
wire _guard5156 = cond_wire980_out;
wire _guard5157 = early_reset_static_par0_go_out;
wire _guard5158 = _guard5156 & _guard5157;
wire _guard5159 = cond_wire984_out;
wire _guard5160 = early_reset_static_par0_go_out;
wire _guard5161 = _guard5159 & _guard5160;
wire _guard5162 = cond_wire948_out;
wire _guard5163 = early_reset_static_par0_go_out;
wire _guard5164 = _guard5162 & _guard5163;
wire _guard5165 = cond_wire976_out;
wire _guard5166 = early_reset_static_par0_go_out;
wire _guard5167 = _guard5165 & _guard5166;
wire _guard5168 = cond_wire936_out;
wire _guard5169 = early_reset_static_par0_go_out;
wire _guard5170 = _guard5168 & _guard5169;
wire _guard5171 = cond_wire960_out;
wire _guard5172 = early_reset_static_par0_go_out;
wire _guard5173 = _guard5171 & _guard5172;
wire _guard5174 = cond_wire968_out;
wire _guard5175 = early_reset_static_par0_go_out;
wire _guard5176 = _guard5174 & _guard5175;
wire _guard5177 = cond_wire956_out;
wire _guard5178 = early_reset_static_par0_go_out;
wire _guard5179 = _guard5177 & _guard5178;
wire _guard5180 = cond_wire972_out;
wire _guard5181 = early_reset_static_par0_go_out;
wire _guard5182 = _guard5180 & _guard5181;
wire _guard5183 = cond_wire944_out;
wire _guard5184 = early_reset_static_par0_go_out;
wire _guard5185 = _guard5183 & _guard5184;
wire _guard5186 = cond_wire952_out;
wire _guard5187 = early_reset_static_par0_go_out;
wire _guard5188 = _guard5186 & _guard5187;
wire _guard5189 = cond_wire964_out;
wire _guard5190 = early_reset_static_par0_go_out;
wire _guard5191 = _guard5189 & _guard5190;
wire _guard5192 = cond_wire980_out;
wire _guard5193 = early_reset_static_par0_go_out;
wire _guard5194 = _guard5192 & _guard5193;
wire _guard5195 = cond_wire932_out;
wire _guard5196 = early_reset_static_par0_go_out;
wire _guard5197 = _guard5195 & _guard5196;
wire _guard5198 = cond_wire956_out;
wire _guard5199 = early_reset_static_par0_go_out;
wire _guard5200 = _guard5198 & _guard5199;
wire _guard5201 = cond_wire960_out;
wire _guard5202 = early_reset_static_par0_go_out;
wire _guard5203 = _guard5201 & _guard5202;
wire _guard5204 = cond_wire964_out;
wire _guard5205 = early_reset_static_par0_go_out;
wire _guard5206 = _guard5204 & _guard5205;
wire _guard5207 = cond_wire984_out;
wire _guard5208 = early_reset_static_par0_go_out;
wire _guard5209 = _guard5207 & _guard5208;
wire _guard5210 = cond_wire944_out;
wire _guard5211 = early_reset_static_par0_go_out;
wire _guard5212 = _guard5210 & _guard5211;
wire _guard5213 = cond_wire976_out;
wire _guard5214 = early_reset_static_par0_go_out;
wire _guard5215 = _guard5213 & _guard5214;
wire _guard5216 = cond_wire988_out;
wire _guard5217 = early_reset_static_par0_go_out;
wire _guard5218 = _guard5216 & _guard5217;
wire _guard5219 = cond_wire928_out;
wire _guard5220 = early_reset_static_par0_go_out;
wire _guard5221 = _guard5219 & _guard5220;
wire _guard5222 = cond_wire948_out;
wire _guard5223 = early_reset_static_par0_go_out;
wire _guard5224 = _guard5222 & _guard5223;
wire _guard5225 = cond_wire952_out;
wire _guard5226 = early_reset_static_par0_go_out;
wire _guard5227 = _guard5225 & _guard5226;
wire _guard5228 = cond_wire940_out;
wire _guard5229 = early_reset_static_par0_go_out;
wire _guard5230 = _guard5228 & _guard5229;
wire _guard5231 = cond_wire968_out;
wire _guard5232 = early_reset_static_par0_go_out;
wire _guard5233 = _guard5231 & _guard5232;
wire _guard5234 = cond_wire936_out;
wire _guard5235 = early_reset_static_par0_go_out;
wire _guard5236 = _guard5234 & _guard5235;
wire _guard5237 = cond_wire972_out;
wire _guard5238 = early_reset_static_par0_go_out;
wire _guard5239 = _guard5237 & _guard5238;
wire _guard5240 = cond_wire1001_out;
wire _guard5241 = early_reset_static_par0_go_out;
wire _guard5242 = _guard5240 & _guard5241;
wire _guard5243 = cond_wire1049_out;
wire _guard5244 = early_reset_static_par0_go_out;
wire _guard5245 = _guard5243 & _guard5244;
wire _guard5246 = cond_wire1029_out;
wire _guard5247 = early_reset_static_par0_go_out;
wire _guard5248 = _guard5246 & _guard5247;
wire _guard5249 = cond_wire1045_out;
wire _guard5250 = early_reset_static_par0_go_out;
wire _guard5251 = _guard5249 & _guard5250;
wire _guard5252 = cond_wire993_out;
wire _guard5253 = early_reset_static_par0_go_out;
wire _guard5254 = _guard5252 & _guard5253;
wire _guard5255 = cond_wire1041_out;
wire _guard5256 = early_reset_static_par0_go_out;
wire _guard5257 = _guard5255 & _guard5256;
wire _guard5258 = cond_wire1037_out;
wire _guard5259 = early_reset_static_par0_go_out;
wire _guard5260 = _guard5258 & _guard5259;
wire _guard5261 = cond_wire1009_out;
wire _guard5262 = early_reset_static_par0_go_out;
wire _guard5263 = _guard5261 & _guard5262;
wire _guard5264 = cond_wire1005_out;
wire _guard5265 = early_reset_static_par0_go_out;
wire _guard5266 = _guard5264 & _guard5265;
wire _guard5267 = cond_wire1017_out;
wire _guard5268 = early_reset_static_par0_go_out;
wire _guard5269 = _guard5267 & _guard5268;
wire _guard5270 = cond_wire1052_out;
wire _guard5271 = early_reset_static_par0_go_out;
wire _guard5272 = _guard5270 & _guard5271;
wire _guard5273 = cond_wire1021_out;
wire _guard5274 = early_reset_static_par0_go_out;
wire _guard5275 = _guard5273 & _guard5274;
wire _guard5276 = cond_wire997_out;
wire _guard5277 = early_reset_static_par0_go_out;
wire _guard5278 = _guard5276 & _guard5277;
wire _guard5279 = cond_wire1013_out;
wire _guard5280 = early_reset_static_par0_go_out;
wire _guard5281 = _guard5279 & _guard5280;
wire _guard5282 = cond_wire1033_out;
wire _guard5283 = early_reset_static_par0_go_out;
wire _guard5284 = _guard5282 & _guard5283;
wire _guard5285 = cond_wire1025_out;
wire _guard5286 = early_reset_static_par0_go_out;
wire _guard5287 = _guard5285 & _guard5286;
wire _guard5288 = fsm_out == 1'd0;
wire _guard5289 = cond_wire993_out;
wire _guard5290 = _guard5288 & _guard5289;
wire _guard5291 = fsm_out == 1'd0;
wire _guard5292 = _guard5290 & _guard5291;
wire _guard5293 = fsm_out == 1'd0;
wire _guard5294 = cond_wire997_out;
wire _guard5295 = _guard5293 & _guard5294;
wire _guard5296 = fsm_out == 1'd0;
wire _guard5297 = _guard5295 & _guard5296;
wire _guard5298 = _guard5292 | _guard5297;
wire _guard5299 = fsm_out == 1'd0;
wire _guard5300 = cond_wire1001_out;
wire _guard5301 = _guard5299 & _guard5300;
wire _guard5302 = fsm_out == 1'd0;
wire _guard5303 = _guard5301 & _guard5302;
wire _guard5304 = _guard5298 | _guard5303;
wire _guard5305 = fsm_out == 1'd0;
wire _guard5306 = cond_wire1005_out;
wire _guard5307 = _guard5305 & _guard5306;
wire _guard5308 = fsm_out == 1'd0;
wire _guard5309 = _guard5307 & _guard5308;
wire _guard5310 = _guard5304 | _guard5309;
wire _guard5311 = fsm_out == 1'd0;
wire _guard5312 = cond_wire1009_out;
wire _guard5313 = _guard5311 & _guard5312;
wire _guard5314 = fsm_out == 1'd0;
wire _guard5315 = _guard5313 & _guard5314;
wire _guard5316 = _guard5310 | _guard5315;
wire _guard5317 = fsm_out == 1'd0;
wire _guard5318 = cond_wire1013_out;
wire _guard5319 = _guard5317 & _guard5318;
wire _guard5320 = fsm_out == 1'd0;
wire _guard5321 = _guard5319 & _guard5320;
wire _guard5322 = _guard5316 | _guard5321;
wire _guard5323 = fsm_out == 1'd0;
wire _guard5324 = cond_wire1017_out;
wire _guard5325 = _guard5323 & _guard5324;
wire _guard5326 = fsm_out == 1'd0;
wire _guard5327 = _guard5325 & _guard5326;
wire _guard5328 = _guard5322 | _guard5327;
wire _guard5329 = fsm_out == 1'd0;
wire _guard5330 = cond_wire1021_out;
wire _guard5331 = _guard5329 & _guard5330;
wire _guard5332 = fsm_out == 1'd0;
wire _guard5333 = _guard5331 & _guard5332;
wire _guard5334 = _guard5328 | _guard5333;
wire _guard5335 = fsm_out == 1'd0;
wire _guard5336 = cond_wire1025_out;
wire _guard5337 = _guard5335 & _guard5336;
wire _guard5338 = fsm_out == 1'd0;
wire _guard5339 = _guard5337 & _guard5338;
wire _guard5340 = _guard5334 | _guard5339;
wire _guard5341 = fsm_out == 1'd0;
wire _guard5342 = cond_wire1029_out;
wire _guard5343 = _guard5341 & _guard5342;
wire _guard5344 = fsm_out == 1'd0;
wire _guard5345 = _guard5343 & _guard5344;
wire _guard5346 = _guard5340 | _guard5345;
wire _guard5347 = fsm_out == 1'd0;
wire _guard5348 = cond_wire1033_out;
wire _guard5349 = _guard5347 & _guard5348;
wire _guard5350 = fsm_out == 1'd0;
wire _guard5351 = _guard5349 & _guard5350;
wire _guard5352 = _guard5346 | _guard5351;
wire _guard5353 = fsm_out == 1'd0;
wire _guard5354 = cond_wire1037_out;
wire _guard5355 = _guard5353 & _guard5354;
wire _guard5356 = fsm_out == 1'd0;
wire _guard5357 = _guard5355 & _guard5356;
wire _guard5358 = _guard5352 | _guard5357;
wire _guard5359 = fsm_out == 1'd0;
wire _guard5360 = cond_wire1041_out;
wire _guard5361 = _guard5359 & _guard5360;
wire _guard5362 = fsm_out == 1'd0;
wire _guard5363 = _guard5361 & _guard5362;
wire _guard5364 = _guard5358 | _guard5363;
wire _guard5365 = fsm_out == 1'd0;
wire _guard5366 = cond_wire1045_out;
wire _guard5367 = _guard5365 & _guard5366;
wire _guard5368 = fsm_out == 1'd0;
wire _guard5369 = _guard5367 & _guard5368;
wire _guard5370 = _guard5364 | _guard5369;
wire _guard5371 = fsm_out == 1'd0;
wire _guard5372 = cond_wire1049_out;
wire _guard5373 = _guard5371 & _guard5372;
wire _guard5374 = fsm_out == 1'd0;
wire _guard5375 = _guard5373 & _guard5374;
wire _guard5376 = _guard5370 | _guard5375;
wire _guard5377 = fsm_out == 1'd0;
wire _guard5378 = cond_wire1052_out;
wire _guard5379 = _guard5377 & _guard5378;
wire _guard5380 = fsm_out == 1'd0;
wire _guard5381 = _guard5379 & _guard5380;
wire _guard5382 = _guard5376 | _guard5381;
wire _guard5383 = early_reset_static_par0_go_out;
wire _guard5384 = _guard5382 & _guard5383;
wire _guard5385 = early_reset_static_par0_go_out;
wire _guard5386 = ~_guard0;
wire _guard5387 = early_reset_static_par0_go_out;
wire _guard5388 = _guard5386 & _guard5387;
wire _guard5389 = early_reset_static_par0_go_out;
wire _guard5390 = ~_guard0;
wire _guard5391 = early_reset_static_par0_go_out;
wire _guard5392 = _guard5390 & _guard5391;
wire _guard5393 = early_reset_static_par0_go_out;
wire _guard5394 = early_reset_static_par0_go_out;
wire _guard5395 = early_reset_static_par0_go_out;
wire _guard5396 = ~_guard0;
wire _guard5397 = early_reset_static_par0_go_out;
wire _guard5398 = _guard5396 & _guard5397;
wire _guard5399 = ~_guard0;
wire _guard5400 = early_reset_static_par0_go_out;
wire _guard5401 = _guard5399 & _guard5400;
wire _guard5402 = early_reset_static_par0_go_out;
wire _guard5403 = early_reset_static_par0_go_out;
wire _guard5404 = early_reset_static_par0_go_out;
wire _guard5405 = early_reset_static_par0_go_out;
wire _guard5406 = ~_guard0;
wire _guard5407 = early_reset_static_par0_go_out;
wire _guard5408 = _guard5406 & _guard5407;
wire _guard5409 = ~_guard0;
wire _guard5410 = early_reset_static_par0_go_out;
wire _guard5411 = _guard5409 & _guard5410;
wire _guard5412 = early_reset_static_par0_go_out;
wire _guard5413 = early_reset_static_par0_go_out;
wire _guard5414 = early_reset_static_par0_go_out;
wire _guard5415 = early_reset_static_par0_go_out;
wire _guard5416 = early_reset_static_par0_go_out;
wire _guard5417 = ~_guard0;
wire _guard5418 = early_reset_static_par0_go_out;
wire _guard5419 = _guard5417 & _guard5418;
wire _guard5420 = early_reset_static_par0_go_out;
wire _guard5421 = early_reset_static_par0_go_out;
wire _guard5422 = early_reset_static_par0_go_out;
wire _guard5423 = early_reset_static_par0_go_out;
wire _guard5424 = early_reset_static_par0_go_out;
wire _guard5425 = early_reset_static_par0_go_out;
wire _guard5426 = early_reset_static_par0_go_out;
wire _guard5427 = early_reset_static_par0_go_out;
wire _guard5428 = ~_guard0;
wire _guard5429 = early_reset_static_par0_go_out;
wire _guard5430 = _guard5428 & _guard5429;
wire _guard5431 = early_reset_static_par0_go_out;
wire _guard5432 = early_reset_static_par0_go_out;
wire _guard5433 = ~_guard0;
wire _guard5434 = early_reset_static_par0_go_out;
wire _guard5435 = _guard5433 & _guard5434;
wire _guard5436 = early_reset_static_par0_go_out;
wire _guard5437 = early_reset_static_par0_go_out;
wire _guard5438 = early_reset_static_par0_go_out;
wire _guard5439 = ~_guard0;
wire _guard5440 = early_reset_static_par0_go_out;
wire _guard5441 = _guard5439 & _guard5440;
wire _guard5442 = early_reset_static_par0_go_out;
wire _guard5443 = ~_guard0;
wire _guard5444 = early_reset_static_par0_go_out;
wire _guard5445 = _guard5443 & _guard5444;
wire _guard5446 = early_reset_static_par0_go_out;
wire _guard5447 = early_reset_static_par0_go_out;
wire _guard5448 = ~_guard0;
wire _guard5449 = early_reset_static_par0_go_out;
wire _guard5450 = _guard5448 & _guard5449;
wire _guard5451 = early_reset_static_par0_go_out;
wire _guard5452 = early_reset_static_par0_go_out;
wire _guard5453 = early_reset_static_par0_go_out;
wire _guard5454 = early_reset_static_par0_go_out;
wire _guard5455 = early_reset_static_par0_go_out;
wire _guard5456 = ~_guard0;
wire _guard5457 = early_reset_static_par0_go_out;
wire _guard5458 = _guard5456 & _guard5457;
wire _guard5459 = early_reset_static_par0_go_out;
wire _guard5460 = early_reset_static_par0_go_out;
wire _guard5461 = early_reset_static_par0_go_out;
wire _guard5462 = early_reset_static_par0_go_out;
wire _guard5463 = early_reset_static_par0_go_out;
wire _guard5464 = early_reset_static_par0_go_out;
wire _guard5465 = ~_guard0;
wire _guard5466 = early_reset_static_par0_go_out;
wire _guard5467 = _guard5465 & _guard5466;
wire _guard5468 = early_reset_static_par0_go_out;
wire _guard5469 = early_reset_static_par0_go_out;
wire _guard5470 = early_reset_static_par0_go_out;
wire _guard5471 = ~_guard0;
wire _guard5472 = early_reset_static_par0_go_out;
wire _guard5473 = _guard5471 & _guard5472;
wire _guard5474 = early_reset_static_par0_go_out;
wire _guard5475 = early_reset_static_par0_go_out;
wire _guard5476 = early_reset_static_par0_go_out;
wire _guard5477 = early_reset_static_par0_go_out;
wire _guard5478 = ~_guard0;
wire _guard5479 = early_reset_static_par0_go_out;
wire _guard5480 = _guard5478 & _guard5479;
wire _guard5481 = early_reset_static_par0_go_out;
wire _guard5482 = early_reset_static_par0_go_out;
wire _guard5483 = early_reset_static_par0_go_out;
wire _guard5484 = early_reset_static_par0_go_out;
wire _guard5485 = early_reset_static_par0_go_out;
wire _guard5486 = ~_guard0;
wire _guard5487 = early_reset_static_par0_go_out;
wire _guard5488 = _guard5486 & _guard5487;
wire _guard5489 = early_reset_static_par0_go_out;
wire _guard5490 = early_reset_static_par0_go_out;
wire _guard5491 = early_reset_static_par0_go_out;
wire _guard5492 = early_reset_static_par0_go_out;
wire _guard5493 = early_reset_static_par0_go_out;
wire _guard5494 = ~_guard0;
wire _guard5495 = early_reset_static_par0_go_out;
wire _guard5496 = _guard5494 & _guard5495;
wire _guard5497 = early_reset_static_par0_go_out;
wire _guard5498 = early_reset_static_par0_go_out;
wire _guard5499 = early_reset_static_par0_go_out;
wire _guard5500 = ~_guard0;
wire _guard5501 = early_reset_static_par0_go_out;
wire _guard5502 = _guard5500 & _guard5501;
wire _guard5503 = early_reset_static_par0_go_out;
wire _guard5504 = ~_guard0;
wire _guard5505 = early_reset_static_par0_go_out;
wire _guard5506 = _guard5504 & _guard5505;
wire _guard5507 = early_reset_static_par0_go_out;
wire _guard5508 = ~_guard0;
wire _guard5509 = early_reset_static_par0_go_out;
wire _guard5510 = _guard5508 & _guard5509;
wire _guard5511 = early_reset_static_par0_go_out;
wire _guard5512 = early_reset_static_par0_go_out;
wire _guard5513 = early_reset_static_par0_go_out;
wire _guard5514 = ~_guard0;
wire _guard5515 = early_reset_static_par0_go_out;
wire _guard5516 = _guard5514 & _guard5515;
wire _guard5517 = early_reset_static_par0_go_out;
wire _guard5518 = ~_guard0;
wire _guard5519 = early_reset_static_par0_go_out;
wire _guard5520 = _guard5518 & _guard5519;
wire _guard5521 = early_reset_static_par0_go_out;
wire _guard5522 = early_reset_static_par0_go_out;
wire _guard5523 = early_reset_static_par0_go_out;
wire _guard5524 = ~_guard0;
wire _guard5525 = early_reset_static_par0_go_out;
wire _guard5526 = _guard5524 & _guard5525;
wire _guard5527 = ~_guard0;
wire _guard5528 = early_reset_static_par0_go_out;
wire _guard5529 = _guard5527 & _guard5528;
wire _guard5530 = early_reset_static_par0_go_out;
wire _guard5531 = early_reset_static_par0_go_out;
wire _guard5532 = early_reset_static_par0_go_out;
wire _guard5533 = early_reset_static_par0_go_out;
wire _guard5534 = ~_guard0;
wire _guard5535 = early_reset_static_par0_go_out;
wire _guard5536 = _guard5534 & _guard5535;
wire _guard5537 = ~_guard0;
wire _guard5538 = early_reset_static_par0_go_out;
wire _guard5539 = _guard5537 & _guard5538;
wire _guard5540 = early_reset_static_par0_go_out;
wire _guard5541 = early_reset_static_par0_go_out;
wire _guard5542 = early_reset_static_par0_go_out;
wire _guard5543 = early_reset_static_par0_go_out;
wire _guard5544 = early_reset_static_par0_go_out;
wire _guard5545 = early_reset_static_par0_go_out;
wire _guard5546 = early_reset_static_par0_go_out;
wire _guard5547 = early_reset_static_par0_go_out;
wire _guard5548 = early_reset_static_par0_go_out;
wire _guard5549 = early_reset_static_par0_go_out;
wire _guard5550 = early_reset_static_par0_go_out;
wire _guard5551 = early_reset_static_par0_go_out;
wire _guard5552 = early_reset_static_par0_go_out;
wire _guard5553 = ~_guard0;
wire _guard5554 = early_reset_static_par0_go_out;
wire _guard5555 = _guard5553 & _guard5554;
wire _guard5556 = early_reset_static_par0_go_out;
wire _guard5557 = early_reset_static_par0_go_out;
wire _guard5558 = early_reset_static_par0_go_out;
wire _guard5559 = early_reset_static_par0_go_out;
wire _guard5560 = early_reset_static_par0_go_out;
wire _guard5561 = early_reset_static_par0_go_out;
wire _guard5562 = ~_guard0;
wire _guard5563 = early_reset_static_par0_go_out;
wire _guard5564 = _guard5562 & _guard5563;
wire _guard5565 = early_reset_static_par0_go_out;
wire _guard5566 = ~_guard0;
wire _guard5567 = early_reset_static_par0_go_out;
wire _guard5568 = _guard5566 & _guard5567;
wire _guard5569 = early_reset_static_par0_go_out;
wire _guard5570 = early_reset_static_par0_go_out;
wire _guard5571 = early_reset_static_par0_go_out;
wire _guard5572 = early_reset_static_par0_go_out;
wire _guard5573 = ~_guard0;
wire _guard5574 = early_reset_static_par0_go_out;
wire _guard5575 = _guard5573 & _guard5574;
wire _guard5576 = early_reset_static_par0_go_out;
wire _guard5577 = early_reset_static_par0_go_out;
wire _guard5578 = ~_guard0;
wire _guard5579 = early_reset_static_par0_go_out;
wire _guard5580 = _guard5578 & _guard5579;
wire _guard5581 = ~_guard0;
wire _guard5582 = early_reset_static_par0_go_out;
wire _guard5583 = _guard5581 & _guard5582;
wire _guard5584 = early_reset_static_par0_go_out;
wire _guard5585 = early_reset_static_par0_go_out;
wire _guard5586 = early_reset_static_par0_go_out;
wire _guard5587 = ~_guard0;
wire _guard5588 = early_reset_static_par0_go_out;
wire _guard5589 = _guard5587 & _guard5588;
wire _guard5590 = early_reset_static_par0_go_out;
wire _guard5591 = early_reset_static_par0_go_out;
wire _guard5592 = ~_guard0;
wire _guard5593 = early_reset_static_par0_go_out;
wire _guard5594 = _guard5592 & _guard5593;
wire _guard5595 = early_reset_static_par0_go_out;
wire _guard5596 = early_reset_static_par0_go_out;
wire _guard5597 = early_reset_static_par0_go_out;
wire _guard5598 = early_reset_static_par0_go_out;
wire _guard5599 = ~_guard0;
wire _guard5600 = early_reset_static_par0_go_out;
wire _guard5601 = _guard5599 & _guard5600;
wire _guard5602 = early_reset_static_par0_go_out;
wire _guard5603 = early_reset_static_par0_go_out;
wire _guard5604 = ~_guard0;
wire _guard5605 = early_reset_static_par0_go_out;
wire _guard5606 = _guard5604 & _guard5605;
wire _guard5607 = ~_guard0;
wire _guard5608 = early_reset_static_par0_go_out;
wire _guard5609 = _guard5607 & _guard5608;
wire _guard5610 = early_reset_static_par0_go_out;
wire _guard5611 = early_reset_static_par0_go_out;
wire _guard5612 = early_reset_static_par0_go_out;
wire _guard5613 = ~_guard0;
wire _guard5614 = early_reset_static_par0_go_out;
wire _guard5615 = _guard5613 & _guard5614;
wire _guard5616 = early_reset_static_par0_go_out;
wire _guard5617 = early_reset_static_par0_go_out;
wire _guard5618 = ~_guard0;
wire _guard5619 = early_reset_static_par0_go_out;
wire _guard5620 = _guard5618 & _guard5619;
wire _guard5621 = early_reset_static_par0_go_out;
wire _guard5622 = early_reset_static_par0_go_out;
wire _guard5623 = early_reset_static_par0_go_out;
wire _guard5624 = ~_guard0;
wire _guard5625 = early_reset_static_par0_go_out;
wire _guard5626 = _guard5624 & _guard5625;
wire _guard5627 = early_reset_static_par0_go_out;
wire _guard5628 = early_reset_static_par0_go_out;
wire _guard5629 = ~_guard0;
wire _guard5630 = early_reset_static_par0_go_out;
wire _guard5631 = _guard5629 & _guard5630;
wire _guard5632 = early_reset_static_par0_go_out;
wire _guard5633 = early_reset_static_par0_go_out;
wire _guard5634 = early_reset_static_par0_go_out;
wire _guard5635 = early_reset_static_par0_go_out;
wire _guard5636 = early_reset_static_par0_go_out;
wire _guard5637 = early_reset_static_par0_go_out;
wire _guard5638 = early_reset_static_par0_go_out;
wire _guard5639 = ~_guard0;
wire _guard5640 = early_reset_static_par0_go_out;
wire _guard5641 = _guard5639 & _guard5640;
wire _guard5642 = early_reset_static_par0_go_out;
wire _guard5643 = early_reset_static_par0_go_out;
wire _guard5644 = early_reset_static_par0_go_out;
wire _guard5645 = early_reset_static_par0_go_out;
wire _guard5646 = early_reset_static_par0_go_out;
wire _guard5647 = early_reset_static_par0_go_out;
wire _guard5648 = ~_guard0;
wire _guard5649 = early_reset_static_par0_go_out;
wire _guard5650 = _guard5648 & _guard5649;
wire _guard5651 = early_reset_static_par0_go_out;
wire _guard5652 = ~_guard0;
wire _guard5653 = early_reset_static_par0_go_out;
wire _guard5654 = _guard5652 & _guard5653;
wire _guard5655 = early_reset_static_par0_go_out;
wire _guard5656 = early_reset_static_par0_go_out;
wire _guard5657 = early_reset_static_par0_go_out;
wire _guard5658 = early_reset_static_par0_go_out;
wire _guard5659 = early_reset_static_par0_go_out;
wire _guard5660 = early_reset_static_par0_go_out;
wire _guard5661 = early_reset_static_par0_go_out;
wire _guard5662 = ~_guard0;
wire _guard5663 = early_reset_static_par0_go_out;
wire _guard5664 = _guard5662 & _guard5663;
wire _guard5665 = early_reset_static_par0_go_out;
wire _guard5666 = ~_guard0;
wire _guard5667 = early_reset_static_par0_go_out;
wire _guard5668 = _guard5666 & _guard5667;
wire _guard5669 = early_reset_static_par0_go_out;
wire _guard5670 = ~_guard0;
wire _guard5671 = early_reset_static_par0_go_out;
wire _guard5672 = _guard5670 & _guard5671;
wire _guard5673 = early_reset_static_par0_go_out;
wire _guard5674 = ~_guard0;
wire _guard5675 = early_reset_static_par0_go_out;
wire _guard5676 = _guard5674 & _guard5675;
wire _guard5677 = early_reset_static_par0_go_out;
wire _guard5678 = early_reset_static_par0_go_out;
wire _guard5679 = early_reset_static_par0_go_out;
wire _guard5680 = early_reset_static_par0_go_out;
wire _guard5681 = early_reset_static_par0_go_out;
wire _guard5682 = early_reset_static_par0_go_out;
wire _guard5683 = early_reset_static_par0_go_out;
wire _guard5684 = early_reset_static_par0_go_out;
wire _guard5685 = ~_guard0;
wire _guard5686 = early_reset_static_par0_go_out;
wire _guard5687 = _guard5685 & _guard5686;
wire _guard5688 = early_reset_static_par0_go_out;
wire _guard5689 = ~_guard0;
wire _guard5690 = early_reset_static_par0_go_out;
wire _guard5691 = _guard5689 & _guard5690;
wire _guard5692 = early_reset_static_par0_go_out;
wire _guard5693 = early_reset_static_par0_go_out;
wire _guard5694 = ~_guard0;
wire _guard5695 = early_reset_static_par0_go_out;
wire _guard5696 = _guard5694 & _guard5695;
wire _guard5697 = early_reset_static_par0_go_out;
wire _guard5698 = early_reset_static_par0_go_out;
wire _guard5699 = early_reset_static_par0_go_out;
wire _guard5700 = early_reset_static_par0_go_out;
wire _guard5701 = early_reset_static_par0_go_out;
wire _guard5702 = early_reset_static_par0_go_out;
wire _guard5703 = early_reset_static_par0_go_out;
wire _guard5704 = early_reset_static_par0_go_out;
wire _guard5705 = early_reset_static_par0_go_out;
wire _guard5706 = early_reset_static_par0_go_out;
wire _guard5707 = early_reset_static_par0_go_out;
wire _guard5708 = early_reset_static_par0_go_out;
wire _guard5709 = early_reset_static_par0_go_out;
wire _guard5710 = early_reset_static_par0_go_out;
wire _guard5711 = ~_guard0;
wire _guard5712 = early_reset_static_par0_go_out;
wire _guard5713 = _guard5711 & _guard5712;
wire _guard5714 = early_reset_static_par0_go_out;
wire _guard5715 = early_reset_static_par0_go_out;
wire _guard5716 = early_reset_static_par0_go_out;
wire _guard5717 = ~_guard0;
wire _guard5718 = early_reset_static_par0_go_out;
wire _guard5719 = _guard5717 & _guard5718;
wire _guard5720 = early_reset_static_par0_go_out;
wire _guard5721 = early_reset_static_par0_go_out;
wire _guard5722 = early_reset_static_par0_go_out;
wire _guard5723 = ~_guard0;
wire _guard5724 = early_reset_static_par0_go_out;
wire _guard5725 = _guard5723 & _guard5724;
wire _guard5726 = early_reset_static_par0_go_out;
wire _guard5727 = early_reset_static_par0_go_out;
wire _guard5728 = early_reset_static_par0_go_out;
wire _guard5729 = early_reset_static_par0_go_out;
wire _guard5730 = ~_guard0;
wire _guard5731 = early_reset_static_par0_go_out;
wire _guard5732 = _guard5730 & _guard5731;
wire _guard5733 = early_reset_static_par0_go_out;
wire _guard5734 = early_reset_static_par0_go_out;
wire _guard5735 = early_reset_static_par0_go_out;
wire _guard5736 = early_reset_static_par0_go_out;
wire _guard5737 = early_reset_static_par0_go_out;
wire _guard5738 = ~_guard0;
wire _guard5739 = early_reset_static_par0_go_out;
wire _guard5740 = _guard5738 & _guard5739;
wire _guard5741 = ~_guard0;
wire _guard5742 = early_reset_static_par0_go_out;
wire _guard5743 = _guard5741 & _guard5742;
wire _guard5744 = early_reset_static_par0_go_out;
wire _guard5745 = early_reset_static_par0_go_out;
wire _guard5746 = ~_guard0;
wire _guard5747 = early_reset_static_par0_go_out;
wire _guard5748 = _guard5746 & _guard5747;
wire _guard5749 = early_reset_static_par0_go_out;
wire _guard5750 = ~_guard0;
wire _guard5751 = early_reset_static_par0_go_out;
wire _guard5752 = _guard5750 & _guard5751;
wire _guard5753 = early_reset_static_par0_go_out;
wire _guard5754 = early_reset_static_par0_go_out;
wire _guard5755 = ~_guard0;
wire _guard5756 = early_reset_static_par0_go_out;
wire _guard5757 = _guard5755 & _guard5756;
wire _guard5758 = early_reset_static_par0_go_out;
wire _guard5759 = ~_guard0;
wire _guard5760 = early_reset_static_par0_go_out;
wire _guard5761 = _guard5759 & _guard5760;
wire _guard5762 = early_reset_static_par0_go_out;
wire _guard5763 = ~_guard0;
wire _guard5764 = early_reset_static_par0_go_out;
wire _guard5765 = _guard5763 & _guard5764;
wire _guard5766 = early_reset_static_par0_go_out;
wire _guard5767 = early_reset_static_par0_go_out;
wire _guard5768 = ~_guard0;
wire _guard5769 = early_reset_static_par0_go_out;
wire _guard5770 = _guard5768 & _guard5769;
wire _guard5771 = early_reset_static_par0_go_out;
wire _guard5772 = early_reset_static_par0_go_out;
wire _guard5773 = early_reset_static_par0_go_out;
wire _guard5774 = early_reset_static_par0_go_out;
wire _guard5775 = early_reset_static_par0_go_out;
wire _guard5776 = early_reset_static_par0_go_out;
wire _guard5777 = early_reset_static_par0_go_out;
wire _guard5778 = early_reset_static_par0_go_out;
wire _guard5779 = ~_guard0;
wire _guard5780 = early_reset_static_par0_go_out;
wire _guard5781 = _guard5779 & _guard5780;
wire _guard5782 = early_reset_static_par0_go_out;
wire _guard5783 = early_reset_static_par0_go_out;
wire _guard5784 = early_reset_static_par0_go_out;
wire _guard5785 = early_reset_static_par0_go_out;
wire _guard5786 = ~_guard0;
wire _guard5787 = early_reset_static_par0_go_out;
wire _guard5788 = _guard5786 & _guard5787;
wire _guard5789 = ~_guard0;
wire _guard5790 = early_reset_static_par0_go_out;
wire _guard5791 = _guard5789 & _guard5790;
wire _guard5792 = early_reset_static_par0_go_out;
wire _guard5793 = early_reset_static_par0_go_out;
wire _guard5794 = early_reset_static_par0_go_out;
wire _guard5795 = early_reset_static_par0_go_out;
wire _guard5796 = ~_guard0;
wire _guard5797 = early_reset_static_par0_go_out;
wire _guard5798 = _guard5796 & _guard5797;
wire _guard5799 = early_reset_static_par0_go_out;
wire _guard5800 = early_reset_static_par0_go_out;
wire _guard5801 = ~_guard0;
wire _guard5802 = early_reset_static_par0_go_out;
wire _guard5803 = _guard5801 & _guard5802;
wire _guard5804 = early_reset_static_par0_go_out;
wire _guard5805 = early_reset_static_par0_go_out;
wire _guard5806 = early_reset_static_par0_go_out;
wire _guard5807 = ~_guard0;
wire _guard5808 = early_reset_static_par0_go_out;
wire _guard5809 = _guard5807 & _guard5808;
wire _guard5810 = early_reset_static_par0_go_out;
wire _guard5811 = early_reset_static_par0_go_out;
wire _guard5812 = ~_guard0;
wire _guard5813 = early_reset_static_par0_go_out;
wire _guard5814 = _guard5812 & _guard5813;
wire _guard5815 = early_reset_static_par0_go_out;
wire _guard5816 = early_reset_static_par0_go_out;
wire _guard5817 = early_reset_static_par0_go_out;
wire _guard5818 = early_reset_static_par0_go_out;
wire _guard5819 = early_reset_static_par0_go_out;
wire _guard5820 = early_reset_static_par0_go_out;
wire _guard5821 = early_reset_static_par0_go_out;
wire _guard5822 = early_reset_static_par0_go_out;
wire _guard5823 = early_reset_static_par0_go_out;
wire _guard5824 = fsm_out == 1'd0;
wire _guard5825 = early_reset_static_par0_go_out;
wire _guard5826 = _guard5824 & _guard5825;
wire _guard5827 = fsm_out != 1'd0;
wire _guard5828 = early_reset_static_par0_go_out;
wire _guard5829 = _guard5827 & _guard5828;
wire _guard5830 = early_reset_static_seq_go_out;
wire _guard5831 = early_reset_static_seq_go_out;
wire _guard5832 = fsm0_out >= 6'd1;
wire _guard5833 = fsm0_out < 6'd53;
wire _guard5834 = _guard5832 & _guard5833;
wire _guard5835 = early_reset_static_seq_go_out;
wire _guard5836 = _guard5834 & _guard5835;
wire _guard5837 = cond_wire29_out;
wire _guard5838 = early_reset_static_par0_go_out;
wire _guard5839 = _guard5837 & _guard5838;
wire _guard5840 = cond_wire29_out;
wire _guard5841 = early_reset_static_par0_go_out;
wire _guard5842 = _guard5840 & _guard5841;
wire _guard5843 = cond_wire74_out;
wire _guard5844 = early_reset_static_par0_go_out;
wire _guard5845 = _guard5843 & _guard5844;
wire _guard5846 = cond_wire74_out;
wire _guard5847 = early_reset_static_par0_go_out;
wire _guard5848 = _guard5846 & _guard5847;
wire _guard5849 = cond_wire93_out;
wire _guard5850 = early_reset_static_par0_go_out;
wire _guard5851 = _guard5849 & _guard5850;
wire _guard5852 = cond_wire93_out;
wire _guard5853 = early_reset_static_par0_go_out;
wire _guard5854 = _guard5852 & _guard5853;
wire _guard5855 = cond_wire26_out;
wire _guard5856 = early_reset_static_par0_go_out;
wire _guard5857 = _guard5855 & _guard5856;
wire _guard5858 = cond_wire26_out;
wire _guard5859 = early_reset_static_par0_go_out;
wire _guard5860 = _guard5858 & _guard5859;
wire _guard5861 = cond_wire97_out;
wire _guard5862 = early_reset_static_par0_go_out;
wire _guard5863 = _guard5861 & _guard5862;
wire _guard5864 = cond_wire97_out;
wire _guard5865 = early_reset_static_par0_go_out;
wire _guard5866 = _guard5864 & _guard5865;
wire _guard5867 = cond_wire113_out;
wire _guard5868 = early_reset_static_par0_go_out;
wire _guard5869 = _guard5867 & _guard5868;
wire _guard5870 = cond_wire113_out;
wire _guard5871 = early_reset_static_par0_go_out;
wire _guard5872 = _guard5870 & _guard5871;
wire _guard5873 = cond_wire203_out;
wire _guard5874 = early_reset_static_par0_go_out;
wire _guard5875 = _guard5873 & _guard5874;
wire _guard5876 = cond_wire201_out;
wire _guard5877 = early_reset_static_par0_go_out;
wire _guard5878 = _guard5876 & _guard5877;
wire _guard5879 = fsm_out == 1'd0;
wire _guard5880 = cond_wire201_out;
wire _guard5881 = _guard5879 & _guard5880;
wire _guard5882 = fsm_out == 1'd0;
wire _guard5883 = _guard5881 & _guard5882;
wire _guard5884 = fsm_out == 1'd0;
wire _guard5885 = cond_wire203_out;
wire _guard5886 = _guard5884 & _guard5885;
wire _guard5887 = fsm_out == 1'd0;
wire _guard5888 = _guard5886 & _guard5887;
wire _guard5889 = _guard5883 | _guard5888;
wire _guard5890 = early_reset_static_par0_go_out;
wire _guard5891 = _guard5889 & _guard5890;
wire _guard5892 = fsm_out == 1'd0;
wire _guard5893 = cond_wire201_out;
wire _guard5894 = _guard5892 & _guard5893;
wire _guard5895 = fsm_out == 1'd0;
wire _guard5896 = _guard5894 & _guard5895;
wire _guard5897 = fsm_out == 1'd0;
wire _guard5898 = cond_wire203_out;
wire _guard5899 = _guard5897 & _guard5898;
wire _guard5900 = fsm_out == 1'd0;
wire _guard5901 = _guard5899 & _guard5900;
wire _guard5902 = _guard5896 | _guard5901;
wire _guard5903 = early_reset_static_par0_go_out;
wire _guard5904 = _guard5902 & _guard5903;
wire _guard5905 = fsm_out == 1'd0;
wire _guard5906 = cond_wire201_out;
wire _guard5907 = _guard5905 & _guard5906;
wire _guard5908 = fsm_out == 1'd0;
wire _guard5909 = _guard5907 & _guard5908;
wire _guard5910 = fsm_out == 1'd0;
wire _guard5911 = cond_wire203_out;
wire _guard5912 = _guard5910 & _guard5911;
wire _guard5913 = fsm_out == 1'd0;
wire _guard5914 = _guard5912 & _guard5913;
wire _guard5915 = _guard5909 | _guard5914;
wire _guard5916 = early_reset_static_par0_go_out;
wire _guard5917 = _guard5915 & _guard5916;
wire _guard5918 = cond_wire202_out;
wire _guard5919 = early_reset_static_par0_go_out;
wire _guard5920 = _guard5918 & _guard5919;
wire _guard5921 = cond_wire202_out;
wire _guard5922 = early_reset_static_par0_go_out;
wire _guard5923 = _guard5921 & _guard5922;
wire _guard5924 = cond_wire228_out;
wire _guard5925 = early_reset_static_par0_go_out;
wire _guard5926 = _guard5924 & _guard5925;
wire _guard5927 = cond_wire226_out;
wire _guard5928 = early_reset_static_par0_go_out;
wire _guard5929 = _guard5927 & _guard5928;
wire _guard5930 = fsm_out == 1'd0;
wire _guard5931 = cond_wire226_out;
wire _guard5932 = _guard5930 & _guard5931;
wire _guard5933 = fsm_out == 1'd0;
wire _guard5934 = _guard5932 & _guard5933;
wire _guard5935 = fsm_out == 1'd0;
wire _guard5936 = cond_wire228_out;
wire _guard5937 = _guard5935 & _guard5936;
wire _guard5938 = fsm_out == 1'd0;
wire _guard5939 = _guard5937 & _guard5938;
wire _guard5940 = _guard5934 | _guard5939;
wire _guard5941 = early_reset_static_par0_go_out;
wire _guard5942 = _guard5940 & _guard5941;
wire _guard5943 = fsm_out == 1'd0;
wire _guard5944 = cond_wire226_out;
wire _guard5945 = _guard5943 & _guard5944;
wire _guard5946 = fsm_out == 1'd0;
wire _guard5947 = _guard5945 & _guard5946;
wire _guard5948 = fsm_out == 1'd0;
wire _guard5949 = cond_wire228_out;
wire _guard5950 = _guard5948 & _guard5949;
wire _guard5951 = fsm_out == 1'd0;
wire _guard5952 = _guard5950 & _guard5951;
wire _guard5953 = _guard5947 | _guard5952;
wire _guard5954 = early_reset_static_par0_go_out;
wire _guard5955 = _guard5953 & _guard5954;
wire _guard5956 = fsm_out == 1'd0;
wire _guard5957 = cond_wire226_out;
wire _guard5958 = _guard5956 & _guard5957;
wire _guard5959 = fsm_out == 1'd0;
wire _guard5960 = _guard5958 & _guard5959;
wire _guard5961 = fsm_out == 1'd0;
wire _guard5962 = cond_wire228_out;
wire _guard5963 = _guard5961 & _guard5962;
wire _guard5964 = fsm_out == 1'd0;
wire _guard5965 = _guard5963 & _guard5964;
wire _guard5966 = _guard5960 | _guard5965;
wire _guard5967 = early_reset_static_par0_go_out;
wire _guard5968 = _guard5966 & _guard5967;
wire _guard5969 = cond_wire240_out;
wire _guard5970 = early_reset_static_par0_go_out;
wire _guard5971 = _guard5969 & _guard5970;
wire _guard5972 = cond_wire238_out;
wire _guard5973 = early_reset_static_par0_go_out;
wire _guard5974 = _guard5972 & _guard5973;
wire _guard5975 = fsm_out == 1'd0;
wire _guard5976 = cond_wire238_out;
wire _guard5977 = _guard5975 & _guard5976;
wire _guard5978 = fsm_out == 1'd0;
wire _guard5979 = _guard5977 & _guard5978;
wire _guard5980 = fsm_out == 1'd0;
wire _guard5981 = cond_wire240_out;
wire _guard5982 = _guard5980 & _guard5981;
wire _guard5983 = fsm_out == 1'd0;
wire _guard5984 = _guard5982 & _guard5983;
wire _guard5985 = _guard5979 | _guard5984;
wire _guard5986 = early_reset_static_par0_go_out;
wire _guard5987 = _guard5985 & _guard5986;
wire _guard5988 = fsm_out == 1'd0;
wire _guard5989 = cond_wire238_out;
wire _guard5990 = _guard5988 & _guard5989;
wire _guard5991 = fsm_out == 1'd0;
wire _guard5992 = _guard5990 & _guard5991;
wire _guard5993 = fsm_out == 1'd0;
wire _guard5994 = cond_wire240_out;
wire _guard5995 = _guard5993 & _guard5994;
wire _guard5996 = fsm_out == 1'd0;
wire _guard5997 = _guard5995 & _guard5996;
wire _guard5998 = _guard5992 | _guard5997;
wire _guard5999 = early_reset_static_par0_go_out;
wire _guard6000 = _guard5998 & _guard5999;
wire _guard6001 = fsm_out == 1'd0;
wire _guard6002 = cond_wire238_out;
wire _guard6003 = _guard6001 & _guard6002;
wire _guard6004 = fsm_out == 1'd0;
wire _guard6005 = _guard6003 & _guard6004;
wire _guard6006 = fsm_out == 1'd0;
wire _guard6007 = cond_wire240_out;
wire _guard6008 = _guard6006 & _guard6007;
wire _guard6009 = fsm_out == 1'd0;
wire _guard6010 = _guard6008 & _guard6009;
wire _guard6011 = _guard6005 | _guard6010;
wire _guard6012 = early_reset_static_par0_go_out;
wire _guard6013 = _guard6011 & _guard6012;
wire _guard6014 = cond_wire178_out;
wire _guard6015 = early_reset_static_par0_go_out;
wire _guard6016 = _guard6014 & _guard6015;
wire _guard6017 = cond_wire178_out;
wire _guard6018 = early_reset_static_par0_go_out;
wire _guard6019 = _guard6017 & _guard6018;
wire _guard6020 = cond_wire243_out;
wire _guard6021 = early_reset_static_par0_go_out;
wire _guard6022 = _guard6020 & _guard6021;
wire _guard6023 = cond_wire243_out;
wire _guard6024 = early_reset_static_par0_go_out;
wire _guard6025 = _guard6023 & _guard6024;
wire _guard6026 = cond_wire190_out;
wire _guard6027 = early_reset_static_par0_go_out;
wire _guard6028 = _guard6026 & _guard6027;
wire _guard6029 = cond_wire190_out;
wire _guard6030 = early_reset_static_par0_go_out;
wire _guard6031 = _guard6029 & _guard6030;
wire _guard6032 = cond_wire255_out;
wire _guard6033 = early_reset_static_par0_go_out;
wire _guard6034 = _guard6032 & _guard6033;
wire _guard6035 = cond_wire255_out;
wire _guard6036 = early_reset_static_par0_go_out;
wire _guard6037 = _guard6035 & _guard6036;
wire _guard6038 = cond_wire277_out;
wire _guard6039 = early_reset_static_par0_go_out;
wire _guard6040 = _guard6038 & _guard6039;
wire _guard6041 = cond_wire275_out;
wire _guard6042 = early_reset_static_par0_go_out;
wire _guard6043 = _guard6041 & _guard6042;
wire _guard6044 = fsm_out == 1'd0;
wire _guard6045 = cond_wire275_out;
wire _guard6046 = _guard6044 & _guard6045;
wire _guard6047 = fsm_out == 1'd0;
wire _guard6048 = _guard6046 & _guard6047;
wire _guard6049 = fsm_out == 1'd0;
wire _guard6050 = cond_wire277_out;
wire _guard6051 = _guard6049 & _guard6050;
wire _guard6052 = fsm_out == 1'd0;
wire _guard6053 = _guard6051 & _guard6052;
wire _guard6054 = _guard6048 | _guard6053;
wire _guard6055 = early_reset_static_par0_go_out;
wire _guard6056 = _guard6054 & _guard6055;
wire _guard6057 = fsm_out == 1'd0;
wire _guard6058 = cond_wire275_out;
wire _guard6059 = _guard6057 & _guard6058;
wire _guard6060 = fsm_out == 1'd0;
wire _guard6061 = _guard6059 & _guard6060;
wire _guard6062 = fsm_out == 1'd0;
wire _guard6063 = cond_wire277_out;
wire _guard6064 = _guard6062 & _guard6063;
wire _guard6065 = fsm_out == 1'd0;
wire _guard6066 = _guard6064 & _guard6065;
wire _guard6067 = _guard6061 | _guard6066;
wire _guard6068 = early_reset_static_par0_go_out;
wire _guard6069 = _guard6067 & _guard6068;
wire _guard6070 = fsm_out == 1'd0;
wire _guard6071 = cond_wire275_out;
wire _guard6072 = _guard6070 & _guard6071;
wire _guard6073 = fsm_out == 1'd0;
wire _guard6074 = _guard6072 & _guard6073;
wire _guard6075 = fsm_out == 1'd0;
wire _guard6076 = cond_wire277_out;
wire _guard6077 = _guard6075 & _guard6076;
wire _guard6078 = fsm_out == 1'd0;
wire _guard6079 = _guard6077 & _guard6078;
wire _guard6080 = _guard6074 | _guard6079;
wire _guard6081 = early_reset_static_par0_go_out;
wire _guard6082 = _guard6080 & _guard6081;
wire _guard6083 = cond_wire280_out;
wire _guard6084 = early_reset_static_par0_go_out;
wire _guard6085 = _guard6083 & _guard6084;
wire _guard6086 = cond_wire280_out;
wire _guard6087 = early_reset_static_par0_go_out;
wire _guard6088 = _guard6086 & _guard6087;
wire _guard6089 = cond_wire342_out;
wire _guard6090 = early_reset_static_par0_go_out;
wire _guard6091 = _guard6089 & _guard6090;
wire _guard6092 = cond_wire340_out;
wire _guard6093 = early_reset_static_par0_go_out;
wire _guard6094 = _guard6092 & _guard6093;
wire _guard6095 = fsm_out == 1'd0;
wire _guard6096 = cond_wire340_out;
wire _guard6097 = _guard6095 & _guard6096;
wire _guard6098 = fsm_out == 1'd0;
wire _guard6099 = _guard6097 & _guard6098;
wire _guard6100 = fsm_out == 1'd0;
wire _guard6101 = cond_wire342_out;
wire _guard6102 = _guard6100 & _guard6101;
wire _guard6103 = fsm_out == 1'd0;
wire _guard6104 = _guard6102 & _guard6103;
wire _guard6105 = _guard6099 | _guard6104;
wire _guard6106 = early_reset_static_par0_go_out;
wire _guard6107 = _guard6105 & _guard6106;
wire _guard6108 = fsm_out == 1'd0;
wire _guard6109 = cond_wire340_out;
wire _guard6110 = _guard6108 & _guard6109;
wire _guard6111 = fsm_out == 1'd0;
wire _guard6112 = _guard6110 & _guard6111;
wire _guard6113 = fsm_out == 1'd0;
wire _guard6114 = cond_wire342_out;
wire _guard6115 = _guard6113 & _guard6114;
wire _guard6116 = fsm_out == 1'd0;
wire _guard6117 = _guard6115 & _guard6116;
wire _guard6118 = _guard6112 | _guard6117;
wire _guard6119 = early_reset_static_par0_go_out;
wire _guard6120 = _guard6118 & _guard6119;
wire _guard6121 = fsm_out == 1'd0;
wire _guard6122 = cond_wire340_out;
wire _guard6123 = _guard6121 & _guard6122;
wire _guard6124 = fsm_out == 1'd0;
wire _guard6125 = _guard6123 & _guard6124;
wire _guard6126 = fsm_out == 1'd0;
wire _guard6127 = cond_wire342_out;
wire _guard6128 = _guard6126 & _guard6127;
wire _guard6129 = fsm_out == 1'd0;
wire _guard6130 = _guard6128 & _guard6129;
wire _guard6131 = _guard6125 | _guard6130;
wire _guard6132 = early_reset_static_par0_go_out;
wire _guard6133 = _guard6131 & _guard6132;
wire _guard6134 = cond_wire361_out;
wire _guard6135 = early_reset_static_par0_go_out;
wire _guard6136 = _guard6134 & _guard6135;
wire _guard6137 = cond_wire361_out;
wire _guard6138 = early_reset_static_par0_go_out;
wire _guard6139 = _guard6137 & _guard6138;
wire _guard6140 = cond_wire336_out;
wire _guard6141 = early_reset_static_par0_go_out;
wire _guard6142 = _guard6140 & _guard6141;
wire _guard6143 = cond_wire336_out;
wire _guard6144 = early_reset_static_par0_go_out;
wire _guard6145 = _guard6143 & _guard6144;
wire _guard6146 = cond_wire422_out;
wire _guard6147 = early_reset_static_par0_go_out;
wire _guard6148 = _guard6146 & _guard6147;
wire _guard6149 = cond_wire422_out;
wire _guard6150 = early_reset_static_par0_go_out;
wire _guard6151 = _guard6149 & _guard6150;
wire _guard6152 = cond_wire365_out;
wire _guard6153 = early_reset_static_par0_go_out;
wire _guard6154 = _guard6152 & _guard6153;
wire _guard6155 = cond_wire365_out;
wire _guard6156 = early_reset_static_par0_go_out;
wire _guard6157 = _guard6155 & _guard6156;
wire _guard6158 = cond_wire451_out;
wire _guard6159 = early_reset_static_par0_go_out;
wire _guard6160 = _guard6158 & _guard6159;
wire _guard6161 = cond_wire449_out;
wire _guard6162 = early_reset_static_par0_go_out;
wire _guard6163 = _guard6161 & _guard6162;
wire _guard6164 = fsm_out == 1'd0;
wire _guard6165 = cond_wire449_out;
wire _guard6166 = _guard6164 & _guard6165;
wire _guard6167 = fsm_out == 1'd0;
wire _guard6168 = _guard6166 & _guard6167;
wire _guard6169 = fsm_out == 1'd0;
wire _guard6170 = cond_wire451_out;
wire _guard6171 = _guard6169 & _guard6170;
wire _guard6172 = fsm_out == 1'd0;
wire _guard6173 = _guard6171 & _guard6172;
wire _guard6174 = _guard6168 | _guard6173;
wire _guard6175 = early_reset_static_par0_go_out;
wire _guard6176 = _guard6174 & _guard6175;
wire _guard6177 = fsm_out == 1'd0;
wire _guard6178 = cond_wire449_out;
wire _guard6179 = _guard6177 & _guard6178;
wire _guard6180 = fsm_out == 1'd0;
wire _guard6181 = _guard6179 & _guard6180;
wire _guard6182 = fsm_out == 1'd0;
wire _guard6183 = cond_wire451_out;
wire _guard6184 = _guard6182 & _guard6183;
wire _guard6185 = fsm_out == 1'd0;
wire _guard6186 = _guard6184 & _guard6185;
wire _guard6187 = _guard6181 | _guard6186;
wire _guard6188 = early_reset_static_par0_go_out;
wire _guard6189 = _guard6187 & _guard6188;
wire _guard6190 = fsm_out == 1'd0;
wire _guard6191 = cond_wire449_out;
wire _guard6192 = _guard6190 & _guard6191;
wire _guard6193 = fsm_out == 1'd0;
wire _guard6194 = _guard6192 & _guard6193;
wire _guard6195 = fsm_out == 1'd0;
wire _guard6196 = cond_wire451_out;
wire _guard6197 = _guard6195 & _guard6196;
wire _guard6198 = fsm_out == 1'd0;
wire _guard6199 = _guard6197 & _guard6198;
wire _guard6200 = _guard6194 | _guard6199;
wire _guard6201 = early_reset_static_par0_go_out;
wire _guard6202 = _guard6200 & _guard6201;
wire _guard6203 = cond_wire515_out;
wire _guard6204 = early_reset_static_par0_go_out;
wire _guard6205 = _guard6203 & _guard6204;
wire _guard6206 = cond_wire515_out;
wire _guard6207 = early_reset_static_par0_go_out;
wire _guard6208 = _guard6206 & _guard6207;
wire _guard6209 = cond_wire532_out;
wire _guard6210 = early_reset_static_par0_go_out;
wire _guard6211 = _guard6209 & _guard6210;
wire _guard6212 = cond_wire530_out;
wire _guard6213 = early_reset_static_par0_go_out;
wire _guard6214 = _guard6212 & _guard6213;
wire _guard6215 = fsm_out == 1'd0;
wire _guard6216 = cond_wire530_out;
wire _guard6217 = _guard6215 & _guard6216;
wire _guard6218 = fsm_out == 1'd0;
wire _guard6219 = _guard6217 & _guard6218;
wire _guard6220 = fsm_out == 1'd0;
wire _guard6221 = cond_wire532_out;
wire _guard6222 = _guard6220 & _guard6221;
wire _guard6223 = fsm_out == 1'd0;
wire _guard6224 = _guard6222 & _guard6223;
wire _guard6225 = _guard6219 | _guard6224;
wire _guard6226 = early_reset_static_par0_go_out;
wire _guard6227 = _guard6225 & _guard6226;
wire _guard6228 = fsm_out == 1'd0;
wire _guard6229 = cond_wire530_out;
wire _guard6230 = _guard6228 & _guard6229;
wire _guard6231 = fsm_out == 1'd0;
wire _guard6232 = _guard6230 & _guard6231;
wire _guard6233 = fsm_out == 1'd0;
wire _guard6234 = cond_wire532_out;
wire _guard6235 = _guard6233 & _guard6234;
wire _guard6236 = fsm_out == 1'd0;
wire _guard6237 = _guard6235 & _guard6236;
wire _guard6238 = _guard6232 | _guard6237;
wire _guard6239 = early_reset_static_par0_go_out;
wire _guard6240 = _guard6238 & _guard6239;
wire _guard6241 = fsm_out == 1'd0;
wire _guard6242 = cond_wire530_out;
wire _guard6243 = _guard6241 & _guard6242;
wire _guard6244 = fsm_out == 1'd0;
wire _guard6245 = _guard6243 & _guard6244;
wire _guard6246 = fsm_out == 1'd0;
wire _guard6247 = cond_wire532_out;
wire _guard6248 = _guard6246 & _guard6247;
wire _guard6249 = fsm_out == 1'd0;
wire _guard6250 = _guard6248 & _guard6249;
wire _guard6251 = _guard6245 | _guard6250;
wire _guard6252 = early_reset_static_par0_go_out;
wire _guard6253 = _guard6251 & _guard6252;
wire _guard6254 = cond_wire499_out;
wire _guard6255 = early_reset_static_par0_go_out;
wire _guard6256 = _guard6254 & _guard6255;
wire _guard6257 = cond_wire499_out;
wire _guard6258 = early_reset_static_par0_go_out;
wire _guard6259 = _guard6257 & _guard6258;
wire _guard6260 = cond_wire572_out;
wire _guard6261 = early_reset_static_par0_go_out;
wire _guard6262 = _guard6260 & _guard6261;
wire _guard6263 = cond_wire572_out;
wire _guard6264 = early_reset_static_par0_go_out;
wire _guard6265 = _guard6263 & _guard6264;
wire _guard6266 = cond_wire630_out;
wire _guard6267 = early_reset_static_par0_go_out;
wire _guard6268 = _guard6266 & _guard6267;
wire _guard6269 = cond_wire628_out;
wire _guard6270 = early_reset_static_par0_go_out;
wire _guard6271 = _guard6269 & _guard6270;
wire _guard6272 = fsm_out == 1'd0;
wire _guard6273 = cond_wire628_out;
wire _guard6274 = _guard6272 & _guard6273;
wire _guard6275 = fsm_out == 1'd0;
wire _guard6276 = _guard6274 & _guard6275;
wire _guard6277 = fsm_out == 1'd0;
wire _guard6278 = cond_wire630_out;
wire _guard6279 = _guard6277 & _guard6278;
wire _guard6280 = fsm_out == 1'd0;
wire _guard6281 = _guard6279 & _guard6280;
wire _guard6282 = _guard6276 | _guard6281;
wire _guard6283 = early_reset_static_par0_go_out;
wire _guard6284 = _guard6282 & _guard6283;
wire _guard6285 = fsm_out == 1'd0;
wire _guard6286 = cond_wire628_out;
wire _guard6287 = _guard6285 & _guard6286;
wire _guard6288 = fsm_out == 1'd0;
wire _guard6289 = _guard6287 & _guard6288;
wire _guard6290 = fsm_out == 1'd0;
wire _guard6291 = cond_wire630_out;
wire _guard6292 = _guard6290 & _guard6291;
wire _guard6293 = fsm_out == 1'd0;
wire _guard6294 = _guard6292 & _guard6293;
wire _guard6295 = _guard6289 | _guard6294;
wire _guard6296 = early_reset_static_par0_go_out;
wire _guard6297 = _guard6295 & _guard6296;
wire _guard6298 = fsm_out == 1'd0;
wire _guard6299 = cond_wire628_out;
wire _guard6300 = _guard6298 & _guard6299;
wire _guard6301 = fsm_out == 1'd0;
wire _guard6302 = _guard6300 & _guard6301;
wire _guard6303 = fsm_out == 1'd0;
wire _guard6304 = cond_wire630_out;
wire _guard6305 = _guard6303 & _guard6304;
wire _guard6306 = fsm_out == 1'd0;
wire _guard6307 = _guard6305 & _guard6306;
wire _guard6308 = _guard6302 | _guard6307;
wire _guard6309 = early_reset_static_par0_go_out;
wire _guard6310 = _guard6308 & _guard6309;
wire _guard6311 = cond_wire686_out;
wire _guard6312 = early_reset_static_par0_go_out;
wire _guard6313 = _guard6311 & _guard6312;
wire _guard6314 = cond_wire686_out;
wire _guard6315 = early_reset_static_par0_go_out;
wire _guard6316 = _guard6314 & _guard6315;
wire _guard6317 = cond_wire764_out;
wire _guard6318 = early_reset_static_par0_go_out;
wire _guard6319 = _guard6317 & _guard6318;
wire _guard6320 = cond_wire762_out;
wire _guard6321 = early_reset_static_par0_go_out;
wire _guard6322 = _guard6320 & _guard6321;
wire _guard6323 = fsm_out == 1'd0;
wire _guard6324 = cond_wire762_out;
wire _guard6325 = _guard6323 & _guard6324;
wire _guard6326 = fsm_out == 1'd0;
wire _guard6327 = _guard6325 & _guard6326;
wire _guard6328 = fsm_out == 1'd0;
wire _guard6329 = cond_wire764_out;
wire _guard6330 = _guard6328 & _guard6329;
wire _guard6331 = fsm_out == 1'd0;
wire _guard6332 = _guard6330 & _guard6331;
wire _guard6333 = _guard6327 | _guard6332;
wire _guard6334 = early_reset_static_par0_go_out;
wire _guard6335 = _guard6333 & _guard6334;
wire _guard6336 = fsm_out == 1'd0;
wire _guard6337 = cond_wire762_out;
wire _guard6338 = _guard6336 & _guard6337;
wire _guard6339 = fsm_out == 1'd0;
wire _guard6340 = _guard6338 & _guard6339;
wire _guard6341 = fsm_out == 1'd0;
wire _guard6342 = cond_wire764_out;
wire _guard6343 = _guard6341 & _guard6342;
wire _guard6344 = fsm_out == 1'd0;
wire _guard6345 = _guard6343 & _guard6344;
wire _guard6346 = _guard6340 | _guard6345;
wire _guard6347 = early_reset_static_par0_go_out;
wire _guard6348 = _guard6346 & _guard6347;
wire _guard6349 = fsm_out == 1'd0;
wire _guard6350 = cond_wire762_out;
wire _guard6351 = _guard6349 & _guard6350;
wire _guard6352 = fsm_out == 1'd0;
wire _guard6353 = _guard6351 & _guard6352;
wire _guard6354 = fsm_out == 1'd0;
wire _guard6355 = cond_wire764_out;
wire _guard6356 = _guard6354 & _guard6355;
wire _guard6357 = fsm_out == 1'd0;
wire _guard6358 = _guard6356 & _guard6357;
wire _guard6359 = _guard6353 | _guard6358;
wire _guard6360 = early_reset_static_par0_go_out;
wire _guard6361 = _guard6359 & _guard6360;
wire _guard6362 = cond_wire710_out;
wire _guard6363 = early_reset_static_par0_go_out;
wire _guard6364 = _guard6362 & _guard6363;
wire _guard6365 = cond_wire710_out;
wire _guard6366 = early_reset_static_par0_go_out;
wire _guard6367 = _guard6365 & _guard6366;
wire _guard6368 = cond_wire792_out;
wire _guard6369 = early_reset_static_par0_go_out;
wire _guard6370 = _guard6368 & _guard6369;
wire _guard6371 = cond_wire790_out;
wire _guard6372 = early_reset_static_par0_go_out;
wire _guard6373 = _guard6371 & _guard6372;
wire _guard6374 = fsm_out == 1'd0;
wire _guard6375 = cond_wire790_out;
wire _guard6376 = _guard6374 & _guard6375;
wire _guard6377 = fsm_out == 1'd0;
wire _guard6378 = _guard6376 & _guard6377;
wire _guard6379 = fsm_out == 1'd0;
wire _guard6380 = cond_wire792_out;
wire _guard6381 = _guard6379 & _guard6380;
wire _guard6382 = fsm_out == 1'd0;
wire _guard6383 = _guard6381 & _guard6382;
wire _guard6384 = _guard6378 | _guard6383;
wire _guard6385 = early_reset_static_par0_go_out;
wire _guard6386 = _guard6384 & _guard6385;
wire _guard6387 = fsm_out == 1'd0;
wire _guard6388 = cond_wire790_out;
wire _guard6389 = _guard6387 & _guard6388;
wire _guard6390 = fsm_out == 1'd0;
wire _guard6391 = _guard6389 & _guard6390;
wire _guard6392 = fsm_out == 1'd0;
wire _guard6393 = cond_wire792_out;
wire _guard6394 = _guard6392 & _guard6393;
wire _guard6395 = fsm_out == 1'd0;
wire _guard6396 = _guard6394 & _guard6395;
wire _guard6397 = _guard6391 | _guard6396;
wire _guard6398 = early_reset_static_par0_go_out;
wire _guard6399 = _guard6397 & _guard6398;
wire _guard6400 = fsm_out == 1'd0;
wire _guard6401 = cond_wire790_out;
wire _guard6402 = _guard6400 & _guard6401;
wire _guard6403 = fsm_out == 1'd0;
wire _guard6404 = _guard6402 & _guard6403;
wire _guard6405 = fsm_out == 1'd0;
wire _guard6406 = cond_wire792_out;
wire _guard6407 = _guard6405 & _guard6406;
wire _guard6408 = fsm_out == 1'd0;
wire _guard6409 = _guard6407 & _guard6408;
wire _guard6410 = _guard6404 | _guard6409;
wire _guard6411 = early_reset_static_par0_go_out;
wire _guard6412 = _guard6410 & _guard6411;
wire _guard6413 = cond_wire812_out;
wire _guard6414 = early_reset_static_par0_go_out;
wire _guard6415 = _guard6413 & _guard6414;
wire _guard6416 = cond_wire812_out;
wire _guard6417 = early_reset_static_par0_go_out;
wire _guard6418 = _guard6416 & _guard6417;
wire _guard6419 = cond_wire833_out;
wire _guard6420 = early_reset_static_par0_go_out;
wire _guard6421 = _guard6419 & _guard6420;
wire _guard6422 = cond_wire831_out;
wire _guard6423 = early_reset_static_par0_go_out;
wire _guard6424 = _guard6422 & _guard6423;
wire _guard6425 = fsm_out == 1'd0;
wire _guard6426 = cond_wire831_out;
wire _guard6427 = _guard6425 & _guard6426;
wire _guard6428 = fsm_out == 1'd0;
wire _guard6429 = _guard6427 & _guard6428;
wire _guard6430 = fsm_out == 1'd0;
wire _guard6431 = cond_wire833_out;
wire _guard6432 = _guard6430 & _guard6431;
wire _guard6433 = fsm_out == 1'd0;
wire _guard6434 = _guard6432 & _guard6433;
wire _guard6435 = _guard6429 | _guard6434;
wire _guard6436 = early_reset_static_par0_go_out;
wire _guard6437 = _guard6435 & _guard6436;
wire _guard6438 = fsm_out == 1'd0;
wire _guard6439 = cond_wire831_out;
wire _guard6440 = _guard6438 & _guard6439;
wire _guard6441 = fsm_out == 1'd0;
wire _guard6442 = _guard6440 & _guard6441;
wire _guard6443 = fsm_out == 1'd0;
wire _guard6444 = cond_wire833_out;
wire _guard6445 = _guard6443 & _guard6444;
wire _guard6446 = fsm_out == 1'd0;
wire _guard6447 = _guard6445 & _guard6446;
wire _guard6448 = _guard6442 | _guard6447;
wire _guard6449 = early_reset_static_par0_go_out;
wire _guard6450 = _guard6448 & _guard6449;
wire _guard6451 = fsm_out == 1'd0;
wire _guard6452 = cond_wire831_out;
wire _guard6453 = _guard6451 & _guard6452;
wire _guard6454 = fsm_out == 1'd0;
wire _guard6455 = _guard6453 & _guard6454;
wire _guard6456 = fsm_out == 1'd0;
wire _guard6457 = cond_wire833_out;
wire _guard6458 = _guard6456 & _guard6457;
wire _guard6459 = fsm_out == 1'd0;
wire _guard6460 = _guard6458 & _guard6459;
wire _guard6461 = _guard6455 | _guard6460;
wire _guard6462 = early_reset_static_par0_go_out;
wire _guard6463 = _guard6461 & _guard6462;
wire _guard6464 = cond_wire845_out;
wire _guard6465 = early_reset_static_par0_go_out;
wire _guard6466 = _guard6464 & _guard6465;
wire _guard6467 = cond_wire843_out;
wire _guard6468 = early_reset_static_par0_go_out;
wire _guard6469 = _guard6467 & _guard6468;
wire _guard6470 = fsm_out == 1'd0;
wire _guard6471 = cond_wire843_out;
wire _guard6472 = _guard6470 & _guard6471;
wire _guard6473 = fsm_out == 1'd0;
wire _guard6474 = _guard6472 & _guard6473;
wire _guard6475 = fsm_out == 1'd0;
wire _guard6476 = cond_wire845_out;
wire _guard6477 = _guard6475 & _guard6476;
wire _guard6478 = fsm_out == 1'd0;
wire _guard6479 = _guard6477 & _guard6478;
wire _guard6480 = _guard6474 | _guard6479;
wire _guard6481 = early_reset_static_par0_go_out;
wire _guard6482 = _guard6480 & _guard6481;
wire _guard6483 = fsm_out == 1'd0;
wire _guard6484 = cond_wire843_out;
wire _guard6485 = _guard6483 & _guard6484;
wire _guard6486 = fsm_out == 1'd0;
wire _guard6487 = _guard6485 & _guard6486;
wire _guard6488 = fsm_out == 1'd0;
wire _guard6489 = cond_wire845_out;
wire _guard6490 = _guard6488 & _guard6489;
wire _guard6491 = fsm_out == 1'd0;
wire _guard6492 = _guard6490 & _guard6491;
wire _guard6493 = _guard6487 | _guard6492;
wire _guard6494 = early_reset_static_par0_go_out;
wire _guard6495 = _guard6493 & _guard6494;
wire _guard6496 = fsm_out == 1'd0;
wire _guard6497 = cond_wire843_out;
wire _guard6498 = _guard6496 & _guard6497;
wire _guard6499 = fsm_out == 1'd0;
wire _guard6500 = _guard6498 & _guard6499;
wire _guard6501 = fsm_out == 1'd0;
wire _guard6502 = cond_wire845_out;
wire _guard6503 = _guard6501 & _guard6502;
wire _guard6504 = fsm_out == 1'd0;
wire _guard6505 = _guard6503 & _guard6504;
wire _guard6506 = _guard6500 | _guard6505;
wire _guard6507 = early_reset_static_par0_go_out;
wire _guard6508 = _guard6506 & _guard6507;
wire _guard6509 = cond_wire787_out;
wire _guard6510 = early_reset_static_par0_go_out;
wire _guard6511 = _guard6509 & _guard6510;
wire _guard6512 = cond_wire787_out;
wire _guard6513 = early_reset_static_par0_go_out;
wire _guard6514 = _guard6512 & _guard6513;
wire _guard6515 = cond_wire796_out;
wire _guard6516 = early_reset_static_par0_go_out;
wire _guard6517 = _guard6515 & _guard6516;
wire _guard6518 = cond_wire796_out;
wire _guard6519 = early_reset_static_par0_go_out;
wire _guard6520 = _guard6518 & _guard6519;
wire _guard6521 = cond_wire836_out;
wire _guard6522 = early_reset_static_par0_go_out;
wire _guard6523 = _guard6521 & _guard6522;
wire _guard6524 = cond_wire836_out;
wire _guard6525 = early_reset_static_par0_go_out;
wire _guard6526 = _guard6524 & _guard6525;
wire _guard6527 = cond_wire954_out;
wire _guard6528 = early_reset_static_par0_go_out;
wire _guard6529 = _guard6527 & _guard6528;
wire _guard6530 = cond_wire954_out;
wire _guard6531 = early_reset_static_par0_go_out;
wire _guard6532 = _guard6530 & _guard6531;
wire _guard6533 = cond_wire909_out;
wire _guard6534 = early_reset_static_par0_go_out;
wire _guard6535 = _guard6533 & _guard6534;
wire _guard6536 = cond_wire909_out;
wire _guard6537 = early_reset_static_par0_go_out;
wire _guard6538 = _guard6536 & _guard6537;
wire _guard6539 = cond_wire979_out;
wire _guard6540 = early_reset_static_par0_go_out;
wire _guard6541 = _guard6539 & _guard6540;
wire _guard6542 = cond_wire977_out;
wire _guard6543 = early_reset_static_par0_go_out;
wire _guard6544 = _guard6542 & _guard6543;
wire _guard6545 = fsm_out == 1'd0;
wire _guard6546 = cond_wire977_out;
wire _guard6547 = _guard6545 & _guard6546;
wire _guard6548 = fsm_out == 1'd0;
wire _guard6549 = _guard6547 & _guard6548;
wire _guard6550 = fsm_out == 1'd0;
wire _guard6551 = cond_wire979_out;
wire _guard6552 = _guard6550 & _guard6551;
wire _guard6553 = fsm_out == 1'd0;
wire _guard6554 = _guard6552 & _guard6553;
wire _guard6555 = _guard6549 | _guard6554;
wire _guard6556 = early_reset_static_par0_go_out;
wire _guard6557 = _guard6555 & _guard6556;
wire _guard6558 = fsm_out == 1'd0;
wire _guard6559 = cond_wire977_out;
wire _guard6560 = _guard6558 & _guard6559;
wire _guard6561 = fsm_out == 1'd0;
wire _guard6562 = _guard6560 & _guard6561;
wire _guard6563 = fsm_out == 1'd0;
wire _guard6564 = cond_wire979_out;
wire _guard6565 = _guard6563 & _guard6564;
wire _guard6566 = fsm_out == 1'd0;
wire _guard6567 = _guard6565 & _guard6566;
wire _guard6568 = _guard6562 | _guard6567;
wire _guard6569 = early_reset_static_par0_go_out;
wire _guard6570 = _guard6568 & _guard6569;
wire _guard6571 = fsm_out == 1'd0;
wire _guard6572 = cond_wire977_out;
wire _guard6573 = _guard6571 & _guard6572;
wire _guard6574 = fsm_out == 1'd0;
wire _guard6575 = _guard6573 & _guard6574;
wire _guard6576 = fsm_out == 1'd0;
wire _guard6577 = cond_wire979_out;
wire _guard6578 = _guard6576 & _guard6577;
wire _guard6579 = fsm_out == 1'd0;
wire _guard6580 = _guard6578 & _guard6579;
wire _guard6581 = _guard6575 | _guard6580;
wire _guard6582 = early_reset_static_par0_go_out;
wire _guard6583 = _guard6581 & _guard6582;
wire _guard6584 = cond_wire917_out;
wire _guard6585 = early_reset_static_par0_go_out;
wire _guard6586 = _guard6584 & _guard6585;
wire _guard6587 = cond_wire917_out;
wire _guard6588 = early_reset_static_par0_go_out;
wire _guard6589 = _guard6587 & _guard6588;
wire _guard6590 = cond_wire1000_out;
wire _guard6591 = early_reset_static_par0_go_out;
wire _guard6592 = _guard6590 & _guard6591;
wire _guard6593 = cond_wire998_out;
wire _guard6594 = early_reset_static_par0_go_out;
wire _guard6595 = _guard6593 & _guard6594;
wire _guard6596 = fsm_out == 1'd0;
wire _guard6597 = cond_wire998_out;
wire _guard6598 = _guard6596 & _guard6597;
wire _guard6599 = fsm_out == 1'd0;
wire _guard6600 = _guard6598 & _guard6599;
wire _guard6601 = fsm_out == 1'd0;
wire _guard6602 = cond_wire1000_out;
wire _guard6603 = _guard6601 & _guard6602;
wire _guard6604 = fsm_out == 1'd0;
wire _guard6605 = _guard6603 & _guard6604;
wire _guard6606 = _guard6600 | _guard6605;
wire _guard6607 = early_reset_static_par0_go_out;
wire _guard6608 = _guard6606 & _guard6607;
wire _guard6609 = fsm_out == 1'd0;
wire _guard6610 = cond_wire998_out;
wire _guard6611 = _guard6609 & _guard6610;
wire _guard6612 = fsm_out == 1'd0;
wire _guard6613 = _guard6611 & _guard6612;
wire _guard6614 = fsm_out == 1'd0;
wire _guard6615 = cond_wire1000_out;
wire _guard6616 = _guard6614 & _guard6615;
wire _guard6617 = fsm_out == 1'd0;
wire _guard6618 = _guard6616 & _guard6617;
wire _guard6619 = _guard6613 | _guard6618;
wire _guard6620 = early_reset_static_par0_go_out;
wire _guard6621 = _guard6619 & _guard6620;
wire _guard6622 = fsm_out == 1'd0;
wire _guard6623 = cond_wire998_out;
wire _guard6624 = _guard6622 & _guard6623;
wire _guard6625 = fsm_out == 1'd0;
wire _guard6626 = _guard6624 & _guard6625;
wire _guard6627 = fsm_out == 1'd0;
wire _guard6628 = cond_wire1000_out;
wire _guard6629 = _guard6627 & _guard6628;
wire _guard6630 = fsm_out == 1'd0;
wire _guard6631 = _guard6629 & _guard6630;
wire _guard6632 = _guard6626 | _guard6631;
wire _guard6633 = early_reset_static_par0_go_out;
wire _guard6634 = _guard6632 & _guard6633;
wire _guard6635 = cond_wire974_out;
wire _guard6636 = early_reset_static_par0_go_out;
wire _guard6637 = _guard6635 & _guard6636;
wire _guard6638 = cond_wire974_out;
wire _guard6639 = early_reset_static_par0_go_out;
wire _guard6640 = _guard6638 & _guard6639;
wire _guard6641 = fsm0_out == 6'd0;
wire _guard6642 = early_reset_static_seq_go_out;
wire _guard6643 = _guard6641 & _guard6642;
wire _guard6644 = cond_wire_out;
wire _guard6645 = early_reset_static_par0_go_out;
wire _guard6646 = _guard6644 & _guard6645;
wire _guard6647 = _guard6643 | _guard6646;
wire _guard6648 = fsm0_out == 6'd0;
wire _guard6649 = early_reset_static_seq_go_out;
wire _guard6650 = _guard6648 & _guard6649;
wire _guard6651 = cond_wire_out;
wire _guard6652 = early_reset_static_par0_go_out;
wire _guard6653 = _guard6651 & _guard6652;
wire _guard6654 = fsm0_out == 6'd0;
wire _guard6655 = early_reset_static_seq_go_out;
wire _guard6656 = _guard6654 & _guard6655;
wire _guard6657 = cond_wire729_out;
wire _guard6658 = early_reset_static_par0_go_out;
wire _guard6659 = _guard6657 & _guard6658;
wire _guard6660 = _guard6656 | _guard6659;
wire _guard6661 = fsm0_out == 6'd0;
wire _guard6662 = early_reset_static_seq_go_out;
wire _guard6663 = _guard6661 & _guard6662;
wire _guard6664 = cond_wire729_out;
wire _guard6665 = early_reset_static_par0_go_out;
wire _guard6666 = _guard6664 & _guard6665;
wire _guard6667 = fsm0_out == 6'd0;
wire _guard6668 = early_reset_static_seq_go_out;
wire _guard6669 = _guard6667 & _guard6668;
wire _guard6670 = early_reset_static_par0_go_out;
wire _guard6671 = _guard6669 | _guard6670;
wire _guard6672 = early_reset_static_par0_go_out;
wire _guard6673 = fsm0_out == 6'd0;
wire _guard6674 = early_reset_static_seq_go_out;
wire _guard6675 = _guard6673 & _guard6674;
wire _guard6676 = fsm0_out == 6'd0;
wire _guard6677 = early_reset_static_seq_go_out;
wire _guard6678 = _guard6676 & _guard6677;
wire _guard6679 = early_reset_static_par0_go_out;
wire _guard6680 = _guard6678 | _guard6679;
wire _guard6681 = fsm0_out == 6'd0;
wire _guard6682 = early_reset_static_seq_go_out;
wire _guard6683 = _guard6681 & _guard6682;
wire _guard6684 = early_reset_static_par0_go_out;
wire _guard6685 = early_reset_static_par0_go_out;
wire _guard6686 = early_reset_static_par0_go_out;
wire _guard6687 = early_reset_static_par0_go_out;
wire _guard6688 = early_reset_static_par0_go_out;
wire _guard6689 = early_reset_static_par0_go_out;
wire _guard6690 = early_reset_static_par0_go_out;
wire _guard6691 = early_reset_static_par0_go_out;
wire _guard6692 = early_reset_static_par0_go_out;
wire _guard6693 = early_reset_static_par0_go_out;
wire _guard6694 = early_reset_static_par0_go_out;
wire _guard6695 = fsm0_out == 6'd0;
wire _guard6696 = early_reset_static_seq_go_out;
wire _guard6697 = _guard6695 & _guard6696;
wire _guard6698 = early_reset_static_par0_go_out;
wire _guard6699 = _guard6697 | _guard6698;
wire _guard6700 = early_reset_static_par0_go_out;
wire _guard6701 = fsm0_out == 6'd0;
wire _guard6702 = early_reset_static_seq_go_out;
wire _guard6703 = _guard6701 & _guard6702;
wire _guard6704 = fsm0_out == 6'd0;
wire _guard6705 = early_reset_static_seq_go_out;
wire _guard6706 = _guard6704 & _guard6705;
wire _guard6707 = early_reset_static_par0_go_out;
wire _guard6708 = _guard6706 | _guard6707;
wire _guard6709 = early_reset_static_par0_go_out;
wire _guard6710 = fsm0_out == 6'd0;
wire _guard6711 = early_reset_static_seq_go_out;
wire _guard6712 = _guard6710 & _guard6711;
wire _guard6713 = early_reset_static_par0_go_out;
wire _guard6714 = early_reset_static_par0_go_out;
wire _guard6715 = early_reset_static_par0_go_out;
wire _guard6716 = early_reset_static_par0_go_out;
wire _guard6717 = fsm0_out == 6'd0;
wire _guard6718 = early_reset_static_seq_go_out;
wire _guard6719 = _guard6717 & _guard6718;
wire _guard6720 = early_reset_static_par0_go_out;
wire _guard6721 = _guard6719 | _guard6720;
wire _guard6722 = fsm0_out == 6'd0;
wire _guard6723 = early_reset_static_seq_go_out;
wire _guard6724 = _guard6722 & _guard6723;
wire _guard6725 = early_reset_static_par0_go_out;
wire _guard6726 = early_reset_static_par0_go_out;
wire _guard6727 = early_reset_static_par0_go_out;
wire _guard6728 = early_reset_static_par0_go_out;
wire _guard6729 = early_reset_static_par0_go_out;
wire _guard6730 = early_reset_static_par0_go_out;
wire _guard6731 = early_reset_static_par0_go_out;
wire _guard6732 = fsm0_out == 6'd0;
wire _guard6733 = early_reset_static_seq_go_out;
wire _guard6734 = _guard6732 & _guard6733;
wire _guard6735 = early_reset_static_par0_go_out;
wire _guard6736 = _guard6734 | _guard6735;
wire _guard6737 = early_reset_static_par0_go_out;
wire _guard6738 = fsm0_out == 6'd0;
wire _guard6739 = early_reset_static_seq_go_out;
wire _guard6740 = _guard6738 & _guard6739;
wire _guard6741 = early_reset_static_par0_go_out;
wire _guard6742 = early_reset_static_par0_go_out;
wire _guard6743 = early_reset_static_par0_go_out;
wire _guard6744 = early_reset_static_par0_go_out;
wire _guard6745 = ~_guard0;
wire _guard6746 = early_reset_static_par0_go_out;
wire _guard6747 = _guard6745 & _guard6746;
wire _guard6748 = early_reset_static_par0_go_out;
wire _guard6749 = early_reset_static_par0_go_out;
wire _guard6750 = early_reset_static_par0_go_out;
wire _guard6751 = ~_guard0;
wire _guard6752 = early_reset_static_par0_go_out;
wire _guard6753 = _guard6751 & _guard6752;
wire _guard6754 = early_reset_static_par0_go_out;
wire _guard6755 = ~_guard0;
wire _guard6756 = early_reset_static_par0_go_out;
wire _guard6757 = _guard6755 & _guard6756;
wire _guard6758 = early_reset_static_par0_go_out;
wire _guard6759 = early_reset_static_par0_go_out;
wire _guard6760 = early_reset_static_par0_go_out;
wire _guard6761 = ~_guard0;
wire _guard6762 = early_reset_static_par0_go_out;
wire _guard6763 = _guard6761 & _guard6762;
wire _guard6764 = early_reset_static_par0_go_out;
wire _guard6765 = early_reset_static_par0_go_out;
wire _guard6766 = ~_guard0;
wire _guard6767 = early_reset_static_par0_go_out;
wire _guard6768 = _guard6766 & _guard6767;
wire _guard6769 = early_reset_static_par0_go_out;
wire _guard6770 = early_reset_static_par0_go_out;
wire _guard6771 = early_reset_static_par0_go_out;
wire _guard6772 = ~_guard0;
wire _guard6773 = early_reset_static_par0_go_out;
wire _guard6774 = _guard6772 & _guard6773;
wire _guard6775 = early_reset_static_par0_go_out;
wire _guard6776 = early_reset_static_par0_go_out;
wire _guard6777 = early_reset_static_par0_go_out;
wire _guard6778 = early_reset_static_par0_go_out;
wire _guard6779 = early_reset_static_par0_go_out;
wire _guard6780 = early_reset_static_par0_go_out;
wire _guard6781 = early_reset_static_par0_go_out;
wire _guard6782 = early_reset_static_par0_go_out;
wire _guard6783 = early_reset_static_par0_go_out;
wire _guard6784 = early_reset_static_par0_go_out;
wire _guard6785 = early_reset_static_par0_go_out;
wire _guard6786 = ~_guard0;
wire _guard6787 = early_reset_static_par0_go_out;
wire _guard6788 = _guard6786 & _guard6787;
wire _guard6789 = early_reset_static_par0_go_out;
wire _guard6790 = ~_guard0;
wire _guard6791 = early_reset_static_par0_go_out;
wire _guard6792 = _guard6790 & _guard6791;
wire _guard6793 = ~_guard0;
wire _guard6794 = early_reset_static_par0_go_out;
wire _guard6795 = _guard6793 & _guard6794;
wire _guard6796 = early_reset_static_par0_go_out;
wire _guard6797 = early_reset_static_par0_go_out;
wire _guard6798 = early_reset_static_par0_go_out;
wire _guard6799 = early_reset_static_par0_go_out;
wire _guard6800 = early_reset_static_par0_go_out;
wire _guard6801 = early_reset_static_par0_go_out;
wire _guard6802 = ~_guard0;
wire _guard6803 = early_reset_static_par0_go_out;
wire _guard6804 = _guard6802 & _guard6803;
wire _guard6805 = ~_guard0;
wire _guard6806 = early_reset_static_par0_go_out;
wire _guard6807 = _guard6805 & _guard6806;
wire _guard6808 = early_reset_static_par0_go_out;
wire _guard6809 = early_reset_static_par0_go_out;
wire _guard6810 = early_reset_static_par0_go_out;
wire _guard6811 = early_reset_static_par0_go_out;
wire _guard6812 = early_reset_static_par0_go_out;
wire _guard6813 = early_reset_static_par0_go_out;
wire _guard6814 = early_reset_static_par0_go_out;
wire _guard6815 = ~_guard0;
wire _guard6816 = early_reset_static_par0_go_out;
wire _guard6817 = _guard6815 & _guard6816;
wire _guard6818 = early_reset_static_par0_go_out;
wire _guard6819 = early_reset_static_par0_go_out;
wire _guard6820 = early_reset_static_par0_go_out;
wire _guard6821 = early_reset_static_par0_go_out;
wire _guard6822 = early_reset_static_par0_go_out;
wire _guard6823 = early_reset_static_par0_go_out;
wire _guard6824 = ~_guard0;
wire _guard6825 = early_reset_static_par0_go_out;
wire _guard6826 = _guard6824 & _guard6825;
wire _guard6827 = ~_guard0;
wire _guard6828 = early_reset_static_par0_go_out;
wire _guard6829 = _guard6827 & _guard6828;
wire _guard6830 = early_reset_static_par0_go_out;
wire _guard6831 = early_reset_static_par0_go_out;
wire _guard6832 = ~_guard0;
wire _guard6833 = early_reset_static_par0_go_out;
wire _guard6834 = _guard6832 & _guard6833;
wire _guard6835 = early_reset_static_par0_go_out;
wire _guard6836 = early_reset_static_par0_go_out;
wire _guard6837 = ~_guard0;
wire _guard6838 = early_reset_static_par0_go_out;
wire _guard6839 = _guard6837 & _guard6838;
wire _guard6840 = early_reset_static_par0_go_out;
wire _guard6841 = early_reset_static_par0_go_out;
wire _guard6842 = early_reset_static_par0_go_out;
wire _guard6843 = early_reset_static_par0_go_out;
wire _guard6844 = early_reset_static_par0_go_out;
wire _guard6845 = early_reset_static_par0_go_out;
wire _guard6846 = early_reset_static_par0_go_out;
wire _guard6847 = early_reset_static_par0_go_out;
wire _guard6848 = early_reset_static_par0_go_out;
wire _guard6849 = early_reset_static_par0_go_out;
wire _guard6850 = ~_guard0;
wire _guard6851 = early_reset_static_par0_go_out;
wire _guard6852 = _guard6850 & _guard6851;
wire _guard6853 = ~_guard0;
wire _guard6854 = early_reset_static_par0_go_out;
wire _guard6855 = _guard6853 & _guard6854;
wire _guard6856 = early_reset_static_par0_go_out;
wire _guard6857 = early_reset_static_par0_go_out;
wire _guard6858 = early_reset_static_par0_go_out;
wire _guard6859 = early_reset_static_par0_go_out;
wire _guard6860 = ~_guard0;
wire _guard6861 = early_reset_static_par0_go_out;
wire _guard6862 = _guard6860 & _guard6861;
wire _guard6863 = early_reset_static_par0_go_out;
wire _guard6864 = early_reset_static_par0_go_out;
wire _guard6865 = ~_guard0;
wire _guard6866 = early_reset_static_par0_go_out;
wire _guard6867 = _guard6865 & _guard6866;
wire _guard6868 = early_reset_static_par0_go_out;
wire _guard6869 = early_reset_static_par0_go_out;
wire _guard6870 = early_reset_static_par0_go_out;
wire _guard6871 = ~_guard0;
wire _guard6872 = early_reset_static_par0_go_out;
wire _guard6873 = _guard6871 & _guard6872;
wire _guard6874 = early_reset_static_par0_go_out;
wire _guard6875 = early_reset_static_par0_go_out;
wire _guard6876 = ~_guard0;
wire _guard6877 = early_reset_static_par0_go_out;
wire _guard6878 = _guard6876 & _guard6877;
wire _guard6879 = ~_guard0;
wire _guard6880 = early_reset_static_par0_go_out;
wire _guard6881 = _guard6879 & _guard6880;
wire _guard6882 = early_reset_static_par0_go_out;
wire _guard6883 = ~_guard0;
wire _guard6884 = early_reset_static_par0_go_out;
wire _guard6885 = _guard6883 & _guard6884;
wire _guard6886 = early_reset_static_par0_go_out;
wire _guard6887 = ~_guard0;
wire _guard6888 = early_reset_static_par0_go_out;
wire _guard6889 = _guard6887 & _guard6888;
wire _guard6890 = early_reset_static_par0_go_out;
wire _guard6891 = early_reset_static_par0_go_out;
wire _guard6892 = early_reset_static_par0_go_out;
wire _guard6893 = ~_guard0;
wire _guard6894 = early_reset_static_par0_go_out;
wire _guard6895 = _guard6893 & _guard6894;
wire _guard6896 = early_reset_static_par0_go_out;
wire _guard6897 = ~_guard0;
wire _guard6898 = early_reset_static_par0_go_out;
wire _guard6899 = _guard6897 & _guard6898;
wire _guard6900 = early_reset_static_par0_go_out;
wire _guard6901 = early_reset_static_par0_go_out;
wire _guard6902 = ~_guard0;
wire _guard6903 = early_reset_static_par0_go_out;
wire _guard6904 = _guard6902 & _guard6903;
wire _guard6905 = ~_guard0;
wire _guard6906 = early_reset_static_par0_go_out;
wire _guard6907 = _guard6905 & _guard6906;
wire _guard6908 = early_reset_static_par0_go_out;
wire _guard6909 = early_reset_static_par0_go_out;
wire _guard6910 = ~_guard0;
wire _guard6911 = early_reset_static_par0_go_out;
wire _guard6912 = _guard6910 & _guard6911;
wire _guard6913 = early_reset_static_par0_go_out;
wire _guard6914 = early_reset_static_par0_go_out;
wire _guard6915 = early_reset_static_par0_go_out;
wire _guard6916 = early_reset_static_par0_go_out;
wire _guard6917 = early_reset_static_par0_go_out;
wire _guard6918 = early_reset_static_par0_go_out;
wire _guard6919 = ~_guard0;
wire _guard6920 = early_reset_static_par0_go_out;
wire _guard6921 = _guard6919 & _guard6920;
wire _guard6922 = early_reset_static_par0_go_out;
wire _guard6923 = early_reset_static_par0_go_out;
wire _guard6924 = early_reset_static_par0_go_out;
wire _guard6925 = ~_guard0;
wire _guard6926 = early_reset_static_par0_go_out;
wire _guard6927 = _guard6925 & _guard6926;
wire _guard6928 = early_reset_static_par0_go_out;
wire _guard6929 = early_reset_static_par0_go_out;
wire _guard6930 = early_reset_static_par0_go_out;
wire _guard6931 = ~_guard0;
wire _guard6932 = early_reset_static_par0_go_out;
wire _guard6933 = _guard6931 & _guard6932;
wire _guard6934 = early_reset_static_par0_go_out;
wire _guard6935 = early_reset_static_par0_go_out;
wire _guard6936 = early_reset_static_par0_go_out;
wire _guard6937 = ~_guard0;
wire _guard6938 = early_reset_static_par0_go_out;
wire _guard6939 = _guard6937 & _guard6938;
wire _guard6940 = early_reset_static_par0_go_out;
wire _guard6941 = early_reset_static_par0_go_out;
wire _guard6942 = ~_guard0;
wire _guard6943 = early_reset_static_par0_go_out;
wire _guard6944 = _guard6942 & _guard6943;
wire _guard6945 = early_reset_static_par0_go_out;
wire _guard6946 = ~_guard0;
wire _guard6947 = early_reset_static_par0_go_out;
wire _guard6948 = _guard6946 & _guard6947;
wire _guard6949 = ~_guard0;
wire _guard6950 = early_reset_static_par0_go_out;
wire _guard6951 = _guard6949 & _guard6950;
wire _guard6952 = early_reset_static_par0_go_out;
wire _guard6953 = early_reset_static_par0_go_out;
wire _guard6954 = ~_guard0;
wire _guard6955 = early_reset_static_par0_go_out;
wire _guard6956 = _guard6954 & _guard6955;
wire _guard6957 = early_reset_static_par0_go_out;
wire _guard6958 = early_reset_static_par0_go_out;
wire _guard6959 = early_reset_static_par0_go_out;
wire _guard6960 = ~_guard0;
wire _guard6961 = early_reset_static_par0_go_out;
wire _guard6962 = _guard6960 & _guard6961;
wire _guard6963 = early_reset_static_par0_go_out;
wire _guard6964 = ~_guard0;
wire _guard6965 = early_reset_static_par0_go_out;
wire _guard6966 = _guard6964 & _guard6965;
wire _guard6967 = early_reset_static_par0_go_out;
wire _guard6968 = early_reset_static_par0_go_out;
wire _guard6969 = early_reset_static_par0_go_out;
wire _guard6970 = early_reset_static_par0_go_out;
wire _guard6971 = early_reset_static_par0_go_out;
wire _guard6972 = early_reset_static_par0_go_out;
wire _guard6973 = early_reset_static_par0_go_out;
wire _guard6974 = early_reset_static_par0_go_out;
wire _guard6975 = early_reset_static_par0_go_out;
wire _guard6976 = early_reset_static_par0_go_out;
wire _guard6977 = early_reset_static_par0_go_out;
wire _guard6978 = ~_guard0;
wire _guard6979 = early_reset_static_par0_go_out;
wire _guard6980 = _guard6978 & _guard6979;
wire _guard6981 = ~_guard0;
wire _guard6982 = early_reset_static_par0_go_out;
wire _guard6983 = _guard6981 & _guard6982;
wire _guard6984 = early_reset_static_par0_go_out;
wire _guard6985 = ~_guard0;
wire _guard6986 = early_reset_static_par0_go_out;
wire _guard6987 = _guard6985 & _guard6986;
wire _guard6988 = early_reset_static_par0_go_out;
wire _guard6989 = early_reset_static_par0_go_out;
wire _guard6990 = ~_guard0;
wire _guard6991 = early_reset_static_par0_go_out;
wire _guard6992 = _guard6990 & _guard6991;
wire _guard6993 = early_reset_static_par0_go_out;
wire _guard6994 = early_reset_static_par0_go_out;
wire _guard6995 = early_reset_static_par0_go_out;
wire _guard6996 = early_reset_static_par0_go_out;
wire _guard6997 = early_reset_static_par0_go_out;
wire _guard6998 = early_reset_static_par0_go_out;
wire _guard6999 = early_reset_static_par0_go_out;
wire _guard7000 = ~_guard0;
wire _guard7001 = early_reset_static_par0_go_out;
wire _guard7002 = _guard7000 & _guard7001;
wire _guard7003 = ~_guard0;
wire _guard7004 = early_reset_static_par0_go_out;
wire _guard7005 = _guard7003 & _guard7004;
wire _guard7006 = early_reset_static_par0_go_out;
wire _guard7007 = early_reset_static_par0_go_out;
wire _guard7008 = early_reset_static_par0_go_out;
wire _guard7009 = early_reset_static_par0_go_out;
wire _guard7010 = early_reset_static_par0_go_out;
wire _guard7011 = ~_guard0;
wire _guard7012 = early_reset_static_par0_go_out;
wire _guard7013 = _guard7011 & _guard7012;
wire _guard7014 = early_reset_static_par0_go_out;
wire _guard7015 = early_reset_static_par0_go_out;
wire _guard7016 = ~_guard0;
wire _guard7017 = early_reset_static_par0_go_out;
wire _guard7018 = _guard7016 & _guard7017;
wire _guard7019 = early_reset_static_par0_go_out;
wire _guard7020 = ~_guard0;
wire _guard7021 = early_reset_static_par0_go_out;
wire _guard7022 = _guard7020 & _guard7021;
wire _guard7023 = ~_guard0;
wire _guard7024 = early_reset_static_par0_go_out;
wire _guard7025 = _guard7023 & _guard7024;
wire _guard7026 = early_reset_static_par0_go_out;
wire _guard7027 = early_reset_static_par0_go_out;
wire _guard7028 = early_reset_static_par0_go_out;
wire _guard7029 = early_reset_static_par0_go_out;
wire _guard7030 = early_reset_static_par0_go_out;
wire _guard7031 = early_reset_static_par0_go_out;
wire _guard7032 = ~_guard0;
wire _guard7033 = early_reset_static_par0_go_out;
wire _guard7034 = _guard7032 & _guard7033;
wire _guard7035 = early_reset_static_par0_go_out;
wire _guard7036 = early_reset_static_par0_go_out;
wire _guard7037 = early_reset_static_par0_go_out;
wire _guard7038 = early_reset_static_par0_go_out;
wire _guard7039 = ~_guard0;
wire _guard7040 = early_reset_static_par0_go_out;
wire _guard7041 = _guard7039 & _guard7040;
wire _guard7042 = early_reset_static_par0_go_out;
wire _guard7043 = early_reset_static_par0_go_out;
wire _guard7044 = early_reset_static_par0_go_out;
wire _guard7045 = early_reset_static_par0_go_out;
wire _guard7046 = early_reset_static_par0_go_out;
wire _guard7047 = early_reset_static_par0_go_out;
wire _guard7048 = ~_guard0;
wire _guard7049 = early_reset_static_par0_go_out;
wire _guard7050 = _guard7048 & _guard7049;
wire _guard7051 = ~_guard0;
wire _guard7052 = early_reset_static_par0_go_out;
wire _guard7053 = _guard7051 & _guard7052;
wire _guard7054 = early_reset_static_par0_go_out;
wire _guard7055 = ~_guard0;
wire _guard7056 = early_reset_static_par0_go_out;
wire _guard7057 = _guard7055 & _guard7056;
wire _guard7058 = early_reset_static_par0_go_out;
wire _guard7059 = early_reset_static_par0_go_out;
wire _guard7060 = ~_guard0;
wire _guard7061 = early_reset_static_par0_go_out;
wire _guard7062 = _guard7060 & _guard7061;
wire _guard7063 = early_reset_static_par0_go_out;
wire _guard7064 = early_reset_static_par0_go_out;
wire _guard7065 = ~_guard0;
wire _guard7066 = early_reset_static_par0_go_out;
wire _guard7067 = _guard7065 & _guard7066;
wire _guard7068 = early_reset_static_par0_go_out;
wire _guard7069 = ~_guard0;
wire _guard7070 = early_reset_static_par0_go_out;
wire _guard7071 = _guard7069 & _guard7070;
wire _guard7072 = early_reset_static_par0_go_out;
wire _guard7073 = early_reset_static_par0_go_out;
wire _guard7074 = early_reset_static_par0_go_out;
wire _guard7075 = early_reset_static_par0_go_out;
wire _guard7076 = early_reset_static_par0_go_out;
wire _guard7077 = early_reset_static_par0_go_out;
wire _guard7078 = ~_guard0;
wire _guard7079 = early_reset_static_par0_go_out;
wire _guard7080 = _guard7078 & _guard7079;
wire _guard7081 = early_reset_static_par0_go_out;
wire _guard7082 = early_reset_static_par0_go_out;
wire _guard7083 = early_reset_static_par0_go_out;
wire _guard7084 = early_reset_static_par0_go_out;
wire _guard7085 = early_reset_static_par0_go_out;
wire _guard7086 = early_reset_static_par0_go_out;
wire _guard7087 = early_reset_static_par0_go_out;
wire _guard7088 = early_reset_static_par0_go_out;
wire _guard7089 = early_reset_static_par0_go_out;
wire _guard7090 = early_reset_static_par0_go_out;
wire _guard7091 = early_reset_static_par0_go_out;
wire _guard7092 = ~_guard0;
wire _guard7093 = early_reset_static_par0_go_out;
wire _guard7094 = _guard7092 & _guard7093;
wire _guard7095 = early_reset_static_par0_go_out;
wire _guard7096 = ~_guard0;
wire _guard7097 = early_reset_static_par0_go_out;
wire _guard7098 = _guard7096 & _guard7097;
wire _guard7099 = early_reset_static_par0_go_out;
wire _guard7100 = early_reset_static_par0_go_out;
wire _guard7101 = early_reset_static_par0_go_out;
wire _guard7102 = early_reset_static_par0_go_out;
wire _guard7103 = early_reset_static_par0_go_out;
wire _guard7104 = ~_guard0;
wire _guard7105 = early_reset_static_par0_go_out;
wire _guard7106 = _guard7104 & _guard7105;
wire _guard7107 = early_reset_static_par0_go_out;
wire _guard7108 = ~_guard0;
wire _guard7109 = early_reset_static_par0_go_out;
wire _guard7110 = _guard7108 & _guard7109;
wire _guard7111 = cond_wire7_out;
wire _guard7112 = early_reset_static_par0_go_out;
wire _guard7113 = _guard7111 & _guard7112;
wire _guard7114 = cond_wire5_out;
wire _guard7115 = early_reset_static_par0_go_out;
wire _guard7116 = _guard7114 & _guard7115;
wire _guard7117 = fsm_out == 1'd0;
wire _guard7118 = cond_wire5_out;
wire _guard7119 = _guard7117 & _guard7118;
wire _guard7120 = fsm_out == 1'd0;
wire _guard7121 = _guard7119 & _guard7120;
wire _guard7122 = fsm_out == 1'd0;
wire _guard7123 = cond_wire7_out;
wire _guard7124 = _guard7122 & _guard7123;
wire _guard7125 = fsm_out == 1'd0;
wire _guard7126 = _guard7124 & _guard7125;
wire _guard7127 = _guard7121 | _guard7126;
wire _guard7128 = early_reset_static_par0_go_out;
wire _guard7129 = _guard7127 & _guard7128;
wire _guard7130 = fsm_out == 1'd0;
wire _guard7131 = cond_wire5_out;
wire _guard7132 = _guard7130 & _guard7131;
wire _guard7133 = fsm_out == 1'd0;
wire _guard7134 = _guard7132 & _guard7133;
wire _guard7135 = fsm_out == 1'd0;
wire _guard7136 = cond_wire7_out;
wire _guard7137 = _guard7135 & _guard7136;
wire _guard7138 = fsm_out == 1'd0;
wire _guard7139 = _guard7137 & _guard7138;
wire _guard7140 = _guard7134 | _guard7139;
wire _guard7141 = early_reset_static_par0_go_out;
wire _guard7142 = _guard7140 & _guard7141;
wire _guard7143 = fsm_out == 1'd0;
wire _guard7144 = cond_wire5_out;
wire _guard7145 = _guard7143 & _guard7144;
wire _guard7146 = fsm_out == 1'd0;
wire _guard7147 = _guard7145 & _guard7146;
wire _guard7148 = fsm_out == 1'd0;
wire _guard7149 = cond_wire7_out;
wire _guard7150 = _guard7148 & _guard7149;
wire _guard7151 = fsm_out == 1'd0;
wire _guard7152 = _guard7150 & _guard7151;
wire _guard7153 = _guard7147 | _guard7152;
wire _guard7154 = early_reset_static_par0_go_out;
wire _guard7155 = _guard7153 & _guard7154;
wire _guard7156 = cond_wire26_out;
wire _guard7157 = early_reset_static_par0_go_out;
wire _guard7158 = _guard7156 & _guard7157;
wire _guard7159 = cond_wire26_out;
wire _guard7160 = early_reset_static_par0_go_out;
wire _guard7161 = _guard7159 & _guard7160;
wire _guard7162 = cond_wire37_out;
wire _guard7163 = early_reset_static_par0_go_out;
wire _guard7164 = _guard7162 & _guard7163;
wire _guard7165 = cond_wire35_out;
wire _guard7166 = early_reset_static_par0_go_out;
wire _guard7167 = _guard7165 & _guard7166;
wire _guard7168 = fsm_out == 1'd0;
wire _guard7169 = cond_wire35_out;
wire _guard7170 = _guard7168 & _guard7169;
wire _guard7171 = fsm_out == 1'd0;
wire _guard7172 = _guard7170 & _guard7171;
wire _guard7173 = fsm_out == 1'd0;
wire _guard7174 = cond_wire37_out;
wire _guard7175 = _guard7173 & _guard7174;
wire _guard7176 = fsm_out == 1'd0;
wire _guard7177 = _guard7175 & _guard7176;
wire _guard7178 = _guard7172 | _guard7177;
wire _guard7179 = early_reset_static_par0_go_out;
wire _guard7180 = _guard7178 & _guard7179;
wire _guard7181 = fsm_out == 1'd0;
wire _guard7182 = cond_wire35_out;
wire _guard7183 = _guard7181 & _guard7182;
wire _guard7184 = fsm_out == 1'd0;
wire _guard7185 = _guard7183 & _guard7184;
wire _guard7186 = fsm_out == 1'd0;
wire _guard7187 = cond_wire37_out;
wire _guard7188 = _guard7186 & _guard7187;
wire _guard7189 = fsm_out == 1'd0;
wire _guard7190 = _guard7188 & _guard7189;
wire _guard7191 = _guard7185 | _guard7190;
wire _guard7192 = early_reset_static_par0_go_out;
wire _guard7193 = _guard7191 & _guard7192;
wire _guard7194 = fsm_out == 1'd0;
wire _guard7195 = cond_wire35_out;
wire _guard7196 = _guard7194 & _guard7195;
wire _guard7197 = fsm_out == 1'd0;
wire _guard7198 = _guard7196 & _guard7197;
wire _guard7199 = fsm_out == 1'd0;
wire _guard7200 = cond_wire37_out;
wire _guard7201 = _guard7199 & _guard7200;
wire _guard7202 = fsm_out == 1'd0;
wire _guard7203 = _guard7201 & _guard7202;
wire _guard7204 = _guard7198 | _guard7203;
wire _guard7205 = early_reset_static_par0_go_out;
wire _guard7206 = _guard7204 & _guard7205;
wire _guard7207 = cond_wire54_out;
wire _guard7208 = early_reset_static_par0_go_out;
wire _guard7209 = _guard7207 & _guard7208;
wire _guard7210 = cond_wire54_out;
wire _guard7211 = early_reset_static_par0_go_out;
wire _guard7212 = _guard7210 & _guard7211;
wire _guard7213 = cond_wire85_out;
wire _guard7214 = early_reset_static_par0_go_out;
wire _guard7215 = _guard7213 & _guard7214;
wire _guard7216 = cond_wire85_out;
wire _guard7217 = early_reset_static_par0_go_out;
wire _guard7218 = _guard7216 & _guard7217;
wire _guard7219 = cond_wire114_out;
wire _guard7220 = early_reset_static_par0_go_out;
wire _guard7221 = _guard7219 & _guard7220;
wire _guard7222 = cond_wire112_out;
wire _guard7223 = early_reset_static_par0_go_out;
wire _guard7224 = _guard7222 & _guard7223;
wire _guard7225 = fsm_out == 1'd0;
wire _guard7226 = cond_wire112_out;
wire _guard7227 = _guard7225 & _guard7226;
wire _guard7228 = fsm_out == 1'd0;
wire _guard7229 = _guard7227 & _guard7228;
wire _guard7230 = fsm_out == 1'd0;
wire _guard7231 = cond_wire114_out;
wire _guard7232 = _guard7230 & _guard7231;
wire _guard7233 = fsm_out == 1'd0;
wire _guard7234 = _guard7232 & _guard7233;
wire _guard7235 = _guard7229 | _guard7234;
wire _guard7236 = early_reset_static_par0_go_out;
wire _guard7237 = _guard7235 & _guard7236;
wire _guard7238 = fsm_out == 1'd0;
wire _guard7239 = cond_wire112_out;
wire _guard7240 = _guard7238 & _guard7239;
wire _guard7241 = fsm_out == 1'd0;
wire _guard7242 = _guard7240 & _guard7241;
wire _guard7243 = fsm_out == 1'd0;
wire _guard7244 = cond_wire114_out;
wire _guard7245 = _guard7243 & _guard7244;
wire _guard7246 = fsm_out == 1'd0;
wire _guard7247 = _guard7245 & _guard7246;
wire _guard7248 = _guard7242 | _guard7247;
wire _guard7249 = early_reset_static_par0_go_out;
wire _guard7250 = _guard7248 & _guard7249;
wire _guard7251 = fsm_out == 1'd0;
wire _guard7252 = cond_wire112_out;
wire _guard7253 = _guard7251 & _guard7252;
wire _guard7254 = fsm_out == 1'd0;
wire _guard7255 = _guard7253 & _guard7254;
wire _guard7256 = fsm_out == 1'd0;
wire _guard7257 = cond_wire114_out;
wire _guard7258 = _guard7256 & _guard7257;
wire _guard7259 = fsm_out == 1'd0;
wire _guard7260 = _guard7258 & _guard7259;
wire _guard7261 = _guard7255 | _guard7260;
wire _guard7262 = early_reset_static_par0_go_out;
wire _guard7263 = _guard7261 & _guard7262;
wire _guard7264 = cond_wire51_out;
wire _guard7265 = early_reset_static_par0_go_out;
wire _guard7266 = _guard7264 & _guard7265;
wire _guard7267 = cond_wire51_out;
wire _guard7268 = early_reset_static_par0_go_out;
wire _guard7269 = _guard7267 & _guard7268;
wire _guard7270 = cond_wire142_out;
wire _guard7271 = early_reset_static_par0_go_out;
wire _guard7272 = _guard7270 & _guard7271;
wire _guard7273 = cond_wire140_out;
wire _guard7274 = early_reset_static_par0_go_out;
wire _guard7275 = _guard7273 & _guard7274;
wire _guard7276 = fsm_out == 1'd0;
wire _guard7277 = cond_wire140_out;
wire _guard7278 = _guard7276 & _guard7277;
wire _guard7279 = fsm_out == 1'd0;
wire _guard7280 = _guard7278 & _guard7279;
wire _guard7281 = fsm_out == 1'd0;
wire _guard7282 = cond_wire142_out;
wire _guard7283 = _guard7281 & _guard7282;
wire _guard7284 = fsm_out == 1'd0;
wire _guard7285 = _guard7283 & _guard7284;
wire _guard7286 = _guard7280 | _guard7285;
wire _guard7287 = early_reset_static_par0_go_out;
wire _guard7288 = _guard7286 & _guard7287;
wire _guard7289 = fsm_out == 1'd0;
wire _guard7290 = cond_wire140_out;
wire _guard7291 = _guard7289 & _guard7290;
wire _guard7292 = fsm_out == 1'd0;
wire _guard7293 = _guard7291 & _guard7292;
wire _guard7294 = fsm_out == 1'd0;
wire _guard7295 = cond_wire142_out;
wire _guard7296 = _guard7294 & _guard7295;
wire _guard7297 = fsm_out == 1'd0;
wire _guard7298 = _guard7296 & _guard7297;
wire _guard7299 = _guard7293 | _guard7298;
wire _guard7300 = early_reset_static_par0_go_out;
wire _guard7301 = _guard7299 & _guard7300;
wire _guard7302 = fsm_out == 1'd0;
wire _guard7303 = cond_wire140_out;
wire _guard7304 = _guard7302 & _guard7303;
wire _guard7305 = fsm_out == 1'd0;
wire _guard7306 = _guard7304 & _guard7305;
wire _guard7307 = fsm_out == 1'd0;
wire _guard7308 = cond_wire142_out;
wire _guard7309 = _guard7307 & _guard7308;
wire _guard7310 = fsm_out == 1'd0;
wire _guard7311 = _guard7309 & _guard7310;
wire _guard7312 = _guard7306 | _guard7311;
wire _guard7313 = early_reset_static_par0_go_out;
wire _guard7314 = _guard7312 & _guard7313;
wire _guard7315 = cond_wire150_out;
wire _guard7316 = early_reset_static_par0_go_out;
wire _guard7317 = _guard7315 & _guard7316;
wire _guard7318 = cond_wire150_out;
wire _guard7319 = early_reset_static_par0_go_out;
wire _guard7320 = _guard7318 & _guard7319;
wire _guard7321 = cond_wire101_out;
wire _guard7322 = early_reset_static_par0_go_out;
wire _guard7323 = _guard7321 & _guard7322;
wire _guard7324 = cond_wire101_out;
wire _guard7325 = early_reset_static_par0_go_out;
wire _guard7326 = _guard7324 & _guard7325;
wire _guard7327 = cond_wire175_out;
wire _guard7328 = early_reset_static_par0_go_out;
wire _guard7329 = _guard7327 & _guard7328;
wire _guard7330 = cond_wire173_out;
wire _guard7331 = early_reset_static_par0_go_out;
wire _guard7332 = _guard7330 & _guard7331;
wire _guard7333 = fsm_out == 1'd0;
wire _guard7334 = cond_wire173_out;
wire _guard7335 = _guard7333 & _guard7334;
wire _guard7336 = fsm_out == 1'd0;
wire _guard7337 = _guard7335 & _guard7336;
wire _guard7338 = fsm_out == 1'd0;
wire _guard7339 = cond_wire175_out;
wire _guard7340 = _guard7338 & _guard7339;
wire _guard7341 = fsm_out == 1'd0;
wire _guard7342 = _guard7340 & _guard7341;
wire _guard7343 = _guard7337 | _guard7342;
wire _guard7344 = early_reset_static_par0_go_out;
wire _guard7345 = _guard7343 & _guard7344;
wire _guard7346 = fsm_out == 1'd0;
wire _guard7347 = cond_wire173_out;
wire _guard7348 = _guard7346 & _guard7347;
wire _guard7349 = fsm_out == 1'd0;
wire _guard7350 = _guard7348 & _guard7349;
wire _guard7351 = fsm_out == 1'd0;
wire _guard7352 = cond_wire175_out;
wire _guard7353 = _guard7351 & _guard7352;
wire _guard7354 = fsm_out == 1'd0;
wire _guard7355 = _guard7353 & _guard7354;
wire _guard7356 = _guard7350 | _guard7355;
wire _guard7357 = early_reset_static_par0_go_out;
wire _guard7358 = _guard7356 & _guard7357;
wire _guard7359 = fsm_out == 1'd0;
wire _guard7360 = cond_wire173_out;
wire _guard7361 = _guard7359 & _guard7360;
wire _guard7362 = fsm_out == 1'd0;
wire _guard7363 = _guard7361 & _guard7362;
wire _guard7364 = fsm_out == 1'd0;
wire _guard7365 = cond_wire175_out;
wire _guard7366 = _guard7364 & _guard7365;
wire _guard7367 = fsm_out == 1'd0;
wire _guard7368 = _guard7366 & _guard7367;
wire _guard7369 = _guard7363 | _guard7368;
wire _guard7370 = early_reset_static_par0_go_out;
wire _guard7371 = _guard7369 & _guard7370;
wire _guard7372 = cond_wire170_out;
wire _guard7373 = early_reset_static_par0_go_out;
wire _guard7374 = _guard7372 & _guard7373;
wire _guard7375 = cond_wire170_out;
wire _guard7376 = early_reset_static_par0_go_out;
wire _guard7377 = _guard7375 & _guard7376;
wire _guard7378 = cond_wire199_out;
wire _guard7379 = early_reset_static_par0_go_out;
wire _guard7380 = _guard7378 & _guard7379;
wire _guard7381 = cond_wire197_out;
wire _guard7382 = early_reset_static_par0_go_out;
wire _guard7383 = _guard7381 & _guard7382;
wire _guard7384 = fsm_out == 1'd0;
wire _guard7385 = cond_wire197_out;
wire _guard7386 = _guard7384 & _guard7385;
wire _guard7387 = fsm_out == 1'd0;
wire _guard7388 = _guard7386 & _guard7387;
wire _guard7389 = fsm_out == 1'd0;
wire _guard7390 = cond_wire199_out;
wire _guard7391 = _guard7389 & _guard7390;
wire _guard7392 = fsm_out == 1'd0;
wire _guard7393 = _guard7391 & _guard7392;
wire _guard7394 = _guard7388 | _guard7393;
wire _guard7395 = early_reset_static_par0_go_out;
wire _guard7396 = _guard7394 & _guard7395;
wire _guard7397 = fsm_out == 1'd0;
wire _guard7398 = cond_wire197_out;
wire _guard7399 = _guard7397 & _guard7398;
wire _guard7400 = fsm_out == 1'd0;
wire _guard7401 = _guard7399 & _guard7400;
wire _guard7402 = fsm_out == 1'd0;
wire _guard7403 = cond_wire199_out;
wire _guard7404 = _guard7402 & _guard7403;
wire _guard7405 = fsm_out == 1'd0;
wire _guard7406 = _guard7404 & _guard7405;
wire _guard7407 = _guard7401 | _guard7406;
wire _guard7408 = early_reset_static_par0_go_out;
wire _guard7409 = _guard7407 & _guard7408;
wire _guard7410 = fsm_out == 1'd0;
wire _guard7411 = cond_wire197_out;
wire _guard7412 = _guard7410 & _guard7411;
wire _guard7413 = fsm_out == 1'd0;
wire _guard7414 = _guard7412 & _guard7413;
wire _guard7415 = fsm_out == 1'd0;
wire _guard7416 = cond_wire199_out;
wire _guard7417 = _guard7415 & _guard7416;
wire _guard7418 = fsm_out == 1'd0;
wire _guard7419 = _guard7417 & _guard7418;
wire _guard7420 = _guard7414 | _guard7419;
wire _guard7421 = early_reset_static_par0_go_out;
wire _guard7422 = _guard7420 & _guard7421;
wire _guard7423 = cond_wire141_out;
wire _guard7424 = early_reset_static_par0_go_out;
wire _guard7425 = _guard7423 & _guard7424;
wire _guard7426 = cond_wire141_out;
wire _guard7427 = early_reset_static_par0_go_out;
wire _guard7428 = _guard7426 & _guard7427;
wire _guard7429 = cond_wire272_out;
wire _guard7430 = early_reset_static_par0_go_out;
wire _guard7431 = _guard7429 & _guard7430;
wire _guard7432 = cond_wire270_out;
wire _guard7433 = early_reset_static_par0_go_out;
wire _guard7434 = _guard7432 & _guard7433;
wire _guard7435 = fsm_out == 1'd0;
wire _guard7436 = cond_wire270_out;
wire _guard7437 = _guard7435 & _guard7436;
wire _guard7438 = fsm_out == 1'd0;
wire _guard7439 = _guard7437 & _guard7438;
wire _guard7440 = fsm_out == 1'd0;
wire _guard7441 = cond_wire272_out;
wire _guard7442 = _guard7440 & _guard7441;
wire _guard7443 = fsm_out == 1'd0;
wire _guard7444 = _guard7442 & _guard7443;
wire _guard7445 = _guard7439 | _guard7444;
wire _guard7446 = early_reset_static_par0_go_out;
wire _guard7447 = _guard7445 & _guard7446;
wire _guard7448 = fsm_out == 1'd0;
wire _guard7449 = cond_wire270_out;
wire _guard7450 = _guard7448 & _guard7449;
wire _guard7451 = fsm_out == 1'd0;
wire _guard7452 = _guard7450 & _guard7451;
wire _guard7453 = fsm_out == 1'd0;
wire _guard7454 = cond_wire272_out;
wire _guard7455 = _guard7453 & _guard7454;
wire _guard7456 = fsm_out == 1'd0;
wire _guard7457 = _guard7455 & _guard7456;
wire _guard7458 = _guard7452 | _guard7457;
wire _guard7459 = early_reset_static_par0_go_out;
wire _guard7460 = _guard7458 & _guard7459;
wire _guard7461 = fsm_out == 1'd0;
wire _guard7462 = cond_wire270_out;
wire _guard7463 = _guard7461 & _guard7462;
wire _guard7464 = fsm_out == 1'd0;
wire _guard7465 = _guard7463 & _guard7464;
wire _guard7466 = fsm_out == 1'd0;
wire _guard7467 = cond_wire272_out;
wire _guard7468 = _guard7466 & _guard7467;
wire _guard7469 = fsm_out == 1'd0;
wire _guard7470 = _guard7468 & _guard7469;
wire _guard7471 = _guard7465 | _guard7470;
wire _guard7472 = early_reset_static_par0_go_out;
wire _guard7473 = _guard7471 & _guard7472;
wire _guard7474 = cond_wire297_out;
wire _guard7475 = early_reset_static_par0_go_out;
wire _guard7476 = _guard7474 & _guard7475;
wire _guard7477 = cond_wire295_out;
wire _guard7478 = early_reset_static_par0_go_out;
wire _guard7479 = _guard7477 & _guard7478;
wire _guard7480 = fsm_out == 1'd0;
wire _guard7481 = cond_wire295_out;
wire _guard7482 = _guard7480 & _guard7481;
wire _guard7483 = fsm_out == 1'd0;
wire _guard7484 = _guard7482 & _guard7483;
wire _guard7485 = fsm_out == 1'd0;
wire _guard7486 = cond_wire297_out;
wire _guard7487 = _guard7485 & _guard7486;
wire _guard7488 = fsm_out == 1'd0;
wire _guard7489 = _guard7487 & _guard7488;
wire _guard7490 = _guard7484 | _guard7489;
wire _guard7491 = early_reset_static_par0_go_out;
wire _guard7492 = _guard7490 & _guard7491;
wire _guard7493 = fsm_out == 1'd0;
wire _guard7494 = cond_wire295_out;
wire _guard7495 = _guard7493 & _guard7494;
wire _guard7496 = fsm_out == 1'd0;
wire _guard7497 = _guard7495 & _guard7496;
wire _guard7498 = fsm_out == 1'd0;
wire _guard7499 = cond_wire297_out;
wire _guard7500 = _guard7498 & _guard7499;
wire _guard7501 = fsm_out == 1'd0;
wire _guard7502 = _guard7500 & _guard7501;
wire _guard7503 = _guard7497 | _guard7502;
wire _guard7504 = early_reset_static_par0_go_out;
wire _guard7505 = _guard7503 & _guard7504;
wire _guard7506 = fsm_out == 1'd0;
wire _guard7507 = cond_wire295_out;
wire _guard7508 = _guard7506 & _guard7507;
wire _guard7509 = fsm_out == 1'd0;
wire _guard7510 = _guard7508 & _guard7509;
wire _guard7511 = fsm_out == 1'd0;
wire _guard7512 = cond_wire297_out;
wire _guard7513 = _guard7511 & _guard7512;
wire _guard7514 = fsm_out == 1'd0;
wire _guard7515 = _guard7513 & _guard7514;
wire _guard7516 = _guard7510 | _guard7515;
wire _guard7517 = early_reset_static_par0_go_out;
wire _guard7518 = _guard7516 & _guard7517;
wire _guard7519 = cond_wire292_out;
wire _guard7520 = early_reset_static_par0_go_out;
wire _guard7521 = _guard7519 & _guard7520;
wire _guard7522 = cond_wire292_out;
wire _guard7523 = early_reset_static_par0_go_out;
wire _guard7524 = _guard7522 & _guard7523;
wire _guard7525 = cond_wire247_out;
wire _guard7526 = early_reset_static_par0_go_out;
wire _guard7527 = _guard7525 & _guard7526;
wire _guard7528 = cond_wire247_out;
wire _guard7529 = early_reset_static_par0_go_out;
wire _guard7530 = _guard7528 & _guard7529;
wire _guard7531 = cond_wire308_out;
wire _guard7532 = early_reset_static_par0_go_out;
wire _guard7533 = _guard7531 & _guard7532;
wire _guard7534 = cond_wire308_out;
wire _guard7535 = early_reset_static_par0_go_out;
wire _guard7536 = _guard7534 & _guard7535;
wire _guard7537 = cond_wire328_out;
wire _guard7538 = early_reset_static_par0_go_out;
wire _guard7539 = _guard7537 & _guard7538;
wire _guard7540 = cond_wire328_out;
wire _guard7541 = early_reset_static_par0_go_out;
wire _guard7542 = _guard7540 & _guard7541;
wire _guard7543 = cond_wire276_out;
wire _guard7544 = early_reset_static_par0_go_out;
wire _guard7545 = _guard7543 & _guard7544;
wire _guard7546 = cond_wire276_out;
wire _guard7547 = early_reset_static_par0_go_out;
wire _guard7548 = _guard7546 & _guard7547;
wire _guard7549 = cond_wire288_out;
wire _guard7550 = early_reset_static_par0_go_out;
wire _guard7551 = _guard7549 & _guard7550;
wire _guard7552 = cond_wire288_out;
wire _guard7553 = early_reset_static_par0_go_out;
wire _guard7554 = _guard7552 & _guard7553;
wire _guard7555 = cond_wire434_out;
wire _guard7556 = early_reset_static_par0_go_out;
wire _guard7557 = _guard7555 & _guard7556;
wire _guard7558 = cond_wire434_out;
wire _guard7559 = early_reset_static_par0_go_out;
wire _guard7560 = _guard7558 & _guard7559;
wire _guard7561 = cond_wire446_out;
wire _guard7562 = early_reset_static_par0_go_out;
wire _guard7563 = _guard7561 & _guard7562;
wire _guard7564 = cond_wire446_out;
wire _guard7565 = early_reset_static_par0_go_out;
wire _guard7566 = _guard7564 & _guard7565;
wire _guard7567 = cond_wire471_out;
wire _guard7568 = early_reset_static_par0_go_out;
wire _guard7569 = _guard7567 & _guard7568;
wire _guard7570 = cond_wire471_out;
wire _guard7571 = early_reset_static_par0_go_out;
wire _guard7572 = _guard7570 & _guard7571;
wire _guard7573 = cond_wire552_out;
wire _guard7574 = early_reset_static_par0_go_out;
wire _guard7575 = _guard7573 & _guard7574;
wire _guard7576 = cond_wire552_out;
wire _guard7577 = early_reset_static_par0_go_out;
wire _guard7578 = _guard7576 & _guard7577;
wire _guard7579 = cond_wire515_out;
wire _guard7580 = early_reset_static_par0_go_out;
wire _guard7581 = _guard7579 & _guard7580;
wire _guard7582 = cond_wire515_out;
wire _guard7583 = early_reset_static_par0_go_out;
wire _guard7584 = _guard7582 & _guard7583;
wire _guard7585 = cond_wire589_out;
wire _guard7586 = early_reset_static_par0_go_out;
wire _guard7587 = _guard7585 & _guard7586;
wire _guard7588 = cond_wire587_out;
wire _guard7589 = early_reset_static_par0_go_out;
wire _guard7590 = _guard7588 & _guard7589;
wire _guard7591 = fsm_out == 1'd0;
wire _guard7592 = cond_wire587_out;
wire _guard7593 = _guard7591 & _guard7592;
wire _guard7594 = fsm_out == 1'd0;
wire _guard7595 = _guard7593 & _guard7594;
wire _guard7596 = fsm_out == 1'd0;
wire _guard7597 = cond_wire589_out;
wire _guard7598 = _guard7596 & _guard7597;
wire _guard7599 = fsm_out == 1'd0;
wire _guard7600 = _guard7598 & _guard7599;
wire _guard7601 = _guard7595 | _guard7600;
wire _guard7602 = early_reset_static_par0_go_out;
wire _guard7603 = _guard7601 & _guard7602;
wire _guard7604 = fsm_out == 1'd0;
wire _guard7605 = cond_wire587_out;
wire _guard7606 = _guard7604 & _guard7605;
wire _guard7607 = fsm_out == 1'd0;
wire _guard7608 = _guard7606 & _guard7607;
wire _guard7609 = fsm_out == 1'd0;
wire _guard7610 = cond_wire589_out;
wire _guard7611 = _guard7609 & _guard7610;
wire _guard7612 = fsm_out == 1'd0;
wire _guard7613 = _guard7611 & _guard7612;
wire _guard7614 = _guard7608 | _guard7613;
wire _guard7615 = early_reset_static_par0_go_out;
wire _guard7616 = _guard7614 & _guard7615;
wire _guard7617 = fsm_out == 1'd0;
wire _guard7618 = cond_wire587_out;
wire _guard7619 = _guard7617 & _guard7618;
wire _guard7620 = fsm_out == 1'd0;
wire _guard7621 = _guard7619 & _guard7620;
wire _guard7622 = fsm_out == 1'd0;
wire _guard7623 = cond_wire589_out;
wire _guard7624 = _guard7622 & _guard7623;
wire _guard7625 = fsm_out == 1'd0;
wire _guard7626 = _guard7624 & _guard7625;
wire _guard7627 = _guard7621 | _guard7626;
wire _guard7628 = early_reset_static_par0_go_out;
wire _guard7629 = _guard7627 & _guard7628;
wire _guard7630 = cond_wire556_out;
wire _guard7631 = early_reset_static_par0_go_out;
wire _guard7632 = _guard7630 & _guard7631;
wire _guard7633 = cond_wire556_out;
wire _guard7634 = early_reset_static_par0_go_out;
wire _guard7635 = _guard7633 & _guard7634;
wire _guard7636 = cond_wire674_out;
wire _guard7637 = early_reset_static_par0_go_out;
wire _guard7638 = _guard7636 & _guard7637;
wire _guard7639 = cond_wire674_out;
wire _guard7640 = early_reset_static_par0_go_out;
wire _guard7641 = _guard7639 & _guard7640;
wire _guard7642 = cond_wire695_out;
wire _guard7643 = early_reset_static_par0_go_out;
wire _guard7644 = _guard7642 & _guard7643;
wire _guard7645 = cond_wire693_out;
wire _guard7646 = early_reset_static_par0_go_out;
wire _guard7647 = _guard7645 & _guard7646;
wire _guard7648 = fsm_out == 1'd0;
wire _guard7649 = cond_wire693_out;
wire _guard7650 = _guard7648 & _guard7649;
wire _guard7651 = fsm_out == 1'd0;
wire _guard7652 = _guard7650 & _guard7651;
wire _guard7653 = fsm_out == 1'd0;
wire _guard7654 = cond_wire695_out;
wire _guard7655 = _guard7653 & _guard7654;
wire _guard7656 = fsm_out == 1'd0;
wire _guard7657 = _guard7655 & _guard7656;
wire _guard7658 = _guard7652 | _guard7657;
wire _guard7659 = early_reset_static_par0_go_out;
wire _guard7660 = _guard7658 & _guard7659;
wire _guard7661 = fsm_out == 1'd0;
wire _guard7662 = cond_wire693_out;
wire _guard7663 = _guard7661 & _guard7662;
wire _guard7664 = fsm_out == 1'd0;
wire _guard7665 = _guard7663 & _guard7664;
wire _guard7666 = fsm_out == 1'd0;
wire _guard7667 = cond_wire695_out;
wire _guard7668 = _guard7666 & _guard7667;
wire _guard7669 = fsm_out == 1'd0;
wire _guard7670 = _guard7668 & _guard7669;
wire _guard7671 = _guard7665 | _guard7670;
wire _guard7672 = early_reset_static_par0_go_out;
wire _guard7673 = _guard7671 & _guard7672;
wire _guard7674 = fsm_out == 1'd0;
wire _guard7675 = cond_wire693_out;
wire _guard7676 = _guard7674 & _guard7675;
wire _guard7677 = fsm_out == 1'd0;
wire _guard7678 = _guard7676 & _guard7677;
wire _guard7679 = fsm_out == 1'd0;
wire _guard7680 = cond_wire695_out;
wire _guard7681 = _guard7679 & _guard7680;
wire _guard7682 = fsm_out == 1'd0;
wire _guard7683 = _guard7681 & _guard7682;
wire _guard7684 = _guard7678 | _guard7683;
wire _guard7685 = early_reset_static_par0_go_out;
wire _guard7686 = _guard7684 & _guard7685;
wire _guard7687 = cond_wire703_out;
wire _guard7688 = early_reset_static_par0_go_out;
wire _guard7689 = _guard7687 & _guard7688;
wire _guard7690 = cond_wire701_out;
wire _guard7691 = early_reset_static_par0_go_out;
wire _guard7692 = _guard7690 & _guard7691;
wire _guard7693 = fsm_out == 1'd0;
wire _guard7694 = cond_wire701_out;
wire _guard7695 = _guard7693 & _guard7694;
wire _guard7696 = fsm_out == 1'd0;
wire _guard7697 = _guard7695 & _guard7696;
wire _guard7698 = fsm_out == 1'd0;
wire _guard7699 = cond_wire703_out;
wire _guard7700 = _guard7698 & _guard7699;
wire _guard7701 = fsm_out == 1'd0;
wire _guard7702 = _guard7700 & _guard7701;
wire _guard7703 = _guard7697 | _guard7702;
wire _guard7704 = early_reset_static_par0_go_out;
wire _guard7705 = _guard7703 & _guard7704;
wire _guard7706 = fsm_out == 1'd0;
wire _guard7707 = cond_wire701_out;
wire _guard7708 = _guard7706 & _guard7707;
wire _guard7709 = fsm_out == 1'd0;
wire _guard7710 = _guard7708 & _guard7709;
wire _guard7711 = fsm_out == 1'd0;
wire _guard7712 = cond_wire703_out;
wire _guard7713 = _guard7711 & _guard7712;
wire _guard7714 = fsm_out == 1'd0;
wire _guard7715 = _guard7713 & _guard7714;
wire _guard7716 = _guard7710 | _guard7715;
wire _guard7717 = early_reset_static_par0_go_out;
wire _guard7718 = _guard7716 & _guard7717;
wire _guard7719 = fsm_out == 1'd0;
wire _guard7720 = cond_wire701_out;
wire _guard7721 = _guard7719 & _guard7720;
wire _guard7722 = fsm_out == 1'd0;
wire _guard7723 = _guard7721 & _guard7722;
wire _guard7724 = fsm_out == 1'd0;
wire _guard7725 = cond_wire703_out;
wire _guard7726 = _guard7724 & _guard7725;
wire _guard7727 = fsm_out == 1'd0;
wire _guard7728 = _guard7726 & _guard7727;
wire _guard7729 = _guard7723 | _guard7728;
wire _guard7730 = early_reset_static_par0_go_out;
wire _guard7731 = _guard7729 & _guard7730;
wire _guard7732 = cond_wire739_out;
wire _guard7733 = early_reset_static_par0_go_out;
wire _guard7734 = _guard7732 & _guard7733;
wire _guard7735 = cond_wire739_out;
wire _guard7736 = early_reset_static_par0_go_out;
wire _guard7737 = _guard7735 & _guard7736;
wire _guard7738 = cond_wire748_out;
wire _guard7739 = early_reset_static_par0_go_out;
wire _guard7740 = _guard7738 & _guard7739;
wire _guard7741 = cond_wire746_out;
wire _guard7742 = early_reset_static_par0_go_out;
wire _guard7743 = _guard7741 & _guard7742;
wire _guard7744 = fsm_out == 1'd0;
wire _guard7745 = cond_wire746_out;
wire _guard7746 = _guard7744 & _guard7745;
wire _guard7747 = fsm_out == 1'd0;
wire _guard7748 = _guard7746 & _guard7747;
wire _guard7749 = fsm_out == 1'd0;
wire _guard7750 = cond_wire748_out;
wire _guard7751 = _guard7749 & _guard7750;
wire _guard7752 = fsm_out == 1'd0;
wire _guard7753 = _guard7751 & _guard7752;
wire _guard7754 = _guard7748 | _guard7753;
wire _guard7755 = early_reset_static_par0_go_out;
wire _guard7756 = _guard7754 & _guard7755;
wire _guard7757 = fsm_out == 1'd0;
wire _guard7758 = cond_wire746_out;
wire _guard7759 = _guard7757 & _guard7758;
wire _guard7760 = fsm_out == 1'd0;
wire _guard7761 = _guard7759 & _guard7760;
wire _guard7762 = fsm_out == 1'd0;
wire _guard7763 = cond_wire748_out;
wire _guard7764 = _guard7762 & _guard7763;
wire _guard7765 = fsm_out == 1'd0;
wire _guard7766 = _guard7764 & _guard7765;
wire _guard7767 = _guard7761 | _guard7766;
wire _guard7768 = early_reset_static_par0_go_out;
wire _guard7769 = _guard7767 & _guard7768;
wire _guard7770 = fsm_out == 1'd0;
wire _guard7771 = cond_wire746_out;
wire _guard7772 = _guard7770 & _guard7771;
wire _guard7773 = fsm_out == 1'd0;
wire _guard7774 = _guard7772 & _guard7773;
wire _guard7775 = fsm_out == 1'd0;
wire _guard7776 = cond_wire748_out;
wire _guard7777 = _guard7775 & _guard7776;
wire _guard7778 = fsm_out == 1'd0;
wire _guard7779 = _guard7777 & _guard7778;
wire _guard7780 = _guard7774 | _guard7779;
wire _guard7781 = early_reset_static_par0_go_out;
wire _guard7782 = _guard7780 & _guard7781;
wire _guard7783 = cond_wire794_out;
wire _guard7784 = early_reset_static_par0_go_out;
wire _guard7785 = _guard7783 & _guard7784;
wire _guard7786 = cond_wire794_out;
wire _guard7787 = early_reset_static_par0_go_out;
wire _guard7788 = _guard7786 & _guard7787;
wire _guard7789 = cond_wire771_out;
wire _guard7790 = early_reset_static_par0_go_out;
wire _guard7791 = _guard7789 & _guard7790;
wire _guard7792 = cond_wire771_out;
wire _guard7793 = early_reset_static_par0_go_out;
wire _guard7794 = _guard7792 & _guard7793;
wire _guard7795 = cond_wire848_out;
wire _guard7796 = early_reset_static_par0_go_out;
wire _guard7797 = _guard7795 & _guard7796;
wire _guard7798 = cond_wire848_out;
wire _guard7799 = early_reset_static_par0_go_out;
wire _guard7800 = _guard7798 & _guard7799;
wire _guard7801 = cond_wire890_out;
wire _guard7802 = early_reset_static_par0_go_out;
wire _guard7803 = _guard7801 & _guard7802;
wire _guard7804 = cond_wire888_out;
wire _guard7805 = early_reset_static_par0_go_out;
wire _guard7806 = _guard7804 & _guard7805;
wire _guard7807 = fsm_out == 1'd0;
wire _guard7808 = cond_wire888_out;
wire _guard7809 = _guard7807 & _guard7808;
wire _guard7810 = fsm_out == 1'd0;
wire _guard7811 = _guard7809 & _guard7810;
wire _guard7812 = fsm_out == 1'd0;
wire _guard7813 = cond_wire890_out;
wire _guard7814 = _guard7812 & _guard7813;
wire _guard7815 = fsm_out == 1'd0;
wire _guard7816 = _guard7814 & _guard7815;
wire _guard7817 = _guard7811 | _guard7816;
wire _guard7818 = early_reset_static_par0_go_out;
wire _guard7819 = _guard7817 & _guard7818;
wire _guard7820 = fsm_out == 1'd0;
wire _guard7821 = cond_wire888_out;
wire _guard7822 = _guard7820 & _guard7821;
wire _guard7823 = fsm_out == 1'd0;
wire _guard7824 = _guard7822 & _guard7823;
wire _guard7825 = fsm_out == 1'd0;
wire _guard7826 = cond_wire890_out;
wire _guard7827 = _guard7825 & _guard7826;
wire _guard7828 = fsm_out == 1'd0;
wire _guard7829 = _guard7827 & _guard7828;
wire _guard7830 = _guard7824 | _guard7829;
wire _guard7831 = early_reset_static_par0_go_out;
wire _guard7832 = _guard7830 & _guard7831;
wire _guard7833 = fsm_out == 1'd0;
wire _guard7834 = cond_wire888_out;
wire _guard7835 = _guard7833 & _guard7834;
wire _guard7836 = fsm_out == 1'd0;
wire _guard7837 = _guard7835 & _guard7836;
wire _guard7838 = fsm_out == 1'd0;
wire _guard7839 = cond_wire890_out;
wire _guard7840 = _guard7838 & _guard7839;
wire _guard7841 = fsm_out == 1'd0;
wire _guard7842 = _guard7840 & _guard7841;
wire _guard7843 = _guard7837 | _guard7842;
wire _guard7844 = early_reset_static_par0_go_out;
wire _guard7845 = _guard7843 & _guard7844;
wire _guard7846 = cond_wire897_out;
wire _guard7847 = early_reset_static_par0_go_out;
wire _guard7848 = _guard7846 & _guard7847;
wire _guard7849 = cond_wire897_out;
wire _guard7850 = early_reset_static_par0_go_out;
wire _guard7851 = _guard7849 & _guard7850;
wire _guard7852 = cond_wire901_out;
wire _guard7853 = early_reset_static_par0_go_out;
wire _guard7854 = _guard7852 & _guard7853;
wire _guard7855 = cond_wire901_out;
wire _guard7856 = early_reset_static_par0_go_out;
wire _guard7857 = _guard7855 & _guard7856;
wire _guard7858 = cond_wire917_out;
wire _guard7859 = early_reset_static_par0_go_out;
wire _guard7860 = _guard7858 & _guard7859;
wire _guard7861 = cond_wire917_out;
wire _guard7862 = early_reset_static_par0_go_out;
wire _guard7863 = _guard7861 & _guard7862;
wire _guard7864 = cond_wire926_out;
wire _guard7865 = early_reset_static_par0_go_out;
wire _guard7866 = _guard7864 & _guard7865;
wire _guard7867 = cond_wire926_out;
wire _guard7868 = early_reset_static_par0_go_out;
wire _guard7869 = _guard7867 & _guard7868;
wire _guard7870 = cond_wire877_out;
wire _guard7871 = early_reset_static_par0_go_out;
wire _guard7872 = _guard7870 & _guard7871;
wire _guard7873 = cond_wire877_out;
wire _guard7874 = early_reset_static_par0_go_out;
wire _guard7875 = _guard7873 & _guard7874;
wire _guard7876 = cond_wire950_out;
wire _guard7877 = early_reset_static_par0_go_out;
wire _guard7878 = _guard7876 & _guard7877;
wire _guard7879 = cond_wire950_out;
wire _guard7880 = early_reset_static_par0_go_out;
wire _guard7881 = _guard7879 & _guard7880;
wire _guard7882 = cond_wire966_out;
wire _guard7883 = early_reset_static_par0_go_out;
wire _guard7884 = _guard7882 & _guard7883;
wire _guard7885 = cond_wire966_out;
wire _guard7886 = early_reset_static_par0_go_out;
wire _guard7887 = _guard7885 & _guard7886;
wire _guard7888 = cond_wire1023_out;
wire _guard7889 = early_reset_static_par0_go_out;
wire _guard7890 = _guard7888 & _guard7889;
wire _guard7891 = cond_wire1023_out;
wire _guard7892 = early_reset_static_par0_go_out;
wire _guard7893 = _guard7891 & _guard7892;
wire _guard7894 = cond_wire1031_out;
wire _guard7895 = early_reset_static_par0_go_out;
wire _guard7896 = _guard7894 & _guard7895;
wire _guard7897 = cond_wire1031_out;
wire _guard7898 = early_reset_static_par0_go_out;
wire _guard7899 = _guard7897 & _guard7898;
wire _guard7900 = cond_wire1048_out;
wire _guard7901 = early_reset_static_par0_go_out;
wire _guard7902 = _guard7900 & _guard7901;
wire _guard7903 = cond_wire1046_out;
wire _guard7904 = early_reset_static_par0_go_out;
wire _guard7905 = _guard7903 & _guard7904;
wire _guard7906 = fsm_out == 1'd0;
wire _guard7907 = cond_wire1046_out;
wire _guard7908 = _guard7906 & _guard7907;
wire _guard7909 = fsm_out == 1'd0;
wire _guard7910 = _guard7908 & _guard7909;
wire _guard7911 = fsm_out == 1'd0;
wire _guard7912 = cond_wire1048_out;
wire _guard7913 = _guard7911 & _guard7912;
wire _guard7914 = fsm_out == 1'd0;
wire _guard7915 = _guard7913 & _guard7914;
wire _guard7916 = _guard7910 | _guard7915;
wire _guard7917 = early_reset_static_par0_go_out;
wire _guard7918 = _guard7916 & _guard7917;
wire _guard7919 = fsm_out == 1'd0;
wire _guard7920 = cond_wire1046_out;
wire _guard7921 = _guard7919 & _guard7920;
wire _guard7922 = fsm_out == 1'd0;
wire _guard7923 = _guard7921 & _guard7922;
wire _guard7924 = fsm_out == 1'd0;
wire _guard7925 = cond_wire1048_out;
wire _guard7926 = _guard7924 & _guard7925;
wire _guard7927 = fsm_out == 1'd0;
wire _guard7928 = _guard7926 & _guard7927;
wire _guard7929 = _guard7923 | _guard7928;
wire _guard7930 = early_reset_static_par0_go_out;
wire _guard7931 = _guard7929 & _guard7930;
wire _guard7932 = fsm_out == 1'd0;
wire _guard7933 = cond_wire1046_out;
wire _guard7934 = _guard7932 & _guard7933;
wire _guard7935 = fsm_out == 1'd0;
wire _guard7936 = _guard7934 & _guard7935;
wire _guard7937 = fsm_out == 1'd0;
wire _guard7938 = cond_wire1048_out;
wire _guard7939 = _guard7937 & _guard7938;
wire _guard7940 = fsm_out == 1'd0;
wire _guard7941 = _guard7939 & _guard7940;
wire _guard7942 = _guard7936 | _guard7941;
wire _guard7943 = early_reset_static_par0_go_out;
wire _guard7944 = _guard7942 & _guard7943;
wire _guard7945 = fsm0_out == 6'd0;
wire _guard7946 = early_reset_static_seq_go_out;
wire _guard7947 = _guard7945 & _guard7946;
wire _guard7948 = cond_wire49_out;
wire _guard7949 = early_reset_static_par0_go_out;
wire _guard7950 = _guard7948 & _guard7949;
wire _guard7951 = _guard7947 | _guard7950;
wire _guard7952 = fsm0_out == 6'd0;
wire _guard7953 = early_reset_static_seq_go_out;
wire _guard7954 = _guard7952 & _guard7953;
wire _guard7955 = cond_wire49_out;
wire _guard7956 = early_reset_static_par0_go_out;
wire _guard7957 = _guard7955 & _guard7956;
wire _guard7958 = cond_wire209_out;
wire _guard7959 = early_reset_static_par0_go_out;
wire _guard7960 = _guard7958 & _guard7959;
wire _guard7961 = cond_wire209_out;
wire _guard7962 = early_reset_static_par0_go_out;
wire _guard7963 = _guard7961 & _guard7962;
wire _guard7964 = cond_wire989_out;
wire _guard7965 = early_reset_static_par0_go_out;
wire _guard7966 = _guard7964 & _guard7965;
wire _guard7967 = cond_wire989_out;
wire _guard7968 = early_reset_static_par0_go_out;
wire _guard7969 = _guard7967 & _guard7968;
wire _guard7970 = early_reset_static_par0_go_out;
wire _guard7971 = early_reset_static_par0_go_out;
wire _guard7972 = early_reset_static_par0_go_out;
wire _guard7973 = early_reset_static_par0_go_out;
wire _guard7974 = early_reset_static_par0_go_out;
wire _guard7975 = early_reset_static_par0_go_out;
wire _guard7976 = early_reset_static_par0_go_out;
wire _guard7977 = early_reset_static_par0_go_out;
wire _guard7978 = early_reset_static_par0_go_out;
wire _guard7979 = early_reset_static_par0_go_out;
wire _guard7980 = fsm0_out == 6'd0;
wire _guard7981 = early_reset_static_seq_go_out;
wire _guard7982 = _guard7980 & _guard7981;
wire _guard7983 = early_reset_static_par0_go_out;
wire _guard7984 = _guard7982 | _guard7983;
wire _guard7985 = fsm0_out == 6'd0;
wire _guard7986 = early_reset_static_seq_go_out;
wire _guard7987 = _guard7985 & _guard7986;
wire _guard7988 = early_reset_static_par0_go_out;
wire _guard7989 = early_reset_static_par0_go_out;
wire _guard7990 = early_reset_static_par0_go_out;
wire _guard7991 = early_reset_static_par0_go_out;
wire _guard7992 = early_reset_static_par0_go_out;
wire _guard7993 = early_reset_static_par0_go_out;
wire _guard7994 = early_reset_static_par0_go_out;
wire _guard7995 = early_reset_static_par0_go_out;
wire _guard7996 = early_reset_static_par0_go_out;
wire _guard7997 = fsm0_out == 6'd0;
wire _guard7998 = early_reset_static_seq_go_out;
wire _guard7999 = _guard7997 & _guard7998;
wire _guard8000 = early_reset_static_par0_go_out;
wire _guard8001 = _guard7999 | _guard8000;
wire _guard8002 = fsm0_out == 6'd0;
wire _guard8003 = early_reset_static_seq_go_out;
wire _guard8004 = _guard8002 & _guard8003;
wire _guard8005 = early_reset_static_par0_go_out;
wire _guard8006 = early_reset_static_par0_go_out;
wire _guard8007 = early_reset_static_par0_go_out;
wire _guard8008 = early_reset_static_par0_go_out;
wire _guard8009 = early_reset_static_par0_go_out;
wire _guard8010 = fsm0_out == 6'd0;
wire _guard8011 = early_reset_static_seq_go_out;
wire _guard8012 = _guard8010 & _guard8011;
wire _guard8013 = early_reset_static_par0_go_out;
wire _guard8014 = _guard8012 | _guard8013;
wire _guard8015 = early_reset_static_par0_go_out;
wire _guard8016 = fsm0_out == 6'd0;
wire _guard8017 = early_reset_static_seq_go_out;
wire _guard8018 = _guard8016 & _guard8017;
wire _guard8019 = early_reset_static_par0_go_out;
wire _guard8020 = early_reset_static_par0_go_out;
wire _guard8021 = early_reset_static_par0_go_out;
wire _guard8022 = early_reset_static_par0_go_out;
wire _guard8023 = early_reset_static_par0_go_out;
wire _guard8024 = early_reset_static_par0_go_out;
wire _guard8025 = early_reset_static_par0_go_out;
wire _guard8026 = early_reset_static_par0_go_out;
wire _guard8027 = early_reset_static_par0_go_out;
wire _guard8028 = early_reset_static_par0_go_out;
wire _guard8029 = early_reset_static_par0_go_out;
wire _guard8030 = early_reset_static_par0_go_out;
wire _guard8031 = early_reset_static_par0_go_out;
wire _guard8032 = ~_guard0;
wire _guard8033 = early_reset_static_par0_go_out;
wire _guard8034 = _guard8032 & _guard8033;
wire _guard8035 = early_reset_static_par0_go_out;
wire _guard8036 = early_reset_static_par0_go_out;
wire _guard8037 = ~_guard0;
wire _guard8038 = early_reset_static_par0_go_out;
wire _guard8039 = _guard8037 & _guard8038;
wire _guard8040 = early_reset_static_par0_go_out;
wire _guard8041 = ~_guard0;
wire _guard8042 = early_reset_static_par0_go_out;
wire _guard8043 = _guard8041 & _guard8042;
wire _guard8044 = early_reset_static_par0_go_out;
wire _guard8045 = ~_guard0;
wire _guard8046 = early_reset_static_par0_go_out;
wire _guard8047 = _guard8045 & _guard8046;
wire _guard8048 = early_reset_static_par0_go_out;
wire _guard8049 = early_reset_static_par0_go_out;
wire _guard8050 = early_reset_static_par0_go_out;
wire _guard8051 = early_reset_static_par0_go_out;
wire _guard8052 = early_reset_static_par0_go_out;
wire _guard8053 = early_reset_static_par0_go_out;
wire _guard8054 = early_reset_static_par0_go_out;
wire _guard8055 = early_reset_static_par0_go_out;
wire _guard8056 = early_reset_static_par0_go_out;
wire _guard8057 = early_reset_static_par0_go_out;
wire _guard8058 = ~_guard0;
wire _guard8059 = early_reset_static_par0_go_out;
wire _guard8060 = _guard8058 & _guard8059;
wire _guard8061 = early_reset_static_par0_go_out;
wire _guard8062 = early_reset_static_par0_go_out;
wire _guard8063 = ~_guard0;
wire _guard8064 = early_reset_static_par0_go_out;
wire _guard8065 = _guard8063 & _guard8064;
wire _guard8066 = early_reset_static_par0_go_out;
wire _guard8067 = ~_guard0;
wire _guard8068 = early_reset_static_par0_go_out;
wire _guard8069 = _guard8067 & _guard8068;
wire _guard8070 = early_reset_static_par0_go_out;
wire _guard8071 = early_reset_static_par0_go_out;
wire _guard8072 = ~_guard0;
wire _guard8073 = early_reset_static_par0_go_out;
wire _guard8074 = _guard8072 & _guard8073;
wire _guard8075 = early_reset_static_par0_go_out;
wire _guard8076 = ~_guard0;
wire _guard8077 = early_reset_static_par0_go_out;
wire _guard8078 = _guard8076 & _guard8077;
wire _guard8079 = early_reset_static_par0_go_out;
wire _guard8080 = early_reset_static_par0_go_out;
wire _guard8081 = early_reset_static_par0_go_out;
wire _guard8082 = ~_guard0;
wire _guard8083 = early_reset_static_par0_go_out;
wire _guard8084 = _guard8082 & _guard8083;
wire _guard8085 = early_reset_static_par0_go_out;
wire _guard8086 = ~_guard0;
wire _guard8087 = early_reset_static_par0_go_out;
wire _guard8088 = _guard8086 & _guard8087;
wire _guard8089 = ~_guard0;
wire _guard8090 = early_reset_static_par0_go_out;
wire _guard8091 = _guard8089 & _guard8090;
wire _guard8092 = early_reset_static_par0_go_out;
wire _guard8093 = early_reset_static_par0_go_out;
wire _guard8094 = early_reset_static_par0_go_out;
wire _guard8095 = early_reset_static_par0_go_out;
wire _guard8096 = early_reset_static_par0_go_out;
wire _guard8097 = early_reset_static_par0_go_out;
wire _guard8098 = early_reset_static_par0_go_out;
wire _guard8099 = early_reset_static_par0_go_out;
wire _guard8100 = ~_guard0;
wire _guard8101 = early_reset_static_par0_go_out;
wire _guard8102 = _guard8100 & _guard8101;
wire _guard8103 = ~_guard0;
wire _guard8104 = early_reset_static_par0_go_out;
wire _guard8105 = _guard8103 & _guard8104;
wire _guard8106 = early_reset_static_par0_go_out;
wire _guard8107 = early_reset_static_par0_go_out;
wire _guard8108 = early_reset_static_par0_go_out;
wire _guard8109 = early_reset_static_par0_go_out;
wire _guard8110 = early_reset_static_par0_go_out;
wire _guard8111 = ~_guard0;
wire _guard8112 = early_reset_static_par0_go_out;
wire _guard8113 = _guard8111 & _guard8112;
wire _guard8114 = early_reset_static_par0_go_out;
wire _guard8115 = early_reset_static_par0_go_out;
wire _guard8116 = early_reset_static_par0_go_out;
wire _guard8117 = early_reset_static_par0_go_out;
wire _guard8118 = ~_guard0;
wire _guard8119 = early_reset_static_par0_go_out;
wire _guard8120 = _guard8118 & _guard8119;
wire _guard8121 = early_reset_static_par0_go_out;
wire _guard8122 = early_reset_static_par0_go_out;
wire _guard8123 = early_reset_static_par0_go_out;
wire _guard8124 = early_reset_static_par0_go_out;
wire _guard8125 = early_reset_static_par0_go_out;
wire _guard8126 = ~_guard0;
wire _guard8127 = early_reset_static_par0_go_out;
wire _guard8128 = _guard8126 & _guard8127;
wire _guard8129 = early_reset_static_par0_go_out;
wire _guard8130 = early_reset_static_par0_go_out;
wire _guard8131 = ~_guard0;
wire _guard8132 = early_reset_static_par0_go_out;
wire _guard8133 = _guard8131 & _guard8132;
wire _guard8134 = early_reset_static_par0_go_out;
wire _guard8135 = early_reset_static_par0_go_out;
wire _guard8136 = early_reset_static_par0_go_out;
wire _guard8137 = early_reset_static_par0_go_out;
wire _guard8138 = ~_guard0;
wire _guard8139 = early_reset_static_par0_go_out;
wire _guard8140 = _guard8138 & _guard8139;
wire _guard8141 = early_reset_static_par0_go_out;
wire _guard8142 = early_reset_static_par0_go_out;
wire _guard8143 = early_reset_static_par0_go_out;
wire _guard8144 = ~_guard0;
wire _guard8145 = early_reset_static_par0_go_out;
wire _guard8146 = _guard8144 & _guard8145;
wire _guard8147 = early_reset_static_par0_go_out;
wire _guard8148 = ~_guard0;
wire _guard8149 = early_reset_static_par0_go_out;
wire _guard8150 = _guard8148 & _guard8149;
wire _guard8151 = early_reset_static_par0_go_out;
wire _guard8152 = early_reset_static_par0_go_out;
wire _guard8153 = ~_guard0;
wire _guard8154 = early_reset_static_par0_go_out;
wire _guard8155 = _guard8153 & _guard8154;
wire _guard8156 = early_reset_static_par0_go_out;
wire _guard8157 = early_reset_static_par0_go_out;
wire _guard8158 = early_reset_static_par0_go_out;
wire _guard8159 = early_reset_static_par0_go_out;
wire _guard8160 = early_reset_static_par0_go_out;
wire _guard8161 = early_reset_static_par0_go_out;
wire _guard8162 = early_reset_static_par0_go_out;
wire _guard8163 = early_reset_static_par0_go_out;
wire _guard8164 = early_reset_static_par0_go_out;
wire _guard8165 = early_reset_static_par0_go_out;
wire _guard8166 = early_reset_static_par0_go_out;
wire _guard8167 = ~_guard0;
wire _guard8168 = early_reset_static_par0_go_out;
wire _guard8169 = _guard8167 & _guard8168;
wire _guard8170 = early_reset_static_par0_go_out;
wire _guard8171 = ~_guard0;
wire _guard8172 = early_reset_static_par0_go_out;
wire _guard8173 = _guard8171 & _guard8172;
wire _guard8174 = early_reset_static_par0_go_out;
wire _guard8175 = early_reset_static_par0_go_out;
wire _guard8176 = early_reset_static_par0_go_out;
wire _guard8177 = early_reset_static_par0_go_out;
wire _guard8178 = early_reset_static_par0_go_out;
wire _guard8179 = early_reset_static_par0_go_out;
wire _guard8180 = early_reset_static_par0_go_out;
wire _guard8181 = early_reset_static_par0_go_out;
wire _guard8182 = early_reset_static_par0_go_out;
wire _guard8183 = early_reset_static_par0_go_out;
wire _guard8184 = ~_guard0;
wire _guard8185 = early_reset_static_par0_go_out;
wire _guard8186 = _guard8184 & _guard8185;
wire _guard8187 = early_reset_static_par0_go_out;
wire _guard8188 = ~_guard0;
wire _guard8189 = early_reset_static_par0_go_out;
wire _guard8190 = _guard8188 & _guard8189;
wire _guard8191 = ~_guard0;
wire _guard8192 = early_reset_static_par0_go_out;
wire _guard8193 = _guard8191 & _guard8192;
wire _guard8194 = early_reset_static_par0_go_out;
wire _guard8195 = early_reset_static_par0_go_out;
wire _guard8196 = ~_guard0;
wire _guard8197 = early_reset_static_par0_go_out;
wire _guard8198 = _guard8196 & _guard8197;
wire _guard8199 = ~_guard0;
wire _guard8200 = early_reset_static_par0_go_out;
wire _guard8201 = _guard8199 & _guard8200;
wire _guard8202 = early_reset_static_par0_go_out;
wire _guard8203 = early_reset_static_par0_go_out;
wire _guard8204 = early_reset_static_par0_go_out;
wire _guard8205 = ~_guard0;
wire _guard8206 = early_reset_static_par0_go_out;
wire _guard8207 = _guard8205 & _guard8206;
wire _guard8208 = early_reset_static_par0_go_out;
wire _guard8209 = early_reset_static_par0_go_out;
wire _guard8210 = early_reset_static_par0_go_out;
wire _guard8211 = early_reset_static_par0_go_out;
wire _guard8212 = early_reset_static_par0_go_out;
wire _guard8213 = ~_guard0;
wire _guard8214 = early_reset_static_par0_go_out;
wire _guard8215 = _guard8213 & _guard8214;
wire _guard8216 = early_reset_static_par0_go_out;
wire _guard8217 = early_reset_static_par0_go_out;
wire _guard8218 = early_reset_static_par0_go_out;
wire _guard8219 = early_reset_static_par0_go_out;
wire _guard8220 = early_reset_static_par0_go_out;
wire _guard8221 = early_reset_static_par0_go_out;
wire _guard8222 = early_reset_static_par0_go_out;
wire _guard8223 = ~_guard0;
wire _guard8224 = early_reset_static_par0_go_out;
wire _guard8225 = _guard8223 & _guard8224;
wire _guard8226 = early_reset_static_par0_go_out;
wire _guard8227 = early_reset_static_par0_go_out;
wire _guard8228 = early_reset_static_par0_go_out;
wire _guard8229 = early_reset_static_par0_go_out;
wire _guard8230 = ~_guard0;
wire _guard8231 = early_reset_static_par0_go_out;
wire _guard8232 = _guard8230 & _guard8231;
wire _guard8233 = early_reset_static_par0_go_out;
wire _guard8234 = early_reset_static_par0_go_out;
wire _guard8235 = early_reset_static_par0_go_out;
wire _guard8236 = ~_guard0;
wire _guard8237 = early_reset_static_par0_go_out;
wire _guard8238 = _guard8236 & _guard8237;
wire _guard8239 = ~_guard0;
wire _guard8240 = early_reset_static_par0_go_out;
wire _guard8241 = _guard8239 & _guard8240;
wire _guard8242 = early_reset_static_par0_go_out;
wire _guard8243 = early_reset_static_par0_go_out;
wire _guard8244 = early_reset_static_par0_go_out;
wire _guard8245 = early_reset_static_par0_go_out;
wire _guard8246 = ~_guard0;
wire _guard8247 = early_reset_static_par0_go_out;
wire _guard8248 = _guard8246 & _guard8247;
wire _guard8249 = ~_guard0;
wire _guard8250 = early_reset_static_par0_go_out;
wire _guard8251 = _guard8249 & _guard8250;
wire _guard8252 = early_reset_static_par0_go_out;
wire _guard8253 = early_reset_static_par0_go_out;
wire _guard8254 = ~_guard0;
wire _guard8255 = early_reset_static_par0_go_out;
wire _guard8256 = _guard8254 & _guard8255;
wire _guard8257 = early_reset_static_par0_go_out;
wire _guard8258 = early_reset_static_par0_go_out;
wire _guard8259 = ~_guard0;
wire _guard8260 = early_reset_static_par0_go_out;
wire _guard8261 = _guard8259 & _guard8260;
wire _guard8262 = early_reset_static_par0_go_out;
wire _guard8263 = ~_guard0;
wire _guard8264 = early_reset_static_par0_go_out;
wire _guard8265 = _guard8263 & _guard8264;
wire _guard8266 = early_reset_static_par0_go_out;
wire _guard8267 = early_reset_static_par0_go_out;
wire _guard8268 = early_reset_static_par0_go_out;
wire _guard8269 = early_reset_static_par0_go_out;
wire _guard8270 = early_reset_static_par0_go_out;
wire _guard8271 = early_reset_static_par0_go_out;
wire _guard8272 = early_reset_static_par0_go_out;
wire _guard8273 = early_reset_static_par0_go_out;
wire _guard8274 = early_reset_static_par0_go_out;
wire _guard8275 = early_reset_static_par0_go_out;
wire _guard8276 = ~_guard0;
wire _guard8277 = early_reset_static_par0_go_out;
wire _guard8278 = _guard8276 & _guard8277;
wire _guard8279 = early_reset_static_par0_go_out;
wire _guard8280 = early_reset_static_par0_go_out;
wire _guard8281 = early_reset_static_par0_go_out;
wire _guard8282 = early_reset_static_par0_go_out;
wire _guard8283 = early_reset_static_par0_go_out;
wire _guard8284 = early_reset_static_par0_go_out;
wire _guard8285 = early_reset_static_par0_go_out;
wire _guard8286 = early_reset_static_par0_go_out;
wire _guard8287 = early_reset_static_par0_go_out;
wire _guard8288 = early_reset_static_par0_go_out;
wire _guard8289 = early_reset_static_par0_go_out;
wire _guard8290 = early_reset_static_par0_go_out;
wire _guard8291 = early_reset_static_par0_go_out;
wire _guard8292 = early_reset_static_par0_go_out;
wire _guard8293 = early_reset_static_par0_go_out;
wire _guard8294 = early_reset_static_par0_go_out;
wire _guard8295 = early_reset_static_par0_go_out;
wire _guard8296 = early_reset_static_par0_go_out;
wire _guard8297 = early_reset_static_par0_go_out;
wire _guard8298 = ~_guard0;
wire _guard8299 = early_reset_static_par0_go_out;
wire _guard8300 = _guard8298 & _guard8299;
wire _guard8301 = early_reset_static_par0_go_out;
wire _guard8302 = early_reset_static_par0_go_out;
wire _guard8303 = ~_guard0;
wire _guard8304 = early_reset_static_par0_go_out;
wire _guard8305 = _guard8303 & _guard8304;
wire _guard8306 = early_reset_static_par0_go_out;
wire _guard8307 = ~_guard0;
wire _guard8308 = early_reset_static_par0_go_out;
wire _guard8309 = _guard8307 & _guard8308;
wire _guard8310 = early_reset_static_par0_go_out;
wire _guard8311 = early_reset_static_par0_go_out;
wire _guard8312 = early_reset_static_par0_go_out;
wire _guard8313 = early_reset_static_par0_go_out;
wire _guard8314 = ~_guard0;
wire _guard8315 = early_reset_static_par0_go_out;
wire _guard8316 = _guard8314 & _guard8315;
wire _guard8317 = early_reset_static_par0_go_out;
wire _guard8318 = early_reset_static_par0_go_out;
wire _guard8319 = early_reset_static_par0_go_out;
wire _guard8320 = ~_guard0;
wire _guard8321 = early_reset_static_par0_go_out;
wire _guard8322 = _guard8320 & _guard8321;
wire _guard8323 = early_reset_static_par0_go_out;
wire _guard8324 = early_reset_static_par0_go_out;
wire _guard8325 = early_reset_static_par0_go_out;
wire _guard8326 = early_reset_static_par0_go_out;
wire _guard8327 = early_reset_static_par0_go_out;
wire _guard8328 = early_reset_static_par0_go_out;
wire _guard8329 = early_reset_static_par0_go_out;
wire _guard8330 = early_reset_static_par0_go_out;
wire _guard8331 = early_reset_static_par0_go_out;
wire _guard8332 = early_reset_static_par0_go_out;
wire _guard8333 = early_reset_static_par0_go_out;
wire _guard8334 = early_reset_static_par0_go_out;
wire _guard8335 = early_reset_static_par0_go_out;
wire _guard8336 = early_reset_static_par0_go_out;
wire _guard8337 = early_reset_static_par0_go_out;
wire _guard8338 = early_reset_static_par0_go_out;
wire _guard8339 = ~_guard0;
wire _guard8340 = early_reset_static_par0_go_out;
wire _guard8341 = _guard8339 & _guard8340;
wire _guard8342 = early_reset_static_par0_go_out;
wire _guard8343 = early_reset_static_par0_go_out;
wire _guard8344 = ~_guard0;
wire _guard8345 = early_reset_static_par0_go_out;
wire _guard8346 = _guard8344 & _guard8345;
wire _guard8347 = early_reset_static_par0_go_out;
wire _guard8348 = ~_guard0;
wire _guard8349 = early_reset_static_par0_go_out;
wire _guard8350 = _guard8348 & _guard8349;
wire _guard8351 = early_reset_static_par0_go_out;
wire _guard8352 = early_reset_static_par0_go_out;
wire _guard8353 = early_reset_static_par0_go_out;
wire _guard8354 = early_reset_static_par0_go_out;
wire _guard8355 = early_reset_static_par0_go_out;
wire _guard8356 = ~_guard0;
wire _guard8357 = early_reset_static_par0_go_out;
wire _guard8358 = _guard8356 & _guard8357;
wire _guard8359 = ~_guard0;
wire _guard8360 = early_reset_static_par0_go_out;
wire _guard8361 = _guard8359 & _guard8360;
wire _guard8362 = early_reset_static_par0_go_out;
wire _guard8363 = ~_guard0;
wire _guard8364 = early_reset_static_par0_go_out;
wire _guard8365 = _guard8363 & _guard8364;
wire _guard8366 = early_reset_static_par0_go_out;
wire _guard8367 = ~_guard0;
wire _guard8368 = early_reset_static_par0_go_out;
wire _guard8369 = _guard8367 & _guard8368;
wire _guard8370 = early_reset_static_par0_go_out;
wire _guard8371 = early_reset_static_par0_go_out;
wire _guard8372 = early_reset_static_par0_go_out;
wire _guard8373 = early_reset_static_par0_go_out;
wire _guard8374 = early_reset_static_par0_go_out;
wire _guard8375 = early_reset_static_par0_go_out;
wire _guard8376 = early_reset_static_par0_go_out;
wire _guard8377 = early_reset_static_par0_go_out;
wire _guard8378 = early_reset_static_par0_go_out;
wire _guard8379 = early_reset_static_par0_go_out;
wire _guard8380 = ~_guard0;
wire _guard8381 = early_reset_static_par0_go_out;
wire _guard8382 = _guard8380 & _guard8381;
wire _guard8383 = ~_guard0;
wire _guard8384 = early_reset_static_par0_go_out;
wire _guard8385 = _guard8383 & _guard8384;
wire _guard8386 = early_reset_static_par0_go_out;
wire _guard8387 = early_reset_static_par0_go_out;
wire _guard8388 = early_reset_static_par0_go_out;
wire _guard8389 = early_reset_static_par0_go_out;
wire _guard8390 = early_reset_static_par0_go_out;
wire _guard8391 = early_reset_static_par0_go_out;
wire _guard8392 = ~_guard0;
wire _guard8393 = early_reset_static_par0_go_out;
wire _guard8394 = _guard8392 & _guard8393;
wire _guard8395 = cond_wire56_out;
wire _guard8396 = early_reset_static_par0_go_out;
wire _guard8397 = _guard8395 & _guard8396;
wire _guard8398 = cond_wire56_out;
wire _guard8399 = early_reset_static_par0_go_out;
wire _guard8400 = _guard8398 & _guard8399;
wire _guard8401 = cond_wire82_out;
wire _guard8402 = early_reset_static_par0_go_out;
wire _guard8403 = _guard8401 & _guard8402;
wire _guard8404 = cond_wire80_out;
wire _guard8405 = early_reset_static_par0_go_out;
wire _guard8406 = _guard8404 & _guard8405;
wire _guard8407 = fsm_out == 1'd0;
wire _guard8408 = cond_wire80_out;
wire _guard8409 = _guard8407 & _guard8408;
wire _guard8410 = fsm_out == 1'd0;
wire _guard8411 = _guard8409 & _guard8410;
wire _guard8412 = fsm_out == 1'd0;
wire _guard8413 = cond_wire82_out;
wire _guard8414 = _guard8412 & _guard8413;
wire _guard8415 = fsm_out == 1'd0;
wire _guard8416 = _guard8414 & _guard8415;
wire _guard8417 = _guard8411 | _guard8416;
wire _guard8418 = early_reset_static_par0_go_out;
wire _guard8419 = _guard8417 & _guard8418;
wire _guard8420 = fsm_out == 1'd0;
wire _guard8421 = cond_wire80_out;
wire _guard8422 = _guard8420 & _guard8421;
wire _guard8423 = fsm_out == 1'd0;
wire _guard8424 = _guard8422 & _guard8423;
wire _guard8425 = fsm_out == 1'd0;
wire _guard8426 = cond_wire82_out;
wire _guard8427 = _guard8425 & _guard8426;
wire _guard8428 = fsm_out == 1'd0;
wire _guard8429 = _guard8427 & _guard8428;
wire _guard8430 = _guard8424 | _guard8429;
wire _guard8431 = early_reset_static_par0_go_out;
wire _guard8432 = _guard8430 & _guard8431;
wire _guard8433 = fsm_out == 1'd0;
wire _guard8434 = cond_wire80_out;
wire _guard8435 = _guard8433 & _guard8434;
wire _guard8436 = fsm_out == 1'd0;
wire _guard8437 = _guard8435 & _guard8436;
wire _guard8438 = fsm_out == 1'd0;
wire _guard8439 = cond_wire82_out;
wire _guard8440 = _guard8438 & _guard8439;
wire _guard8441 = fsm_out == 1'd0;
wire _guard8442 = _guard8440 & _guard8441;
wire _guard8443 = _guard8437 | _guard8442;
wire _guard8444 = early_reset_static_par0_go_out;
wire _guard8445 = _guard8443 & _guard8444;
wire _guard8446 = cond_wire79_out;
wire _guard8447 = early_reset_static_par0_go_out;
wire _guard8448 = _guard8446 & _guard8447;
wire _guard8449 = cond_wire79_out;
wire _guard8450 = early_reset_static_par0_go_out;
wire _guard8451 = _guard8449 & _guard8450;
wire _guard8452 = cond_wire81_out;
wire _guard8453 = early_reset_static_par0_go_out;
wire _guard8454 = _guard8452 & _guard8453;
wire _guard8455 = cond_wire81_out;
wire _guard8456 = early_reset_static_par0_go_out;
wire _guard8457 = _guard8455 & _guard8456;
wire _guard8458 = cond_wire11_out;
wire _guard8459 = early_reset_static_par0_go_out;
wire _guard8460 = _guard8458 & _guard8459;
wire _guard8461 = cond_wire11_out;
wire _guard8462 = early_reset_static_par0_go_out;
wire _guard8463 = _guard8461 & _guard8462;
wire _guard8464 = cond_wire121_out;
wire _guard8465 = early_reset_static_par0_go_out;
wire _guard8466 = _guard8464 & _guard8465;
wire _guard8467 = cond_wire121_out;
wire _guard8468 = early_reset_static_par0_go_out;
wire _guard8469 = _guard8467 & _guard8468;
wire _guard8470 = cond_wire76_out;
wire _guard8471 = early_reset_static_par0_go_out;
wire _guard8472 = _guard8470 & _guard8471;
wire _guard8473 = cond_wire76_out;
wire _guard8474 = early_reset_static_par0_go_out;
wire _guard8475 = _guard8473 & _guard8474;
wire _guard8476 = cond_wire144_out;
wire _guard8477 = early_reset_static_par0_go_out;
wire _guard8478 = _guard8476 & _guard8477;
wire _guard8479 = cond_wire144_out;
wire _guard8480 = early_reset_static_par0_go_out;
wire _guard8481 = _guard8479 & _guard8480;
wire _guard8482 = cond_wire178_out;
wire _guard8483 = early_reset_static_par0_go_out;
wire _guard8484 = _guard8482 & _guard8483;
wire _guard8485 = cond_wire178_out;
wire _guard8486 = early_reset_static_par0_go_out;
wire _guard8487 = _guard8485 & _guard8486;
wire _guard8488 = cond_wire129_out;
wire _guard8489 = early_reset_static_par0_go_out;
wire _guard8490 = _guard8488 & _guard8489;
wire _guard8491 = cond_wire129_out;
wire _guard8492 = early_reset_static_par0_go_out;
wire _guard8493 = _guard8491 & _guard8492;
wire _guard8494 = cond_wire211_out;
wire _guard8495 = early_reset_static_par0_go_out;
wire _guard8496 = _guard8494 & _guard8495;
wire _guard8497 = cond_wire211_out;
wire _guard8498 = early_reset_static_par0_go_out;
wire _guard8499 = _guard8497 & _guard8498;
wire _guard8500 = cond_wire220_out;
wire _guard8501 = early_reset_static_par0_go_out;
wire _guard8502 = _guard8500 & _guard8501;
wire _guard8503 = cond_wire218_out;
wire _guard8504 = early_reset_static_par0_go_out;
wire _guard8505 = _guard8503 & _guard8504;
wire _guard8506 = fsm_out == 1'd0;
wire _guard8507 = cond_wire218_out;
wire _guard8508 = _guard8506 & _guard8507;
wire _guard8509 = fsm_out == 1'd0;
wire _guard8510 = _guard8508 & _guard8509;
wire _guard8511 = fsm_out == 1'd0;
wire _guard8512 = cond_wire220_out;
wire _guard8513 = _guard8511 & _guard8512;
wire _guard8514 = fsm_out == 1'd0;
wire _guard8515 = _guard8513 & _guard8514;
wire _guard8516 = _guard8510 | _guard8515;
wire _guard8517 = early_reset_static_par0_go_out;
wire _guard8518 = _guard8516 & _guard8517;
wire _guard8519 = fsm_out == 1'd0;
wire _guard8520 = cond_wire218_out;
wire _guard8521 = _guard8519 & _guard8520;
wire _guard8522 = fsm_out == 1'd0;
wire _guard8523 = _guard8521 & _guard8522;
wire _guard8524 = fsm_out == 1'd0;
wire _guard8525 = cond_wire220_out;
wire _guard8526 = _guard8524 & _guard8525;
wire _guard8527 = fsm_out == 1'd0;
wire _guard8528 = _guard8526 & _guard8527;
wire _guard8529 = _guard8523 | _guard8528;
wire _guard8530 = early_reset_static_par0_go_out;
wire _guard8531 = _guard8529 & _guard8530;
wire _guard8532 = fsm_out == 1'd0;
wire _guard8533 = cond_wire218_out;
wire _guard8534 = _guard8532 & _guard8533;
wire _guard8535 = fsm_out == 1'd0;
wire _guard8536 = _guard8534 & _guard8535;
wire _guard8537 = fsm_out == 1'd0;
wire _guard8538 = cond_wire220_out;
wire _guard8539 = _guard8537 & _guard8538;
wire _guard8540 = fsm_out == 1'd0;
wire _guard8541 = _guard8539 & _guard8540;
wire _guard8542 = _guard8536 | _guard8541;
wire _guard8543 = early_reset_static_par0_go_out;
wire _guard8544 = _guard8542 & _guard8543;
wire _guard8545 = cond_wire232_out;
wire _guard8546 = early_reset_static_par0_go_out;
wire _guard8547 = _guard8545 & _guard8546;
wire _guard8548 = cond_wire230_out;
wire _guard8549 = early_reset_static_par0_go_out;
wire _guard8550 = _guard8548 & _guard8549;
wire _guard8551 = fsm_out == 1'd0;
wire _guard8552 = cond_wire230_out;
wire _guard8553 = _guard8551 & _guard8552;
wire _guard8554 = fsm_out == 1'd0;
wire _guard8555 = _guard8553 & _guard8554;
wire _guard8556 = fsm_out == 1'd0;
wire _guard8557 = cond_wire232_out;
wire _guard8558 = _guard8556 & _guard8557;
wire _guard8559 = fsm_out == 1'd0;
wire _guard8560 = _guard8558 & _guard8559;
wire _guard8561 = _guard8555 | _guard8560;
wire _guard8562 = early_reset_static_par0_go_out;
wire _guard8563 = _guard8561 & _guard8562;
wire _guard8564 = fsm_out == 1'd0;
wire _guard8565 = cond_wire230_out;
wire _guard8566 = _guard8564 & _guard8565;
wire _guard8567 = fsm_out == 1'd0;
wire _guard8568 = _guard8566 & _guard8567;
wire _guard8569 = fsm_out == 1'd0;
wire _guard8570 = cond_wire232_out;
wire _guard8571 = _guard8569 & _guard8570;
wire _guard8572 = fsm_out == 1'd0;
wire _guard8573 = _guard8571 & _guard8572;
wire _guard8574 = _guard8568 | _guard8573;
wire _guard8575 = early_reset_static_par0_go_out;
wire _guard8576 = _guard8574 & _guard8575;
wire _guard8577 = fsm_out == 1'd0;
wire _guard8578 = cond_wire230_out;
wire _guard8579 = _guard8577 & _guard8578;
wire _guard8580 = fsm_out == 1'd0;
wire _guard8581 = _guard8579 & _guard8580;
wire _guard8582 = fsm_out == 1'd0;
wire _guard8583 = cond_wire232_out;
wire _guard8584 = _guard8582 & _guard8583;
wire _guard8585 = fsm_out == 1'd0;
wire _guard8586 = _guard8584 & _guard8585;
wire _guard8587 = _guard8581 | _guard8586;
wire _guard8588 = early_reset_static_par0_go_out;
wire _guard8589 = _guard8587 & _guard8588;
wire _guard8590 = cond_wire236_out;
wire _guard8591 = early_reset_static_par0_go_out;
wire _guard8592 = _guard8590 & _guard8591;
wire _guard8593 = cond_wire234_out;
wire _guard8594 = early_reset_static_par0_go_out;
wire _guard8595 = _guard8593 & _guard8594;
wire _guard8596 = fsm_out == 1'd0;
wire _guard8597 = cond_wire234_out;
wire _guard8598 = _guard8596 & _guard8597;
wire _guard8599 = fsm_out == 1'd0;
wire _guard8600 = _guard8598 & _guard8599;
wire _guard8601 = fsm_out == 1'd0;
wire _guard8602 = cond_wire236_out;
wire _guard8603 = _guard8601 & _guard8602;
wire _guard8604 = fsm_out == 1'd0;
wire _guard8605 = _guard8603 & _guard8604;
wire _guard8606 = _guard8600 | _guard8605;
wire _guard8607 = early_reset_static_par0_go_out;
wire _guard8608 = _guard8606 & _guard8607;
wire _guard8609 = fsm_out == 1'd0;
wire _guard8610 = cond_wire234_out;
wire _guard8611 = _guard8609 & _guard8610;
wire _guard8612 = fsm_out == 1'd0;
wire _guard8613 = _guard8611 & _guard8612;
wire _guard8614 = fsm_out == 1'd0;
wire _guard8615 = cond_wire236_out;
wire _guard8616 = _guard8614 & _guard8615;
wire _guard8617 = fsm_out == 1'd0;
wire _guard8618 = _guard8616 & _guard8617;
wire _guard8619 = _guard8613 | _guard8618;
wire _guard8620 = early_reset_static_par0_go_out;
wire _guard8621 = _guard8619 & _guard8620;
wire _guard8622 = fsm_out == 1'd0;
wire _guard8623 = cond_wire234_out;
wire _guard8624 = _guard8622 & _guard8623;
wire _guard8625 = fsm_out == 1'd0;
wire _guard8626 = _guard8624 & _guard8625;
wire _guard8627 = fsm_out == 1'd0;
wire _guard8628 = cond_wire236_out;
wire _guard8629 = _guard8627 & _guard8628;
wire _guard8630 = fsm_out == 1'd0;
wire _guard8631 = _guard8629 & _guard8630;
wire _guard8632 = _guard8626 | _guard8631;
wire _guard8633 = early_reset_static_par0_go_out;
wire _guard8634 = _guard8632 & _guard8633;
wire _guard8635 = cond_wire235_out;
wire _guard8636 = early_reset_static_par0_go_out;
wire _guard8637 = _guard8635 & _guard8636;
wire _guard8638 = cond_wire235_out;
wire _guard8639 = early_reset_static_par0_go_out;
wire _guard8640 = _guard8638 & _guard8639;
wire _guard8641 = cond_wire251_out;
wire _guard8642 = early_reset_static_par0_go_out;
wire _guard8643 = _guard8641 & _guard8642;
wire _guard8644 = cond_wire251_out;
wire _guard8645 = early_reset_static_par0_go_out;
wire _guard8646 = _guard8644 & _guard8645;
wire _guard8647 = cond_wire259_out;
wire _guard8648 = early_reset_static_par0_go_out;
wire _guard8649 = _guard8647 & _guard8648;
wire _guard8650 = cond_wire259_out;
wire _guard8651 = early_reset_static_par0_go_out;
wire _guard8652 = _guard8650 & _guard8651;
wire _guard8653 = cond_wire231_out;
wire _guard8654 = early_reset_static_par0_go_out;
wire _guard8655 = _guard8653 & _guard8654;
wire _guard8656 = cond_wire231_out;
wire _guard8657 = early_reset_static_par0_go_out;
wire _guard8658 = _guard8656 & _guard8657;
wire _guard8659 = cond_wire358_out;
wire _guard8660 = early_reset_static_par0_go_out;
wire _guard8661 = _guard8659 & _guard8660;
wire _guard8662 = cond_wire356_out;
wire _guard8663 = early_reset_static_par0_go_out;
wire _guard8664 = _guard8662 & _guard8663;
wire _guard8665 = fsm_out == 1'd0;
wire _guard8666 = cond_wire356_out;
wire _guard8667 = _guard8665 & _guard8666;
wire _guard8668 = fsm_out == 1'd0;
wire _guard8669 = _guard8667 & _guard8668;
wire _guard8670 = fsm_out == 1'd0;
wire _guard8671 = cond_wire358_out;
wire _guard8672 = _guard8670 & _guard8671;
wire _guard8673 = fsm_out == 1'd0;
wire _guard8674 = _guard8672 & _guard8673;
wire _guard8675 = _guard8669 | _guard8674;
wire _guard8676 = early_reset_static_par0_go_out;
wire _guard8677 = _guard8675 & _guard8676;
wire _guard8678 = fsm_out == 1'd0;
wire _guard8679 = cond_wire356_out;
wire _guard8680 = _guard8678 & _guard8679;
wire _guard8681 = fsm_out == 1'd0;
wire _guard8682 = _guard8680 & _guard8681;
wire _guard8683 = fsm_out == 1'd0;
wire _guard8684 = cond_wire358_out;
wire _guard8685 = _guard8683 & _guard8684;
wire _guard8686 = fsm_out == 1'd0;
wire _guard8687 = _guard8685 & _guard8686;
wire _guard8688 = _guard8682 | _guard8687;
wire _guard8689 = early_reset_static_par0_go_out;
wire _guard8690 = _guard8688 & _guard8689;
wire _guard8691 = fsm_out == 1'd0;
wire _guard8692 = cond_wire356_out;
wire _guard8693 = _guard8691 & _guard8692;
wire _guard8694 = fsm_out == 1'd0;
wire _guard8695 = _guard8693 & _guard8694;
wire _guard8696 = fsm_out == 1'd0;
wire _guard8697 = cond_wire358_out;
wire _guard8698 = _guard8696 & _guard8697;
wire _guard8699 = fsm_out == 1'd0;
wire _guard8700 = _guard8698 & _guard8699;
wire _guard8701 = _guard8695 | _guard8700;
wire _guard8702 = early_reset_static_par0_go_out;
wire _guard8703 = _guard8701 & _guard8702;
wire _guard8704 = cond_wire414_out;
wire _guard8705 = early_reset_static_par0_go_out;
wire _guard8706 = _guard8704 & _guard8705;
wire _guard8707 = cond_wire414_out;
wire _guard8708 = early_reset_static_par0_go_out;
wire _guard8709 = _guard8707 & _guard8708;
wire _guard8710 = cond_wire488_out;
wire _guard8711 = early_reset_static_par0_go_out;
wire _guard8712 = _guard8710 & _guard8711;
wire _guard8713 = cond_wire486_out;
wire _guard8714 = early_reset_static_par0_go_out;
wire _guard8715 = _guard8713 & _guard8714;
wire _guard8716 = fsm_out == 1'd0;
wire _guard8717 = cond_wire486_out;
wire _guard8718 = _guard8716 & _guard8717;
wire _guard8719 = fsm_out == 1'd0;
wire _guard8720 = _guard8718 & _guard8719;
wire _guard8721 = fsm_out == 1'd0;
wire _guard8722 = cond_wire488_out;
wire _guard8723 = _guard8721 & _guard8722;
wire _guard8724 = fsm_out == 1'd0;
wire _guard8725 = _guard8723 & _guard8724;
wire _guard8726 = _guard8720 | _guard8725;
wire _guard8727 = early_reset_static_par0_go_out;
wire _guard8728 = _guard8726 & _guard8727;
wire _guard8729 = fsm_out == 1'd0;
wire _guard8730 = cond_wire486_out;
wire _guard8731 = _guard8729 & _guard8730;
wire _guard8732 = fsm_out == 1'd0;
wire _guard8733 = _guard8731 & _guard8732;
wire _guard8734 = fsm_out == 1'd0;
wire _guard8735 = cond_wire488_out;
wire _guard8736 = _guard8734 & _guard8735;
wire _guard8737 = fsm_out == 1'd0;
wire _guard8738 = _guard8736 & _guard8737;
wire _guard8739 = _guard8733 | _guard8738;
wire _guard8740 = early_reset_static_par0_go_out;
wire _guard8741 = _guard8739 & _guard8740;
wire _guard8742 = fsm_out == 1'd0;
wire _guard8743 = cond_wire486_out;
wire _guard8744 = _guard8742 & _guard8743;
wire _guard8745 = fsm_out == 1'd0;
wire _guard8746 = _guard8744 & _guard8745;
wire _guard8747 = fsm_out == 1'd0;
wire _guard8748 = cond_wire488_out;
wire _guard8749 = _guard8747 & _guard8748;
wire _guard8750 = fsm_out == 1'd0;
wire _guard8751 = _guard8749 & _guard8750;
wire _guard8752 = _guard8746 | _guard8751;
wire _guard8753 = early_reset_static_par0_go_out;
wire _guard8754 = _guard8752 & _guard8753;
wire _guard8755 = cond_wire499_out;
wire _guard8756 = early_reset_static_par0_go_out;
wire _guard8757 = _guard8755 & _guard8756;
wire _guard8758 = cond_wire499_out;
wire _guard8759 = early_reset_static_par0_go_out;
wire _guard8760 = _guard8758 & _guard8759;
wire _guard8761 = cond_wire450_out;
wire _guard8762 = early_reset_static_par0_go_out;
wire _guard8763 = _guard8761 & _guard8762;
wire _guard8764 = cond_wire450_out;
wire _guard8765 = early_reset_static_par0_go_out;
wire _guard8766 = _guard8764 & _guard8765;
wire _guard8767 = cond_wire541_out;
wire _guard8768 = early_reset_static_par0_go_out;
wire _guard8769 = _guard8767 & _guard8768;
wire _guard8770 = cond_wire539_out;
wire _guard8771 = early_reset_static_par0_go_out;
wire _guard8772 = _guard8770 & _guard8771;
wire _guard8773 = fsm_out == 1'd0;
wire _guard8774 = cond_wire539_out;
wire _guard8775 = _guard8773 & _guard8774;
wire _guard8776 = fsm_out == 1'd0;
wire _guard8777 = _guard8775 & _guard8776;
wire _guard8778 = fsm_out == 1'd0;
wire _guard8779 = cond_wire541_out;
wire _guard8780 = _guard8778 & _guard8779;
wire _guard8781 = fsm_out == 1'd0;
wire _guard8782 = _guard8780 & _guard8781;
wire _guard8783 = _guard8777 | _guard8782;
wire _guard8784 = early_reset_static_par0_go_out;
wire _guard8785 = _guard8783 & _guard8784;
wire _guard8786 = fsm_out == 1'd0;
wire _guard8787 = cond_wire539_out;
wire _guard8788 = _guard8786 & _guard8787;
wire _guard8789 = fsm_out == 1'd0;
wire _guard8790 = _guard8788 & _guard8789;
wire _guard8791 = fsm_out == 1'd0;
wire _guard8792 = cond_wire541_out;
wire _guard8793 = _guard8791 & _guard8792;
wire _guard8794 = fsm_out == 1'd0;
wire _guard8795 = _guard8793 & _guard8794;
wire _guard8796 = _guard8790 | _guard8795;
wire _guard8797 = early_reset_static_par0_go_out;
wire _guard8798 = _guard8796 & _guard8797;
wire _guard8799 = fsm_out == 1'd0;
wire _guard8800 = cond_wire539_out;
wire _guard8801 = _guard8799 & _guard8800;
wire _guard8802 = fsm_out == 1'd0;
wire _guard8803 = _guard8801 & _guard8802;
wire _guard8804 = fsm_out == 1'd0;
wire _guard8805 = cond_wire541_out;
wire _guard8806 = _guard8804 & _guard8805;
wire _guard8807 = fsm_out == 1'd0;
wire _guard8808 = _guard8806 & _guard8807;
wire _guard8809 = _guard8803 | _guard8808;
wire _guard8810 = early_reset_static_par0_go_out;
wire _guard8811 = _guard8809 & _guard8810;
wire _guard8812 = cond_wire540_out;
wire _guard8813 = early_reset_static_par0_go_out;
wire _guard8814 = _guard8812 & _guard8813;
wire _guard8815 = cond_wire540_out;
wire _guard8816 = early_reset_static_par0_go_out;
wire _guard8817 = _guard8815 & _guard8816;
wire _guard8818 = cond_wire560_out;
wire _guard8819 = early_reset_static_par0_go_out;
wire _guard8820 = _guard8818 & _guard8819;
wire _guard8821 = cond_wire560_out;
wire _guard8822 = early_reset_static_par0_go_out;
wire _guard8823 = _guard8821 & _guard8822;
wire _guard8824 = cond_wire552_out;
wire _guard8825 = early_reset_static_par0_go_out;
wire _guard8826 = _guard8824 & _guard8825;
wire _guard8827 = cond_wire552_out;
wire _guard8828 = early_reset_static_par0_go_out;
wire _guard8829 = _guard8827 & _guard8828;
wire _guard8830 = cond_wire613_out;
wire _guard8831 = early_reset_static_par0_go_out;
wire _guard8832 = _guard8830 & _guard8831;
wire _guard8833 = cond_wire613_out;
wire _guard8834 = early_reset_static_par0_go_out;
wire _guard8835 = _guard8833 & _guard8834;
wire _guard8836 = cond_wire638_out;
wire _guard8837 = early_reset_static_par0_go_out;
wire _guard8838 = _guard8836 & _guard8837;
wire _guard8839 = cond_wire636_out;
wire _guard8840 = early_reset_static_par0_go_out;
wire _guard8841 = _guard8839 & _guard8840;
wire _guard8842 = fsm_out == 1'd0;
wire _guard8843 = cond_wire636_out;
wire _guard8844 = _guard8842 & _guard8843;
wire _guard8845 = fsm_out == 1'd0;
wire _guard8846 = _guard8844 & _guard8845;
wire _guard8847 = fsm_out == 1'd0;
wire _guard8848 = cond_wire638_out;
wire _guard8849 = _guard8847 & _guard8848;
wire _guard8850 = fsm_out == 1'd0;
wire _guard8851 = _guard8849 & _guard8850;
wire _guard8852 = _guard8846 | _guard8851;
wire _guard8853 = early_reset_static_par0_go_out;
wire _guard8854 = _guard8852 & _guard8853;
wire _guard8855 = fsm_out == 1'd0;
wire _guard8856 = cond_wire636_out;
wire _guard8857 = _guard8855 & _guard8856;
wire _guard8858 = fsm_out == 1'd0;
wire _guard8859 = _guard8857 & _guard8858;
wire _guard8860 = fsm_out == 1'd0;
wire _guard8861 = cond_wire638_out;
wire _guard8862 = _guard8860 & _guard8861;
wire _guard8863 = fsm_out == 1'd0;
wire _guard8864 = _guard8862 & _guard8863;
wire _guard8865 = _guard8859 | _guard8864;
wire _guard8866 = early_reset_static_par0_go_out;
wire _guard8867 = _guard8865 & _guard8866;
wire _guard8868 = fsm_out == 1'd0;
wire _guard8869 = cond_wire636_out;
wire _guard8870 = _guard8868 & _guard8869;
wire _guard8871 = fsm_out == 1'd0;
wire _guard8872 = _guard8870 & _guard8871;
wire _guard8873 = fsm_out == 1'd0;
wire _guard8874 = cond_wire638_out;
wire _guard8875 = _guard8873 & _guard8874;
wire _guard8876 = fsm_out == 1'd0;
wire _guard8877 = _guard8875 & _guard8876;
wire _guard8878 = _guard8872 | _guard8877;
wire _guard8879 = early_reset_static_par0_go_out;
wire _guard8880 = _guard8878 & _guard8879;
wire _guard8881 = cond_wire584_out;
wire _guard8882 = early_reset_static_par0_go_out;
wire _guard8883 = _guard8881 & _guard8882;
wire _guard8884 = cond_wire584_out;
wire _guard8885 = early_reset_static_par0_go_out;
wire _guard8886 = _guard8884 & _guard8885;
wire _guard8887 = cond_wire654_out;
wire _guard8888 = early_reset_static_par0_go_out;
wire _guard8889 = _guard8887 & _guard8888;
wire _guard8890 = cond_wire652_out;
wire _guard8891 = early_reset_static_par0_go_out;
wire _guard8892 = _guard8890 & _guard8891;
wire _guard8893 = fsm_out == 1'd0;
wire _guard8894 = cond_wire652_out;
wire _guard8895 = _guard8893 & _guard8894;
wire _guard8896 = fsm_out == 1'd0;
wire _guard8897 = _guard8895 & _guard8896;
wire _guard8898 = fsm_out == 1'd0;
wire _guard8899 = cond_wire654_out;
wire _guard8900 = _guard8898 & _guard8899;
wire _guard8901 = fsm_out == 1'd0;
wire _guard8902 = _guard8900 & _guard8901;
wire _guard8903 = _guard8897 | _guard8902;
wire _guard8904 = early_reset_static_par0_go_out;
wire _guard8905 = _guard8903 & _guard8904;
wire _guard8906 = fsm_out == 1'd0;
wire _guard8907 = cond_wire652_out;
wire _guard8908 = _guard8906 & _guard8907;
wire _guard8909 = fsm_out == 1'd0;
wire _guard8910 = _guard8908 & _guard8909;
wire _guard8911 = fsm_out == 1'd0;
wire _guard8912 = cond_wire654_out;
wire _guard8913 = _guard8911 & _guard8912;
wire _guard8914 = fsm_out == 1'd0;
wire _guard8915 = _guard8913 & _guard8914;
wire _guard8916 = _guard8910 | _guard8915;
wire _guard8917 = early_reset_static_par0_go_out;
wire _guard8918 = _guard8916 & _guard8917;
wire _guard8919 = fsm_out == 1'd0;
wire _guard8920 = cond_wire652_out;
wire _guard8921 = _guard8919 & _guard8920;
wire _guard8922 = fsm_out == 1'd0;
wire _guard8923 = _guard8921 & _guard8922;
wire _guard8924 = fsm_out == 1'd0;
wire _guard8925 = cond_wire654_out;
wire _guard8926 = _guard8924 & _guard8925;
wire _guard8927 = fsm_out == 1'd0;
wire _guard8928 = _guard8926 & _guard8927;
wire _guard8929 = _guard8923 | _guard8928;
wire _guard8930 = early_reset_static_par0_go_out;
wire _guard8931 = _guard8929 & _guard8930;
wire _guard8932 = cond_wire609_out;
wire _guard8933 = early_reset_static_par0_go_out;
wire _guard8934 = _guard8932 & _guard8933;
wire _guard8935 = cond_wire609_out;
wire _guard8936 = early_reset_static_par0_go_out;
wire _guard8937 = _guard8935 & _guard8936;
wire _guard8938 = cond_wire699_out;
wire _guard8939 = early_reset_static_par0_go_out;
wire _guard8940 = _guard8938 & _guard8939;
wire _guard8941 = cond_wire697_out;
wire _guard8942 = early_reset_static_par0_go_out;
wire _guard8943 = _guard8941 & _guard8942;
wire _guard8944 = fsm_out == 1'd0;
wire _guard8945 = cond_wire697_out;
wire _guard8946 = _guard8944 & _guard8945;
wire _guard8947 = fsm_out == 1'd0;
wire _guard8948 = _guard8946 & _guard8947;
wire _guard8949 = fsm_out == 1'd0;
wire _guard8950 = cond_wire699_out;
wire _guard8951 = _guard8949 & _guard8950;
wire _guard8952 = fsm_out == 1'd0;
wire _guard8953 = _guard8951 & _guard8952;
wire _guard8954 = _guard8948 | _guard8953;
wire _guard8955 = early_reset_static_par0_go_out;
wire _guard8956 = _guard8954 & _guard8955;
wire _guard8957 = fsm_out == 1'd0;
wire _guard8958 = cond_wire697_out;
wire _guard8959 = _guard8957 & _guard8958;
wire _guard8960 = fsm_out == 1'd0;
wire _guard8961 = _guard8959 & _guard8960;
wire _guard8962 = fsm_out == 1'd0;
wire _guard8963 = cond_wire699_out;
wire _guard8964 = _guard8962 & _guard8963;
wire _guard8965 = fsm_out == 1'd0;
wire _guard8966 = _guard8964 & _guard8965;
wire _guard8967 = _guard8961 | _guard8966;
wire _guard8968 = early_reset_static_par0_go_out;
wire _guard8969 = _guard8967 & _guard8968;
wire _guard8970 = fsm_out == 1'd0;
wire _guard8971 = cond_wire697_out;
wire _guard8972 = _guard8970 & _guard8971;
wire _guard8973 = fsm_out == 1'd0;
wire _guard8974 = _guard8972 & _guard8973;
wire _guard8975 = fsm_out == 1'd0;
wire _guard8976 = cond_wire699_out;
wire _guard8977 = _guard8975 & _guard8976;
wire _guard8978 = fsm_out == 1'd0;
wire _guard8979 = _guard8977 & _guard8978;
wire _guard8980 = _guard8974 | _guard8979;
wire _guard8981 = early_reset_static_par0_go_out;
wire _guard8982 = _guard8980 & _guard8981;
wire _guard8983 = cond_wire719_out;
wire _guard8984 = early_reset_static_par0_go_out;
wire _guard8985 = _guard8983 & _guard8984;
wire _guard8986 = cond_wire717_out;
wire _guard8987 = early_reset_static_par0_go_out;
wire _guard8988 = _guard8986 & _guard8987;
wire _guard8989 = fsm_out == 1'd0;
wire _guard8990 = cond_wire717_out;
wire _guard8991 = _guard8989 & _guard8990;
wire _guard8992 = fsm_out == 1'd0;
wire _guard8993 = _guard8991 & _guard8992;
wire _guard8994 = fsm_out == 1'd0;
wire _guard8995 = cond_wire719_out;
wire _guard8996 = _guard8994 & _guard8995;
wire _guard8997 = fsm_out == 1'd0;
wire _guard8998 = _guard8996 & _guard8997;
wire _guard8999 = _guard8993 | _guard8998;
wire _guard9000 = early_reset_static_par0_go_out;
wire _guard9001 = _guard8999 & _guard9000;
wire _guard9002 = fsm_out == 1'd0;
wire _guard9003 = cond_wire717_out;
wire _guard9004 = _guard9002 & _guard9003;
wire _guard9005 = fsm_out == 1'd0;
wire _guard9006 = _guard9004 & _guard9005;
wire _guard9007 = fsm_out == 1'd0;
wire _guard9008 = cond_wire719_out;
wire _guard9009 = _guard9007 & _guard9008;
wire _guard9010 = fsm_out == 1'd0;
wire _guard9011 = _guard9009 & _guard9010;
wire _guard9012 = _guard9006 | _guard9011;
wire _guard9013 = early_reset_static_par0_go_out;
wire _guard9014 = _guard9012 & _guard9013;
wire _guard9015 = fsm_out == 1'd0;
wire _guard9016 = cond_wire717_out;
wire _guard9017 = _guard9015 & _guard9016;
wire _guard9018 = fsm_out == 1'd0;
wire _guard9019 = _guard9017 & _guard9018;
wire _guard9020 = fsm_out == 1'd0;
wire _guard9021 = cond_wire719_out;
wire _guard9022 = _guard9020 & _guard9021;
wire _guard9023 = fsm_out == 1'd0;
wire _guard9024 = _guard9022 & _guard9023;
wire _guard9025 = _guard9019 | _guard9024;
wire _guard9026 = early_reset_static_par0_go_out;
wire _guard9027 = _guard9025 & _guard9026;
wire _guard9028 = cond_wire698_out;
wire _guard9029 = early_reset_static_par0_go_out;
wire _guard9030 = _guard9028 & _guard9029;
wire _guard9031 = cond_wire698_out;
wire _guard9032 = early_reset_static_par0_go_out;
wire _guard9033 = _guard9031 & _guard9032;
wire _guard9034 = cond_wire759_out;
wire _guard9035 = early_reset_static_par0_go_out;
wire _guard9036 = _guard9034 & _guard9035;
wire _guard9037 = cond_wire759_out;
wire _guard9038 = early_reset_static_par0_go_out;
wire _guard9039 = _guard9037 & _guard9038;
wire _guard9040 = cond_wire844_out;
wire _guard9041 = early_reset_static_par0_go_out;
wire _guard9042 = _guard9040 & _guard9041;
wire _guard9043 = cond_wire844_out;
wire _guard9044 = early_reset_static_par0_go_out;
wire _guard9045 = _guard9043 & _guard9044;
wire _guard9046 = cond_wire816_out;
wire _guard9047 = early_reset_static_par0_go_out;
wire _guard9048 = _guard9046 & _guard9047;
wire _guard9049 = cond_wire816_out;
wire _guard9050 = early_reset_static_par0_go_out;
wire _guard9051 = _guard9049 & _guard9050;
wire _guard9052 = cond_wire931_out;
wire _guard9053 = early_reset_static_par0_go_out;
wire _guard9054 = _guard9052 & _guard9053;
wire _guard9055 = cond_wire929_out;
wire _guard9056 = early_reset_static_par0_go_out;
wire _guard9057 = _guard9055 & _guard9056;
wire _guard9058 = fsm_out == 1'd0;
wire _guard9059 = cond_wire929_out;
wire _guard9060 = _guard9058 & _guard9059;
wire _guard9061 = fsm_out == 1'd0;
wire _guard9062 = _guard9060 & _guard9061;
wire _guard9063 = fsm_out == 1'd0;
wire _guard9064 = cond_wire931_out;
wire _guard9065 = _guard9063 & _guard9064;
wire _guard9066 = fsm_out == 1'd0;
wire _guard9067 = _guard9065 & _guard9066;
wire _guard9068 = _guard9062 | _guard9067;
wire _guard9069 = early_reset_static_par0_go_out;
wire _guard9070 = _guard9068 & _guard9069;
wire _guard9071 = fsm_out == 1'd0;
wire _guard9072 = cond_wire929_out;
wire _guard9073 = _guard9071 & _guard9072;
wire _guard9074 = fsm_out == 1'd0;
wire _guard9075 = _guard9073 & _guard9074;
wire _guard9076 = fsm_out == 1'd0;
wire _guard9077 = cond_wire931_out;
wire _guard9078 = _guard9076 & _guard9077;
wire _guard9079 = fsm_out == 1'd0;
wire _guard9080 = _guard9078 & _guard9079;
wire _guard9081 = _guard9075 | _guard9080;
wire _guard9082 = early_reset_static_par0_go_out;
wire _guard9083 = _guard9081 & _guard9082;
wire _guard9084 = fsm_out == 1'd0;
wire _guard9085 = cond_wire929_out;
wire _guard9086 = _guard9084 & _guard9085;
wire _guard9087 = fsm_out == 1'd0;
wire _guard9088 = _guard9086 & _guard9087;
wire _guard9089 = fsm_out == 1'd0;
wire _guard9090 = cond_wire931_out;
wire _guard9091 = _guard9089 & _guard9090;
wire _guard9092 = fsm_out == 1'd0;
wire _guard9093 = _guard9091 & _guard9092;
wire _guard9094 = _guard9088 | _guard9093;
wire _guard9095 = early_reset_static_par0_go_out;
wire _guard9096 = _guard9094 & _guard9095;
wire _guard9097 = cond_wire955_out;
wire _guard9098 = early_reset_static_par0_go_out;
wire _guard9099 = _guard9097 & _guard9098;
wire _guard9100 = cond_wire953_out;
wire _guard9101 = early_reset_static_par0_go_out;
wire _guard9102 = _guard9100 & _guard9101;
wire _guard9103 = fsm_out == 1'd0;
wire _guard9104 = cond_wire953_out;
wire _guard9105 = _guard9103 & _guard9104;
wire _guard9106 = fsm_out == 1'd0;
wire _guard9107 = _guard9105 & _guard9106;
wire _guard9108 = fsm_out == 1'd0;
wire _guard9109 = cond_wire955_out;
wire _guard9110 = _guard9108 & _guard9109;
wire _guard9111 = fsm_out == 1'd0;
wire _guard9112 = _guard9110 & _guard9111;
wire _guard9113 = _guard9107 | _guard9112;
wire _guard9114 = early_reset_static_par0_go_out;
wire _guard9115 = _guard9113 & _guard9114;
wire _guard9116 = fsm_out == 1'd0;
wire _guard9117 = cond_wire953_out;
wire _guard9118 = _guard9116 & _guard9117;
wire _guard9119 = fsm_out == 1'd0;
wire _guard9120 = _guard9118 & _guard9119;
wire _guard9121 = fsm_out == 1'd0;
wire _guard9122 = cond_wire955_out;
wire _guard9123 = _guard9121 & _guard9122;
wire _guard9124 = fsm_out == 1'd0;
wire _guard9125 = _guard9123 & _guard9124;
wire _guard9126 = _guard9120 | _guard9125;
wire _guard9127 = early_reset_static_par0_go_out;
wire _guard9128 = _guard9126 & _guard9127;
wire _guard9129 = fsm_out == 1'd0;
wire _guard9130 = cond_wire953_out;
wire _guard9131 = _guard9129 & _guard9130;
wire _guard9132 = fsm_out == 1'd0;
wire _guard9133 = _guard9131 & _guard9132;
wire _guard9134 = fsm_out == 1'd0;
wire _guard9135 = cond_wire955_out;
wire _guard9136 = _guard9134 & _guard9135;
wire _guard9137 = fsm_out == 1'd0;
wire _guard9138 = _guard9136 & _guard9137;
wire _guard9139 = _guard9133 | _guard9138;
wire _guard9140 = early_reset_static_par0_go_out;
wire _guard9141 = _guard9139 & _guard9140;
wire _guard9142 = cond_wire959_out;
wire _guard9143 = early_reset_static_par0_go_out;
wire _guard9144 = _guard9142 & _guard9143;
wire _guard9145 = cond_wire957_out;
wire _guard9146 = early_reset_static_par0_go_out;
wire _guard9147 = _guard9145 & _guard9146;
wire _guard9148 = fsm_out == 1'd0;
wire _guard9149 = cond_wire957_out;
wire _guard9150 = _guard9148 & _guard9149;
wire _guard9151 = fsm_out == 1'd0;
wire _guard9152 = _guard9150 & _guard9151;
wire _guard9153 = fsm_out == 1'd0;
wire _guard9154 = cond_wire959_out;
wire _guard9155 = _guard9153 & _guard9154;
wire _guard9156 = fsm_out == 1'd0;
wire _guard9157 = _guard9155 & _guard9156;
wire _guard9158 = _guard9152 | _guard9157;
wire _guard9159 = early_reset_static_par0_go_out;
wire _guard9160 = _guard9158 & _guard9159;
wire _guard9161 = fsm_out == 1'd0;
wire _guard9162 = cond_wire957_out;
wire _guard9163 = _guard9161 & _guard9162;
wire _guard9164 = fsm_out == 1'd0;
wire _guard9165 = _guard9163 & _guard9164;
wire _guard9166 = fsm_out == 1'd0;
wire _guard9167 = cond_wire959_out;
wire _guard9168 = _guard9166 & _guard9167;
wire _guard9169 = fsm_out == 1'd0;
wire _guard9170 = _guard9168 & _guard9169;
wire _guard9171 = _guard9165 | _guard9170;
wire _guard9172 = early_reset_static_par0_go_out;
wire _guard9173 = _guard9171 & _guard9172;
wire _guard9174 = fsm_out == 1'd0;
wire _guard9175 = cond_wire957_out;
wire _guard9176 = _guard9174 & _guard9175;
wire _guard9177 = fsm_out == 1'd0;
wire _guard9178 = _guard9176 & _guard9177;
wire _guard9179 = fsm_out == 1'd0;
wire _guard9180 = cond_wire959_out;
wire _guard9181 = _guard9179 & _guard9180;
wire _guard9182 = fsm_out == 1'd0;
wire _guard9183 = _guard9181 & _guard9182;
wire _guard9184 = _guard9178 | _guard9183;
wire _guard9185 = early_reset_static_par0_go_out;
wire _guard9186 = _guard9184 & _guard9185;
wire _guard9187 = cond_wire963_out;
wire _guard9188 = early_reset_static_par0_go_out;
wire _guard9189 = _guard9187 & _guard9188;
wire _guard9190 = cond_wire961_out;
wire _guard9191 = early_reset_static_par0_go_out;
wire _guard9192 = _guard9190 & _guard9191;
wire _guard9193 = fsm_out == 1'd0;
wire _guard9194 = cond_wire961_out;
wire _guard9195 = _guard9193 & _guard9194;
wire _guard9196 = fsm_out == 1'd0;
wire _guard9197 = _guard9195 & _guard9196;
wire _guard9198 = fsm_out == 1'd0;
wire _guard9199 = cond_wire963_out;
wire _guard9200 = _guard9198 & _guard9199;
wire _guard9201 = fsm_out == 1'd0;
wire _guard9202 = _guard9200 & _guard9201;
wire _guard9203 = _guard9197 | _guard9202;
wire _guard9204 = early_reset_static_par0_go_out;
wire _guard9205 = _guard9203 & _guard9204;
wire _guard9206 = fsm_out == 1'd0;
wire _guard9207 = cond_wire961_out;
wire _guard9208 = _guard9206 & _guard9207;
wire _guard9209 = fsm_out == 1'd0;
wire _guard9210 = _guard9208 & _guard9209;
wire _guard9211 = fsm_out == 1'd0;
wire _guard9212 = cond_wire963_out;
wire _guard9213 = _guard9211 & _guard9212;
wire _guard9214 = fsm_out == 1'd0;
wire _guard9215 = _guard9213 & _guard9214;
wire _guard9216 = _guard9210 | _guard9215;
wire _guard9217 = early_reset_static_par0_go_out;
wire _guard9218 = _guard9216 & _guard9217;
wire _guard9219 = fsm_out == 1'd0;
wire _guard9220 = cond_wire961_out;
wire _guard9221 = _guard9219 & _guard9220;
wire _guard9222 = fsm_out == 1'd0;
wire _guard9223 = _guard9221 & _guard9222;
wire _guard9224 = fsm_out == 1'd0;
wire _guard9225 = cond_wire963_out;
wire _guard9226 = _guard9224 & _guard9225;
wire _guard9227 = fsm_out == 1'd0;
wire _guard9228 = _guard9226 & _guard9227;
wire _guard9229 = _guard9223 | _guard9228;
wire _guard9230 = early_reset_static_par0_go_out;
wire _guard9231 = _guard9229 & _guard9230;
wire _guard9232 = cond_wire897_out;
wire _guard9233 = early_reset_static_par0_go_out;
wire _guard9234 = _guard9232 & _guard9233;
wire _guard9235 = cond_wire897_out;
wire _guard9236 = early_reset_static_par0_go_out;
wire _guard9237 = _guard9235 & _guard9236;
wire _guard9238 = cond_wire905_out;
wire _guard9239 = early_reset_static_par0_go_out;
wire _guard9240 = _guard9238 & _guard9239;
wire _guard9241 = cond_wire905_out;
wire _guard9242 = early_reset_static_par0_go_out;
wire _guard9243 = _guard9241 & _guard9242;
wire _guard9244 = cond_wire983_out;
wire _guard9245 = early_reset_static_par0_go_out;
wire _guard9246 = _guard9244 & _guard9245;
wire _guard9247 = cond_wire981_out;
wire _guard9248 = early_reset_static_par0_go_out;
wire _guard9249 = _guard9247 & _guard9248;
wire _guard9250 = fsm_out == 1'd0;
wire _guard9251 = cond_wire981_out;
wire _guard9252 = _guard9250 & _guard9251;
wire _guard9253 = fsm_out == 1'd0;
wire _guard9254 = _guard9252 & _guard9253;
wire _guard9255 = fsm_out == 1'd0;
wire _guard9256 = cond_wire983_out;
wire _guard9257 = _guard9255 & _guard9256;
wire _guard9258 = fsm_out == 1'd0;
wire _guard9259 = _guard9257 & _guard9258;
wire _guard9260 = _guard9254 | _guard9259;
wire _guard9261 = early_reset_static_par0_go_out;
wire _guard9262 = _guard9260 & _guard9261;
wire _guard9263 = fsm_out == 1'd0;
wire _guard9264 = cond_wire981_out;
wire _guard9265 = _guard9263 & _guard9264;
wire _guard9266 = fsm_out == 1'd0;
wire _guard9267 = _guard9265 & _guard9266;
wire _guard9268 = fsm_out == 1'd0;
wire _guard9269 = cond_wire983_out;
wire _guard9270 = _guard9268 & _guard9269;
wire _guard9271 = fsm_out == 1'd0;
wire _guard9272 = _guard9270 & _guard9271;
wire _guard9273 = _guard9267 | _guard9272;
wire _guard9274 = early_reset_static_par0_go_out;
wire _guard9275 = _guard9273 & _guard9274;
wire _guard9276 = fsm_out == 1'd0;
wire _guard9277 = cond_wire981_out;
wire _guard9278 = _guard9276 & _guard9277;
wire _guard9279 = fsm_out == 1'd0;
wire _guard9280 = _guard9278 & _guard9279;
wire _guard9281 = fsm_out == 1'd0;
wire _guard9282 = cond_wire983_out;
wire _guard9283 = _guard9281 & _guard9282;
wire _guard9284 = fsm_out == 1'd0;
wire _guard9285 = _guard9283 & _guard9284;
wire _guard9286 = _guard9280 | _guard9285;
wire _guard9287 = early_reset_static_par0_go_out;
wire _guard9288 = _guard9286 & _guard9287;
wire _guard9289 = cond_wire982_out;
wire _guard9290 = early_reset_static_par0_go_out;
wire _guard9291 = _guard9289 & _guard9290;
wire _guard9292 = cond_wire982_out;
wire _guard9293 = early_reset_static_par0_go_out;
wire _guard9294 = _guard9292 & _guard9293;
wire _guard9295 = cond_wire1028_out;
wire _guard9296 = early_reset_static_par0_go_out;
wire _guard9297 = _guard9295 & _guard9296;
wire _guard9298 = cond_wire1026_out;
wire _guard9299 = early_reset_static_par0_go_out;
wire _guard9300 = _guard9298 & _guard9299;
wire _guard9301 = fsm_out == 1'd0;
wire _guard9302 = cond_wire1026_out;
wire _guard9303 = _guard9301 & _guard9302;
wire _guard9304 = fsm_out == 1'd0;
wire _guard9305 = _guard9303 & _guard9304;
wire _guard9306 = fsm_out == 1'd0;
wire _guard9307 = cond_wire1028_out;
wire _guard9308 = _guard9306 & _guard9307;
wire _guard9309 = fsm_out == 1'd0;
wire _guard9310 = _guard9308 & _guard9309;
wire _guard9311 = _guard9305 | _guard9310;
wire _guard9312 = early_reset_static_par0_go_out;
wire _guard9313 = _guard9311 & _guard9312;
wire _guard9314 = fsm_out == 1'd0;
wire _guard9315 = cond_wire1026_out;
wire _guard9316 = _guard9314 & _guard9315;
wire _guard9317 = fsm_out == 1'd0;
wire _guard9318 = _guard9316 & _guard9317;
wire _guard9319 = fsm_out == 1'd0;
wire _guard9320 = cond_wire1028_out;
wire _guard9321 = _guard9319 & _guard9320;
wire _guard9322 = fsm_out == 1'd0;
wire _guard9323 = _guard9321 & _guard9322;
wire _guard9324 = _guard9318 | _guard9323;
wire _guard9325 = early_reset_static_par0_go_out;
wire _guard9326 = _guard9324 & _guard9325;
wire _guard9327 = fsm_out == 1'd0;
wire _guard9328 = cond_wire1026_out;
wire _guard9329 = _guard9327 & _guard9328;
wire _guard9330 = fsm_out == 1'd0;
wire _guard9331 = _guard9329 & _guard9330;
wire _guard9332 = fsm_out == 1'd0;
wire _guard9333 = cond_wire1028_out;
wire _guard9334 = _guard9332 & _guard9333;
wire _guard9335 = fsm_out == 1'd0;
wire _guard9336 = _guard9334 & _guard9335;
wire _guard9337 = _guard9331 | _guard9336;
wire _guard9338 = early_reset_static_par0_go_out;
wire _guard9339 = _guard9337 & _guard9338;
wire _guard9340 = cond_wire962_out;
wire _guard9341 = early_reset_static_par0_go_out;
wire _guard9342 = _guard9340 & _guard9341;
wire _guard9343 = cond_wire962_out;
wire _guard9344 = early_reset_static_par0_go_out;
wire _guard9345 = _guard9343 & _guard9344;
wire _guard9346 = cond_wire970_out;
wire _guard9347 = early_reset_static_par0_go_out;
wire _guard9348 = _guard9346 & _guard9347;
wire _guard9349 = cond_wire970_out;
wire _guard9350 = early_reset_static_par0_go_out;
wire _guard9351 = _guard9349 & _guard9350;
wire _guard9352 = cond_wire1043_out;
wire _guard9353 = early_reset_static_par0_go_out;
wire _guard9354 = _guard9352 & _guard9353;
wire _guard9355 = cond_wire1043_out;
wire _guard9356 = early_reset_static_par0_go_out;
wire _guard9357 = _guard9355 & _guard9356;
wire _guard9358 = fsm0_out == 6'd0;
wire _guard9359 = early_reset_static_seq_go_out;
wire _guard9360 = _guard9358 & _guard9359;
wire _guard9361 = cond_wire4_out;
wire _guard9362 = early_reset_static_par0_go_out;
wire _guard9363 = _guard9361 & _guard9362;
wire _guard9364 = _guard9360 | _guard9363;
wire _guard9365 = fsm0_out == 6'd0;
wire _guard9366 = early_reset_static_seq_go_out;
wire _guard9367 = _guard9365 & _guard9366;
wire _guard9368 = cond_wire4_out;
wire _guard9369 = early_reset_static_par0_go_out;
wire _guard9370 = _guard9368 & _guard9369;
wire _guard9371 = fsm0_out == 6'd0;
wire _guard9372 = early_reset_static_seq_go_out;
wire _guard9373 = _guard9371 & _guard9372;
wire _guard9374 = cond_wire34_out;
wire _guard9375 = early_reset_static_par0_go_out;
wire _guard9376 = _guard9374 & _guard9375;
wire _guard9377 = _guard9373 | _guard9376;
wire _guard9378 = fsm0_out == 6'd0;
wire _guard9379 = early_reset_static_seq_go_out;
wire _guard9380 = _guard9378 & _guard9379;
wire _guard9381 = cond_wire34_out;
wire _guard9382 = early_reset_static_par0_go_out;
wire _guard9383 = _guard9381 & _guard9382;
wire _guard9384 = fsm0_out == 6'd0;
wire _guard9385 = early_reset_static_seq_go_out;
wire _guard9386 = _guard9384 & _guard9385;
wire _guard9387 = cond_wire44_out;
wire _guard9388 = early_reset_static_par0_go_out;
wire _guard9389 = _guard9387 & _guard9388;
wire _guard9390 = _guard9386 | _guard9389;
wire _guard9391 = fsm0_out == 6'd0;
wire _guard9392 = early_reset_static_seq_go_out;
wire _guard9393 = _guard9391 & _guard9392;
wire _guard9394 = cond_wire44_out;
wire _guard9395 = early_reset_static_par0_go_out;
wire _guard9396 = _guard9394 & _guard9395;
wire _guard9397 = fsm0_out == 6'd0;
wire _guard9398 = early_reset_static_seq_go_out;
wire _guard9399 = _guard9397 & _guard9398;
wire _guard9400 = cond_wire599_out;
wire _guard9401 = early_reset_static_par0_go_out;
wire _guard9402 = _guard9400 & _guard9401;
wire _guard9403 = _guard9399 | _guard9402;
wire _guard9404 = fsm0_out == 6'd0;
wire _guard9405 = early_reset_static_seq_go_out;
wire _guard9406 = _guard9404 & _guard9405;
wire _guard9407 = cond_wire599_out;
wire _guard9408 = early_reset_static_par0_go_out;
wire _guard9409 = _guard9407 & _guard9408;
wire _guard9410 = cond_wire859_out;
wire _guard9411 = early_reset_static_par0_go_out;
wire _guard9412 = _guard9410 & _guard9411;
wire _guard9413 = cond_wire859_out;
wire _guard9414 = early_reset_static_par0_go_out;
wire _guard9415 = _guard9413 & _guard9414;
wire _guard9416 = early_reset_static_par0_go_out;
wire _guard9417 = early_reset_static_par0_go_out;
wire _guard9418 = early_reset_static_par0_go_out;
wire _guard9419 = early_reset_static_par0_go_out;
wire _guard9420 = early_reset_static_par0_go_out;
wire _guard9421 = early_reset_static_par0_go_out;
wire _guard9422 = fsm0_out == 6'd0;
wire _guard9423 = early_reset_static_seq_go_out;
wire _guard9424 = _guard9422 & _guard9423;
wire _guard9425 = early_reset_static_par0_go_out;
wire _guard9426 = _guard9424 | _guard9425;
wire _guard9427 = fsm0_out == 6'd0;
wire _guard9428 = early_reset_static_seq_go_out;
wire _guard9429 = _guard9427 & _guard9428;
wire _guard9430 = early_reset_static_par0_go_out;
wire _guard9431 = early_reset_static_par0_go_out;
wire _guard9432 = early_reset_static_par0_go_out;
wire _guard9433 = fsm0_out == 6'd0;
wire _guard9434 = early_reset_static_seq_go_out;
wire _guard9435 = _guard9433 & _guard9434;
wire _guard9436 = early_reset_static_par0_go_out;
wire _guard9437 = _guard9435 | _guard9436;
wire _guard9438 = fsm0_out == 6'd0;
wire _guard9439 = early_reset_static_seq_go_out;
wire _guard9440 = _guard9438 & _guard9439;
wire _guard9441 = early_reset_static_par0_go_out;
wire _guard9442 = early_reset_static_par0_go_out;
wire _guard9443 = early_reset_static_par0_go_out;
wire _guard9444 = early_reset_static_par0_go_out;
wire _guard9445 = early_reset_static_par0_go_out;
wire _guard9446 = early_reset_static_par0_go_out;
wire _guard9447 = early_reset_static_par0_go_out;
wire _guard9448 = fsm0_out == 6'd0;
wire _guard9449 = early_reset_static_seq_go_out;
wire _guard9450 = _guard9448 & _guard9449;
wire _guard9451 = early_reset_static_par0_go_out;
wire _guard9452 = _guard9450 | _guard9451;
wire _guard9453 = early_reset_static_par0_go_out;
wire _guard9454 = fsm0_out == 6'd0;
wire _guard9455 = early_reset_static_seq_go_out;
wire _guard9456 = _guard9454 & _guard9455;
wire _guard9457 = early_reset_static_par0_go_out;
wire _guard9458 = early_reset_static_par0_go_out;
wire _guard9459 = early_reset_static_par0_go_out;
wire _guard9460 = ~_guard0;
wire _guard9461 = early_reset_static_par0_go_out;
wire _guard9462 = _guard9460 & _guard9461;
wire _guard9463 = early_reset_static_par0_go_out;
wire _guard9464 = ~_guard0;
wire _guard9465 = early_reset_static_par0_go_out;
wire _guard9466 = _guard9464 & _guard9465;
wire _guard9467 = ~_guard0;
wire _guard9468 = early_reset_static_par0_go_out;
wire _guard9469 = _guard9467 & _guard9468;
wire _guard9470 = early_reset_static_par0_go_out;
wire _guard9471 = ~_guard0;
wire _guard9472 = early_reset_static_par0_go_out;
wire _guard9473 = _guard9471 & _guard9472;
wire _guard9474 = early_reset_static_par0_go_out;
wire _guard9475 = ~_guard0;
wire _guard9476 = early_reset_static_par0_go_out;
wire _guard9477 = _guard9475 & _guard9476;
wire _guard9478 = early_reset_static_par0_go_out;
wire _guard9479 = early_reset_static_par0_go_out;
wire _guard9480 = ~_guard0;
wire _guard9481 = early_reset_static_par0_go_out;
wire _guard9482 = _guard9480 & _guard9481;
wire _guard9483 = ~_guard0;
wire _guard9484 = early_reset_static_par0_go_out;
wire _guard9485 = _guard9483 & _guard9484;
wire _guard9486 = early_reset_static_par0_go_out;
wire _guard9487 = early_reset_static_par0_go_out;
wire _guard9488 = early_reset_static_par0_go_out;
wire _guard9489 = ~_guard0;
wire _guard9490 = early_reset_static_par0_go_out;
wire _guard9491 = _guard9489 & _guard9490;
wire _guard9492 = early_reset_static_par0_go_out;
wire _guard9493 = early_reset_static_par0_go_out;
wire _guard9494 = early_reset_static_par0_go_out;
wire _guard9495 = early_reset_static_par0_go_out;
wire _guard9496 = ~_guard0;
wire _guard9497 = early_reset_static_par0_go_out;
wire _guard9498 = _guard9496 & _guard9497;
wire _guard9499 = early_reset_static_par0_go_out;
wire _guard9500 = early_reset_static_par0_go_out;
wire _guard9501 = early_reset_static_par0_go_out;
wire _guard9502 = ~_guard0;
wire _guard9503 = early_reset_static_par0_go_out;
wire _guard9504 = _guard9502 & _guard9503;
wire _guard9505 = ~_guard0;
wire _guard9506 = early_reset_static_par0_go_out;
wire _guard9507 = _guard9505 & _guard9506;
wire _guard9508 = early_reset_static_par0_go_out;
wire _guard9509 = ~_guard0;
wire _guard9510 = early_reset_static_par0_go_out;
wire _guard9511 = _guard9509 & _guard9510;
wire _guard9512 = early_reset_static_par0_go_out;
wire _guard9513 = early_reset_static_par0_go_out;
wire _guard9514 = early_reset_static_par0_go_out;
wire _guard9515 = early_reset_static_par0_go_out;
wire _guard9516 = early_reset_static_par0_go_out;
wire _guard9517 = early_reset_static_par0_go_out;
wire _guard9518 = ~_guard0;
wire _guard9519 = early_reset_static_par0_go_out;
wire _guard9520 = _guard9518 & _guard9519;
wire _guard9521 = early_reset_static_par0_go_out;
wire _guard9522 = ~_guard0;
wire _guard9523 = early_reset_static_par0_go_out;
wire _guard9524 = _guard9522 & _guard9523;
wire _guard9525 = early_reset_static_par0_go_out;
wire _guard9526 = early_reset_static_par0_go_out;
wire _guard9527 = early_reset_static_par0_go_out;
wire _guard9528 = early_reset_static_par0_go_out;
wire _guard9529 = ~_guard0;
wire _guard9530 = early_reset_static_par0_go_out;
wire _guard9531 = _guard9529 & _guard9530;
wire _guard9532 = early_reset_static_par0_go_out;
wire _guard9533 = ~_guard0;
wire _guard9534 = early_reset_static_par0_go_out;
wire _guard9535 = _guard9533 & _guard9534;
wire _guard9536 = early_reset_static_par0_go_out;
wire _guard9537 = early_reset_static_par0_go_out;
wire _guard9538 = early_reset_static_par0_go_out;
wire _guard9539 = ~_guard0;
wire _guard9540 = early_reset_static_par0_go_out;
wire _guard9541 = _guard9539 & _guard9540;
wire _guard9542 = early_reset_static_par0_go_out;
wire _guard9543 = early_reset_static_par0_go_out;
wire _guard9544 = early_reset_static_par0_go_out;
wire _guard9545 = early_reset_static_par0_go_out;
wire _guard9546 = early_reset_static_par0_go_out;
wire _guard9547 = early_reset_static_par0_go_out;
wire _guard9548 = early_reset_static_par0_go_out;
wire _guard9549 = early_reset_static_par0_go_out;
wire _guard9550 = early_reset_static_par0_go_out;
wire _guard9551 = early_reset_static_par0_go_out;
wire _guard9552 = ~_guard0;
wire _guard9553 = early_reset_static_par0_go_out;
wire _guard9554 = _guard9552 & _guard9553;
wire _guard9555 = early_reset_static_par0_go_out;
wire _guard9556 = early_reset_static_par0_go_out;
wire _guard9557 = early_reset_static_par0_go_out;
wire _guard9558 = early_reset_static_par0_go_out;
wire _guard9559 = early_reset_static_par0_go_out;
wire _guard9560 = early_reset_static_par0_go_out;
wire _guard9561 = early_reset_static_par0_go_out;
wire _guard9562 = early_reset_static_par0_go_out;
wire _guard9563 = ~_guard0;
wire _guard9564 = early_reset_static_par0_go_out;
wire _guard9565 = _guard9563 & _guard9564;
wire _guard9566 = early_reset_static_par0_go_out;
wire _guard9567 = early_reset_static_par0_go_out;
wire _guard9568 = ~_guard0;
wire _guard9569 = early_reset_static_par0_go_out;
wire _guard9570 = _guard9568 & _guard9569;
wire _guard9571 = early_reset_static_par0_go_out;
wire _guard9572 = early_reset_static_par0_go_out;
wire _guard9573 = early_reset_static_par0_go_out;
wire _guard9574 = ~_guard0;
wire _guard9575 = early_reset_static_par0_go_out;
wire _guard9576 = _guard9574 & _guard9575;
wire _guard9577 = early_reset_static_par0_go_out;
wire _guard9578 = early_reset_static_par0_go_out;
wire _guard9579 = early_reset_static_par0_go_out;
wire _guard9580 = early_reset_static_par0_go_out;
wire _guard9581 = early_reset_static_par0_go_out;
wire _guard9582 = ~_guard0;
wire _guard9583 = early_reset_static_par0_go_out;
wire _guard9584 = _guard9582 & _guard9583;
wire _guard9585 = early_reset_static_par0_go_out;
wire _guard9586 = early_reset_static_par0_go_out;
wire _guard9587 = ~_guard0;
wire _guard9588 = early_reset_static_par0_go_out;
wire _guard9589 = _guard9587 & _guard9588;
wire _guard9590 = early_reset_static_par0_go_out;
wire _guard9591 = ~_guard0;
wire _guard9592 = early_reset_static_par0_go_out;
wire _guard9593 = _guard9591 & _guard9592;
wire _guard9594 = early_reset_static_par0_go_out;
wire _guard9595 = ~_guard0;
wire _guard9596 = early_reset_static_par0_go_out;
wire _guard9597 = _guard9595 & _guard9596;
wire _guard9598 = early_reset_static_par0_go_out;
wire _guard9599 = ~_guard0;
wire _guard9600 = early_reset_static_par0_go_out;
wire _guard9601 = _guard9599 & _guard9600;
wire _guard9602 = early_reset_static_par0_go_out;
wire _guard9603 = early_reset_static_par0_go_out;
wire _guard9604 = early_reset_static_par0_go_out;
wire _guard9605 = early_reset_static_par0_go_out;
wire _guard9606 = ~_guard0;
wire _guard9607 = early_reset_static_par0_go_out;
wire _guard9608 = _guard9606 & _guard9607;
wire _guard9609 = early_reset_static_par0_go_out;
wire _guard9610 = ~_guard0;
wire _guard9611 = early_reset_static_par0_go_out;
wire _guard9612 = _guard9610 & _guard9611;
wire _guard9613 = early_reset_static_par0_go_out;
wire _guard9614 = early_reset_static_par0_go_out;
wire _guard9615 = ~_guard0;
wire _guard9616 = early_reset_static_par0_go_out;
wire _guard9617 = _guard9615 & _guard9616;
wire _guard9618 = early_reset_static_par0_go_out;
wire _guard9619 = early_reset_static_par0_go_out;
wire _guard9620 = ~_guard0;
wire _guard9621 = early_reset_static_par0_go_out;
wire _guard9622 = _guard9620 & _guard9621;
wire _guard9623 = early_reset_static_par0_go_out;
wire _guard9624 = ~_guard0;
wire _guard9625 = early_reset_static_par0_go_out;
wire _guard9626 = _guard9624 & _guard9625;
wire _guard9627 = early_reset_static_par0_go_out;
wire _guard9628 = ~_guard0;
wire _guard9629 = early_reset_static_par0_go_out;
wire _guard9630 = _guard9628 & _guard9629;
wire _guard9631 = early_reset_static_par0_go_out;
wire _guard9632 = ~_guard0;
wire _guard9633 = early_reset_static_par0_go_out;
wire _guard9634 = _guard9632 & _guard9633;
wire _guard9635 = ~_guard0;
wire _guard9636 = early_reset_static_par0_go_out;
wire _guard9637 = _guard9635 & _guard9636;
wire _guard9638 = early_reset_static_par0_go_out;
wire _guard9639 = early_reset_static_par0_go_out;
wire _guard9640 = early_reset_static_par0_go_out;
wire _guard9641 = early_reset_static_par0_go_out;
wire _guard9642 = early_reset_static_par0_go_out;
wire _guard9643 = early_reset_static_par0_go_out;
wire _guard9644 = ~_guard0;
wire _guard9645 = early_reset_static_par0_go_out;
wire _guard9646 = _guard9644 & _guard9645;
wire _guard9647 = early_reset_static_par0_go_out;
wire _guard9648 = ~_guard0;
wire _guard9649 = early_reset_static_par0_go_out;
wire _guard9650 = _guard9648 & _guard9649;
wire _guard9651 = ~_guard0;
wire _guard9652 = early_reset_static_par0_go_out;
wire _guard9653 = _guard9651 & _guard9652;
wire _guard9654 = early_reset_static_par0_go_out;
wire _guard9655 = early_reset_static_par0_go_out;
wire _guard9656 = early_reset_static_par0_go_out;
wire _guard9657 = early_reset_static_par0_go_out;
wire _guard9658 = early_reset_static_par0_go_out;
wire _guard9659 = early_reset_static_par0_go_out;
wire _guard9660 = ~_guard0;
wire _guard9661 = early_reset_static_par0_go_out;
wire _guard9662 = _guard9660 & _guard9661;
wire _guard9663 = early_reset_static_par0_go_out;
wire _guard9664 = early_reset_static_par0_go_out;
wire _guard9665 = ~_guard0;
wire _guard9666 = early_reset_static_par0_go_out;
wire _guard9667 = _guard9665 & _guard9666;
wire _guard9668 = early_reset_static_par0_go_out;
wire _guard9669 = ~_guard0;
wire _guard9670 = early_reset_static_par0_go_out;
wire _guard9671 = _guard9669 & _guard9670;
wire _guard9672 = early_reset_static_par0_go_out;
wire _guard9673 = early_reset_static_par0_go_out;
wire _guard9674 = ~_guard0;
wire _guard9675 = early_reset_static_par0_go_out;
wire _guard9676 = _guard9674 & _guard9675;
wire _guard9677 = early_reset_static_par0_go_out;
wire _guard9678 = ~_guard0;
wire _guard9679 = early_reset_static_par0_go_out;
wire _guard9680 = _guard9678 & _guard9679;
wire _guard9681 = early_reset_static_par0_go_out;
wire _guard9682 = ~_guard0;
wire _guard9683 = early_reset_static_par0_go_out;
wire _guard9684 = _guard9682 & _guard9683;
wire _guard9685 = early_reset_static_par0_go_out;
wire _guard9686 = early_reset_static_par0_go_out;
wire _guard9687 = early_reset_static_par0_go_out;
wire _guard9688 = ~_guard0;
wire _guard9689 = early_reset_static_par0_go_out;
wire _guard9690 = _guard9688 & _guard9689;
wire _guard9691 = early_reset_static_par0_go_out;
wire _guard9692 = ~_guard0;
wire _guard9693 = early_reset_static_par0_go_out;
wire _guard9694 = _guard9692 & _guard9693;
wire _guard9695 = early_reset_static_par0_go_out;
wire _guard9696 = early_reset_static_par0_go_out;
wire _guard9697 = early_reset_static_par0_go_out;
wire _guard9698 = ~_guard0;
wire _guard9699 = early_reset_static_par0_go_out;
wire _guard9700 = _guard9698 & _guard9699;
wire _guard9701 = ~_guard0;
wire _guard9702 = early_reset_static_par0_go_out;
wire _guard9703 = _guard9701 & _guard9702;
wire _guard9704 = early_reset_static_par0_go_out;
wire _guard9705 = early_reset_static_par0_go_out;
wire _guard9706 = early_reset_static_par0_go_out;
wire _guard9707 = early_reset_static_par0_go_out;
wire _guard9708 = ~_guard0;
wire _guard9709 = early_reset_static_par0_go_out;
wire _guard9710 = _guard9708 & _guard9709;
wire _guard9711 = early_reset_static_par0_go_out;
wire _guard9712 = early_reset_static_par0_go_out;
wire _guard9713 = early_reset_static_par0_go_out;
wire _guard9714 = early_reset_static_par0_go_out;
wire _guard9715 = ~_guard0;
wire _guard9716 = early_reset_static_par0_go_out;
wire _guard9717 = _guard9715 & _guard9716;
wire _guard9718 = early_reset_static_par0_go_out;
wire _guard9719 = early_reset_static_par0_go_out;
wire _guard9720 = ~_guard0;
wire _guard9721 = early_reset_static_par0_go_out;
wire _guard9722 = _guard9720 & _guard9721;
wire _guard9723 = early_reset_static_par0_go_out;
wire _guard9724 = ~_guard0;
wire _guard9725 = early_reset_static_par0_go_out;
wire _guard9726 = _guard9724 & _guard9725;
wire _guard9727 = ~_guard0;
wire _guard9728 = early_reset_static_par0_go_out;
wire _guard9729 = _guard9727 & _guard9728;
wire _guard9730 = early_reset_static_par0_go_out;
wire _guard9731 = early_reset_static_par0_go_out;
wire _guard9732 = early_reset_static_par0_go_out;
wire _guard9733 = early_reset_static_par0_go_out;
wire _guard9734 = early_reset_static_par0_go_out;
wire _guard9735 = ~_guard0;
wire _guard9736 = early_reset_static_par0_go_out;
wire _guard9737 = _guard9735 & _guard9736;
wire _guard9738 = early_reset_static_par0_go_out;
wire _guard9739 = early_reset_static_par0_go_out;
wire _guard9740 = early_reset_static_par0_go_out;
wire _guard9741 = ~_guard0;
wire _guard9742 = early_reset_static_par0_go_out;
wire _guard9743 = _guard9741 & _guard9742;
wire _guard9744 = early_reset_static_par0_go_out;
wire _guard9745 = early_reset_static_par0_go_out;
wire _guard9746 = early_reset_static_par0_go_out;
wire _guard9747 = early_reset_static_par0_go_out;
wire _guard9748 = early_reset_static_par0_go_out;
wire _guard9749 = ~_guard0;
wire _guard9750 = early_reset_static_par0_go_out;
wire _guard9751 = _guard9749 & _guard9750;
wire _guard9752 = early_reset_static_par0_go_out;
wire _guard9753 = ~_guard0;
wire _guard9754 = early_reset_static_par0_go_out;
wire _guard9755 = _guard9753 & _guard9754;
wire _guard9756 = early_reset_static_par0_go_out;
wire _guard9757 = early_reset_static_par0_go_out;
wire _guard9758 = early_reset_static_par0_go_out;
wire _guard9759 = early_reset_static_par0_go_out;
wire _guard9760 = ~_guard0;
wire _guard9761 = early_reset_static_par0_go_out;
wire _guard9762 = _guard9760 & _guard9761;
wire _guard9763 = early_reset_static_par0_go_out;
wire _guard9764 = ~_guard0;
wire _guard9765 = early_reset_static_par0_go_out;
wire _guard9766 = _guard9764 & _guard9765;
wire _guard9767 = ~_guard0;
wire _guard9768 = early_reset_static_par0_go_out;
wire _guard9769 = _guard9767 & _guard9768;
wire _guard9770 = early_reset_static_par0_go_out;
wire _guard9771 = early_reset_static_par0_go_out;
wire _guard9772 = ~_guard0;
wire _guard9773 = early_reset_static_par0_go_out;
wire _guard9774 = _guard9772 & _guard9773;
wire _guard9775 = early_reset_static_par0_go_out;
wire _guard9776 = early_reset_static_par0_go_out;
wire _guard9777 = early_reset_static_par0_go_out;
wire _guard9778 = early_reset_static_par0_go_out;
wire _guard9779 = ~_guard0;
wire _guard9780 = early_reset_static_par0_go_out;
wire _guard9781 = _guard9779 & _guard9780;
wire _guard9782 = early_reset_static_par0_go_out;
wire _guard9783 = ~_guard0;
wire _guard9784 = early_reset_static_par0_go_out;
wire _guard9785 = _guard9783 & _guard9784;
wire _guard9786 = early_reset_static_par0_go_out;
wire _guard9787 = ~_guard0;
wire _guard9788 = early_reset_static_par0_go_out;
wire _guard9789 = _guard9787 & _guard9788;
wire _guard9790 = early_reset_static_par0_go_out;
wire _guard9791 = early_reset_static_par0_go_out;
wire _guard9792 = early_reset_static_par0_go_out;
wire _guard9793 = early_reset_static_par0_go_out;
wire _guard9794 = ~_guard0;
wire _guard9795 = early_reset_static_par0_go_out;
wire _guard9796 = _guard9794 & _guard9795;
wire _guard9797 = early_reset_static_par0_go_out;
wire _guard9798 = ~_guard0;
wire _guard9799 = early_reset_static_par0_go_out;
wire _guard9800 = _guard9798 & _guard9799;
wire _guard9801 = early_reset_static_par0_go_out;
wire _guard9802 = ~_guard0;
wire _guard9803 = early_reset_static_par0_go_out;
wire _guard9804 = _guard9802 & _guard9803;
wire _guard9805 = ~_guard0;
wire _guard9806 = early_reset_static_par0_go_out;
wire _guard9807 = _guard9805 & _guard9806;
wire _guard9808 = early_reset_static_par0_go_out;
wire _guard9809 = ~_guard0;
wire _guard9810 = early_reset_static_par0_go_out;
wire _guard9811 = _guard9809 & _guard9810;
wire _guard9812 = early_reset_static_par0_go_out;
wire _guard9813 = early_reset_static_par0_go_out;
wire _guard9814 = ~_guard0;
wire _guard9815 = early_reset_static_par0_go_out;
wire _guard9816 = _guard9814 & _guard9815;
wire _guard9817 = early_reset_static_par0_go_out;
wire _guard9818 = ~_guard0;
wire _guard9819 = early_reset_static_par0_go_out;
wire _guard9820 = _guard9818 & _guard9819;
wire _guard9821 = early_reset_static_par0_go_out;
wire _guard9822 = early_reset_static_par0_go_out;
wire _guard9823 = early_reset_static_par0_go_out;
wire _guard9824 = early_reset_static_par0_go_out;
wire _guard9825 = early_reset_static_par0_go_out;
wire _guard9826 = early_reset_static_par0_go_out;
wire _guard9827 = ~_guard0;
wire _guard9828 = early_reset_static_par0_go_out;
wire _guard9829 = _guard9827 & _guard9828;
wire _guard9830 = early_reset_static_par0_go_out;
wire _guard9831 = early_reset_static_par0_go_out;
wire _guard9832 = early_reset_static_par0_go_out;
wire _guard9833 = early_reset_static_par0_go_out;
wire _guard9834 = early_reset_static_par0_go_out;
wire _guard9835 = early_reset_static_par0_go_out;
wire _guard9836 = early_reset_static_par0_go_out;
wire _guard9837 = early_reset_static_par0_go_out;
wire _guard9838 = early_reset_static_par0_go_out;
wire _guard9839 = ~_guard0;
wire _guard9840 = early_reset_static_par0_go_out;
wire _guard9841 = _guard9839 & _guard9840;
wire _guard9842 = early_reset_static_par0_go_out;
wire _guard9843 = early_reset_static_par0_go_out;
wire _guard9844 = early_reset_static_par0_go_out;
wire _guard9845 = early_reset_static_par0_go_out;
wire _guard9846 = early_reset_static_par0_go_out;
wire _guard9847 = ~_guard0;
wire _guard9848 = early_reset_static_par0_go_out;
wire _guard9849 = _guard9847 & _guard9848;
wire _guard9850 = early_reset_static_par0_go_out;
wire _guard9851 = ~_guard0;
wire _guard9852 = early_reset_static_par0_go_out;
wire _guard9853 = _guard9851 & _guard9852;
wire _guard9854 = early_reset_static_par0_go_out;
wire _guard9855 = early_reset_static_par0_go_out;
wire _guard9856 = early_reset_static_par0_go_out;
wire _guard9857 = early_reset_static_par0_go_out;
wire _guard9858 = early_reset_static_par0_go_out;
wire _guard9859 = early_reset_static_par0_go_out;
wire _guard9860 = early_reset_static_par0_go_out;
wire _guard9861 = early_reset_static_par0_go_out;
wire _guard9862 = ~_guard0;
wire _guard9863 = early_reset_static_par0_go_out;
wire _guard9864 = _guard9862 & _guard9863;
wire _guard9865 = cond_wire_out;
wire _guard9866 = early_reset_static_par0_go_out;
wire _guard9867 = _guard9865 & _guard9866;
wire _guard9868 = cond_wire_out;
wire _guard9869 = early_reset_static_par0_go_out;
wire _guard9870 = _guard9868 & _guard9869;
wire _guard9871 = cond_wire17_out;
wire _guard9872 = early_reset_static_par0_go_out;
wire _guard9873 = _guard9871 & _guard9872;
wire _guard9874 = cond_wire15_out;
wire _guard9875 = early_reset_static_par0_go_out;
wire _guard9876 = _guard9874 & _guard9875;
wire _guard9877 = fsm_out == 1'd0;
wire _guard9878 = cond_wire15_out;
wire _guard9879 = _guard9877 & _guard9878;
wire _guard9880 = fsm_out == 1'd0;
wire _guard9881 = _guard9879 & _guard9880;
wire _guard9882 = fsm_out == 1'd0;
wire _guard9883 = cond_wire17_out;
wire _guard9884 = _guard9882 & _guard9883;
wire _guard9885 = fsm_out == 1'd0;
wire _guard9886 = _guard9884 & _guard9885;
wire _guard9887 = _guard9881 | _guard9886;
wire _guard9888 = early_reset_static_par0_go_out;
wire _guard9889 = _guard9887 & _guard9888;
wire _guard9890 = fsm_out == 1'd0;
wire _guard9891 = cond_wire15_out;
wire _guard9892 = _guard9890 & _guard9891;
wire _guard9893 = fsm_out == 1'd0;
wire _guard9894 = _guard9892 & _guard9893;
wire _guard9895 = fsm_out == 1'd0;
wire _guard9896 = cond_wire17_out;
wire _guard9897 = _guard9895 & _guard9896;
wire _guard9898 = fsm_out == 1'd0;
wire _guard9899 = _guard9897 & _guard9898;
wire _guard9900 = _guard9894 | _guard9899;
wire _guard9901 = early_reset_static_par0_go_out;
wire _guard9902 = _guard9900 & _guard9901;
wire _guard9903 = fsm_out == 1'd0;
wire _guard9904 = cond_wire15_out;
wire _guard9905 = _guard9903 & _guard9904;
wire _guard9906 = fsm_out == 1'd0;
wire _guard9907 = _guard9905 & _guard9906;
wire _guard9908 = fsm_out == 1'd0;
wire _guard9909 = cond_wire17_out;
wire _guard9910 = _guard9908 & _guard9909;
wire _guard9911 = fsm_out == 1'd0;
wire _guard9912 = _guard9910 & _guard9911;
wire _guard9913 = _guard9907 | _guard9912;
wire _guard9914 = early_reset_static_par0_go_out;
wire _guard9915 = _guard9913 & _guard9914;
wire _guard9916 = cond_wire27_out;
wire _guard9917 = early_reset_static_par0_go_out;
wire _guard9918 = _guard9916 & _guard9917;
wire _guard9919 = cond_wire25_out;
wire _guard9920 = early_reset_static_par0_go_out;
wire _guard9921 = _guard9919 & _guard9920;
wire _guard9922 = fsm_out == 1'd0;
wire _guard9923 = cond_wire25_out;
wire _guard9924 = _guard9922 & _guard9923;
wire _guard9925 = fsm_out == 1'd0;
wire _guard9926 = _guard9924 & _guard9925;
wire _guard9927 = fsm_out == 1'd0;
wire _guard9928 = cond_wire27_out;
wire _guard9929 = _guard9927 & _guard9928;
wire _guard9930 = fsm_out == 1'd0;
wire _guard9931 = _guard9929 & _guard9930;
wire _guard9932 = _guard9926 | _guard9931;
wire _guard9933 = early_reset_static_par0_go_out;
wire _guard9934 = _guard9932 & _guard9933;
wire _guard9935 = fsm_out == 1'd0;
wire _guard9936 = cond_wire25_out;
wire _guard9937 = _guard9935 & _guard9936;
wire _guard9938 = fsm_out == 1'd0;
wire _guard9939 = _guard9937 & _guard9938;
wire _guard9940 = fsm_out == 1'd0;
wire _guard9941 = cond_wire27_out;
wire _guard9942 = _guard9940 & _guard9941;
wire _guard9943 = fsm_out == 1'd0;
wire _guard9944 = _guard9942 & _guard9943;
wire _guard9945 = _guard9939 | _guard9944;
wire _guard9946 = early_reset_static_par0_go_out;
wire _guard9947 = _guard9945 & _guard9946;
wire _guard9948 = fsm_out == 1'd0;
wire _guard9949 = cond_wire25_out;
wire _guard9950 = _guard9948 & _guard9949;
wire _guard9951 = fsm_out == 1'd0;
wire _guard9952 = _guard9950 & _guard9951;
wire _guard9953 = fsm_out == 1'd0;
wire _guard9954 = cond_wire27_out;
wire _guard9955 = _guard9953 & _guard9954;
wire _guard9956 = fsm_out == 1'd0;
wire _guard9957 = _guard9955 & _guard9956;
wire _guard9958 = _guard9952 | _guard9957;
wire _guard9959 = early_reset_static_par0_go_out;
wire _guard9960 = _guard9958 & _guard9959;
wire _guard9961 = cond_wire42_out;
wire _guard9962 = early_reset_static_par0_go_out;
wire _guard9963 = _guard9961 & _guard9962;
wire _guard9964 = cond_wire40_out;
wire _guard9965 = early_reset_static_par0_go_out;
wire _guard9966 = _guard9964 & _guard9965;
wire _guard9967 = fsm_out == 1'd0;
wire _guard9968 = cond_wire40_out;
wire _guard9969 = _guard9967 & _guard9968;
wire _guard9970 = fsm_out == 1'd0;
wire _guard9971 = _guard9969 & _guard9970;
wire _guard9972 = fsm_out == 1'd0;
wire _guard9973 = cond_wire42_out;
wire _guard9974 = _guard9972 & _guard9973;
wire _guard9975 = fsm_out == 1'd0;
wire _guard9976 = _guard9974 & _guard9975;
wire _guard9977 = _guard9971 | _guard9976;
wire _guard9978 = early_reset_static_par0_go_out;
wire _guard9979 = _guard9977 & _guard9978;
wire _guard9980 = fsm_out == 1'd0;
wire _guard9981 = cond_wire40_out;
wire _guard9982 = _guard9980 & _guard9981;
wire _guard9983 = fsm_out == 1'd0;
wire _guard9984 = _guard9982 & _guard9983;
wire _guard9985 = fsm_out == 1'd0;
wire _guard9986 = cond_wire42_out;
wire _guard9987 = _guard9985 & _guard9986;
wire _guard9988 = fsm_out == 1'd0;
wire _guard9989 = _guard9987 & _guard9988;
wire _guard9990 = _guard9984 | _guard9989;
wire _guard9991 = early_reset_static_par0_go_out;
wire _guard9992 = _guard9990 & _guard9991;
wire _guard9993 = fsm_out == 1'd0;
wire _guard9994 = cond_wire40_out;
wire _guard9995 = _guard9993 & _guard9994;
wire _guard9996 = fsm_out == 1'd0;
wire _guard9997 = _guard9995 & _guard9996;
wire _guard9998 = fsm_out == 1'd0;
wire _guard9999 = cond_wire42_out;
wire _guard10000 = _guard9998 & _guard9999;
wire _guard10001 = fsm_out == 1'd0;
wire _guard10002 = _guard10000 & _guard10001;
wire _guard10003 = _guard9997 | _guard10002;
wire _guard10004 = early_reset_static_par0_go_out;
wire _guard10005 = _guard10003 & _guard10004;
wire _guard10006 = cond_wire47_out;
wire _guard10007 = early_reset_static_par0_go_out;
wire _guard10008 = _guard10006 & _guard10007;
wire _guard10009 = cond_wire45_out;
wire _guard10010 = early_reset_static_par0_go_out;
wire _guard10011 = _guard10009 & _guard10010;
wire _guard10012 = fsm_out == 1'd0;
wire _guard10013 = cond_wire45_out;
wire _guard10014 = _guard10012 & _guard10013;
wire _guard10015 = fsm_out == 1'd0;
wire _guard10016 = _guard10014 & _guard10015;
wire _guard10017 = fsm_out == 1'd0;
wire _guard10018 = cond_wire47_out;
wire _guard10019 = _guard10017 & _guard10018;
wire _guard10020 = fsm_out == 1'd0;
wire _guard10021 = _guard10019 & _guard10020;
wire _guard10022 = _guard10016 | _guard10021;
wire _guard10023 = early_reset_static_par0_go_out;
wire _guard10024 = _guard10022 & _guard10023;
wire _guard10025 = fsm_out == 1'd0;
wire _guard10026 = cond_wire45_out;
wire _guard10027 = _guard10025 & _guard10026;
wire _guard10028 = fsm_out == 1'd0;
wire _guard10029 = _guard10027 & _guard10028;
wire _guard10030 = fsm_out == 1'd0;
wire _guard10031 = cond_wire47_out;
wire _guard10032 = _guard10030 & _guard10031;
wire _guard10033 = fsm_out == 1'd0;
wire _guard10034 = _guard10032 & _guard10033;
wire _guard10035 = _guard10029 | _guard10034;
wire _guard10036 = early_reset_static_par0_go_out;
wire _guard10037 = _guard10035 & _guard10036;
wire _guard10038 = fsm_out == 1'd0;
wire _guard10039 = cond_wire45_out;
wire _guard10040 = _guard10038 & _guard10039;
wire _guard10041 = fsm_out == 1'd0;
wire _guard10042 = _guard10040 & _guard10041;
wire _guard10043 = fsm_out == 1'd0;
wire _guard10044 = cond_wire47_out;
wire _guard10045 = _guard10043 & _guard10044;
wire _guard10046 = fsm_out == 1'd0;
wire _guard10047 = _guard10045 & _guard10046;
wire _guard10048 = _guard10042 | _guard10047;
wire _guard10049 = early_reset_static_par0_go_out;
wire _guard10050 = _guard10048 & _guard10049;
wire _guard10051 = cond_wire59_out;
wire _guard10052 = early_reset_static_par0_go_out;
wire _guard10053 = _guard10051 & _guard10052;
wire _guard10054 = cond_wire59_out;
wire _guard10055 = early_reset_static_par0_go_out;
wire _guard10056 = _guard10054 & _guard10055;
wire _guard10057 = cond_wire16_out;
wire _guard10058 = early_reset_static_par0_go_out;
wire _guard10059 = _guard10057 & _guard10058;
wire _guard10060 = cond_wire16_out;
wire _guard10061 = early_reset_static_par0_go_out;
wire _guard10062 = _guard10060 & _guard10061;
wire _guard10063 = cond_wire21_out;
wire _guard10064 = early_reset_static_par0_go_out;
wire _guard10065 = _guard10063 & _guard10064;
wire _guard10066 = cond_wire21_out;
wire _guard10067 = early_reset_static_par0_go_out;
wire _guard10068 = _guard10066 & _guard10067;
wire _guard10069 = cond_wire41_out;
wire _guard10070 = early_reset_static_par0_go_out;
wire _guard10071 = _guard10069 & _guard10070;
wire _guard10072 = cond_wire41_out;
wire _guard10073 = early_reset_static_par0_go_out;
wire _guard10074 = _guard10072 & _guard10073;
wire _guard10075 = cond_wire154_out;
wire _guard10076 = early_reset_static_par0_go_out;
wire _guard10077 = _guard10075 & _guard10076;
wire _guard10078 = cond_wire154_out;
wire _guard10079 = early_reset_static_par0_go_out;
wire _guard10080 = _guard10078 & _guard10079;
wire _guard10081 = cond_wire163_out;
wire _guard10082 = early_reset_static_par0_go_out;
wire _guard10083 = _guard10081 & _guard10082;
wire _guard10084 = cond_wire161_out;
wire _guard10085 = early_reset_static_par0_go_out;
wire _guard10086 = _guard10084 & _guard10085;
wire _guard10087 = fsm_out == 1'd0;
wire _guard10088 = cond_wire161_out;
wire _guard10089 = _guard10087 & _guard10088;
wire _guard10090 = fsm_out == 1'd0;
wire _guard10091 = _guard10089 & _guard10090;
wire _guard10092 = fsm_out == 1'd0;
wire _guard10093 = cond_wire163_out;
wire _guard10094 = _guard10092 & _guard10093;
wire _guard10095 = fsm_out == 1'd0;
wire _guard10096 = _guard10094 & _guard10095;
wire _guard10097 = _guard10091 | _guard10096;
wire _guard10098 = early_reset_static_par0_go_out;
wire _guard10099 = _guard10097 & _guard10098;
wire _guard10100 = fsm_out == 1'd0;
wire _guard10101 = cond_wire161_out;
wire _guard10102 = _guard10100 & _guard10101;
wire _guard10103 = fsm_out == 1'd0;
wire _guard10104 = _guard10102 & _guard10103;
wire _guard10105 = fsm_out == 1'd0;
wire _guard10106 = cond_wire163_out;
wire _guard10107 = _guard10105 & _guard10106;
wire _guard10108 = fsm_out == 1'd0;
wire _guard10109 = _guard10107 & _guard10108;
wire _guard10110 = _guard10104 | _guard10109;
wire _guard10111 = early_reset_static_par0_go_out;
wire _guard10112 = _guard10110 & _guard10111;
wire _guard10113 = fsm_out == 1'd0;
wire _guard10114 = cond_wire161_out;
wire _guard10115 = _guard10113 & _guard10114;
wire _guard10116 = fsm_out == 1'd0;
wire _guard10117 = _guard10115 & _guard10116;
wire _guard10118 = fsm_out == 1'd0;
wire _guard10119 = cond_wire163_out;
wire _guard10120 = _guard10118 & _guard10119;
wire _guard10121 = fsm_out == 1'd0;
wire _guard10122 = _guard10120 & _guard10121;
wire _guard10123 = _guard10117 | _guard10122;
wire _guard10124 = early_reset_static_par0_go_out;
wire _guard10125 = _guard10123 & _guard10124;
wire _guard10126 = cond_wire105_out;
wire _guard10127 = early_reset_static_par0_go_out;
wire _guard10128 = _guard10126 & _guard10127;
wire _guard10129 = cond_wire105_out;
wire _guard10130 = early_reset_static_par0_go_out;
wire _guard10131 = _guard10129 & _guard10130;
wire _guard10132 = cond_wire125_out;
wire _guard10133 = early_reset_static_par0_go_out;
wire _guard10134 = _guard10132 & _guard10133;
wire _guard10135 = cond_wire125_out;
wire _guard10136 = early_reset_static_par0_go_out;
wire _guard10137 = _guard10135 & _guard10136;
wire _guard10138 = cond_wire207_out;
wire _guard10139 = early_reset_static_par0_go_out;
wire _guard10140 = _guard10138 & _guard10139;
wire _guard10141 = cond_wire205_out;
wire _guard10142 = early_reset_static_par0_go_out;
wire _guard10143 = _guard10141 & _guard10142;
wire _guard10144 = fsm_out == 1'd0;
wire _guard10145 = cond_wire205_out;
wire _guard10146 = _guard10144 & _guard10145;
wire _guard10147 = fsm_out == 1'd0;
wire _guard10148 = _guard10146 & _guard10147;
wire _guard10149 = fsm_out == 1'd0;
wire _guard10150 = cond_wire207_out;
wire _guard10151 = _guard10149 & _guard10150;
wire _guard10152 = fsm_out == 1'd0;
wire _guard10153 = _guard10151 & _guard10152;
wire _guard10154 = _guard10148 | _guard10153;
wire _guard10155 = early_reset_static_par0_go_out;
wire _guard10156 = _guard10154 & _guard10155;
wire _guard10157 = fsm_out == 1'd0;
wire _guard10158 = cond_wire205_out;
wire _guard10159 = _guard10157 & _guard10158;
wire _guard10160 = fsm_out == 1'd0;
wire _guard10161 = _guard10159 & _guard10160;
wire _guard10162 = fsm_out == 1'd0;
wire _guard10163 = cond_wire207_out;
wire _guard10164 = _guard10162 & _guard10163;
wire _guard10165 = fsm_out == 1'd0;
wire _guard10166 = _guard10164 & _guard10165;
wire _guard10167 = _guard10161 | _guard10166;
wire _guard10168 = early_reset_static_par0_go_out;
wire _guard10169 = _guard10167 & _guard10168;
wire _guard10170 = fsm_out == 1'd0;
wire _guard10171 = cond_wire205_out;
wire _guard10172 = _guard10170 & _guard10171;
wire _guard10173 = fsm_out == 1'd0;
wire _guard10174 = _guard10172 & _guard10173;
wire _guard10175 = fsm_out == 1'd0;
wire _guard10176 = cond_wire207_out;
wire _guard10177 = _guard10175 & _guard10176;
wire _guard10178 = fsm_out == 1'd0;
wire _guard10179 = _guard10177 & _guard10178;
wire _guard10180 = _guard10174 | _guard10179;
wire _guard10181 = early_reset_static_par0_go_out;
wire _guard10182 = _guard10180 & _guard10181;
wire _guard10183 = cond_wire212_out;
wire _guard10184 = early_reset_static_par0_go_out;
wire _guard10185 = _guard10183 & _guard10184;
wire _guard10186 = cond_wire210_out;
wire _guard10187 = early_reset_static_par0_go_out;
wire _guard10188 = _guard10186 & _guard10187;
wire _guard10189 = fsm_out == 1'd0;
wire _guard10190 = cond_wire210_out;
wire _guard10191 = _guard10189 & _guard10190;
wire _guard10192 = fsm_out == 1'd0;
wire _guard10193 = _guard10191 & _guard10192;
wire _guard10194 = fsm_out == 1'd0;
wire _guard10195 = cond_wire212_out;
wire _guard10196 = _guard10194 & _guard10195;
wire _guard10197 = fsm_out == 1'd0;
wire _guard10198 = _guard10196 & _guard10197;
wire _guard10199 = _guard10193 | _guard10198;
wire _guard10200 = early_reset_static_par0_go_out;
wire _guard10201 = _guard10199 & _guard10200;
wire _guard10202 = fsm_out == 1'd0;
wire _guard10203 = cond_wire210_out;
wire _guard10204 = _guard10202 & _guard10203;
wire _guard10205 = fsm_out == 1'd0;
wire _guard10206 = _guard10204 & _guard10205;
wire _guard10207 = fsm_out == 1'd0;
wire _guard10208 = cond_wire212_out;
wire _guard10209 = _guard10207 & _guard10208;
wire _guard10210 = fsm_out == 1'd0;
wire _guard10211 = _guard10209 & _guard10210;
wire _guard10212 = _guard10206 | _guard10211;
wire _guard10213 = early_reset_static_par0_go_out;
wire _guard10214 = _guard10212 & _guard10213;
wire _guard10215 = fsm_out == 1'd0;
wire _guard10216 = cond_wire210_out;
wire _guard10217 = _guard10215 & _guard10216;
wire _guard10218 = fsm_out == 1'd0;
wire _guard10219 = _guard10217 & _guard10218;
wire _guard10220 = fsm_out == 1'd0;
wire _guard10221 = cond_wire212_out;
wire _guard10222 = _guard10220 & _guard10221;
wire _guard10223 = fsm_out == 1'd0;
wire _guard10224 = _guard10222 & _guard10223;
wire _guard10225 = _guard10219 | _guard10224;
wire _guard10226 = early_reset_static_par0_go_out;
wire _guard10227 = _guard10225 & _guard10226;
wire _guard10228 = cond_wire154_out;
wire _guard10229 = early_reset_static_par0_go_out;
wire _guard10230 = _guard10228 & _guard10229;
wire _guard10231 = cond_wire154_out;
wire _guard10232 = early_reset_static_par0_go_out;
wire _guard10233 = _guard10231 & _guard10232;
wire _guard10234 = cond_wire202_out;
wire _guard10235 = early_reset_static_par0_go_out;
wire _guard10236 = _guard10234 & _guard10235;
wire _guard10237 = cond_wire202_out;
wire _guard10238 = early_reset_static_par0_go_out;
wire _guard10239 = _guard10237 & _guard10238;
wire _guard10240 = cond_wire211_out;
wire _guard10241 = early_reset_static_par0_go_out;
wire _guard10242 = _guard10240 & _guard10241;
wire _guard10243 = cond_wire211_out;
wire _guard10244 = early_reset_static_par0_go_out;
wire _guard10245 = _guard10243 & _guard10244;
wire _guard10246 = cond_wire296_out;
wire _guard10247 = early_reset_static_par0_go_out;
wire _guard10248 = _guard10246 & _guard10247;
wire _guard10249 = cond_wire296_out;
wire _guard10250 = early_reset_static_par0_go_out;
wire _guard10251 = _guard10249 & _guard10250;
wire _guard10252 = cond_wire300_out;
wire _guard10253 = early_reset_static_par0_go_out;
wire _guard10254 = _guard10252 & _guard10253;
wire _guard10255 = cond_wire300_out;
wire _guard10256 = early_reset_static_par0_go_out;
wire _guard10257 = _guard10255 & _guard10256;
wire _guard10258 = cond_wire346_out;
wire _guard10259 = early_reset_static_par0_go_out;
wire _guard10260 = _guard10258 & _guard10259;
wire _guard10261 = cond_wire344_out;
wire _guard10262 = early_reset_static_par0_go_out;
wire _guard10263 = _guard10261 & _guard10262;
wire _guard10264 = fsm_out == 1'd0;
wire _guard10265 = cond_wire344_out;
wire _guard10266 = _guard10264 & _guard10265;
wire _guard10267 = fsm_out == 1'd0;
wire _guard10268 = _guard10266 & _guard10267;
wire _guard10269 = fsm_out == 1'd0;
wire _guard10270 = cond_wire346_out;
wire _guard10271 = _guard10269 & _guard10270;
wire _guard10272 = fsm_out == 1'd0;
wire _guard10273 = _guard10271 & _guard10272;
wire _guard10274 = _guard10268 | _guard10273;
wire _guard10275 = early_reset_static_par0_go_out;
wire _guard10276 = _guard10274 & _guard10275;
wire _guard10277 = fsm_out == 1'd0;
wire _guard10278 = cond_wire344_out;
wire _guard10279 = _guard10277 & _guard10278;
wire _guard10280 = fsm_out == 1'd0;
wire _guard10281 = _guard10279 & _guard10280;
wire _guard10282 = fsm_out == 1'd0;
wire _guard10283 = cond_wire346_out;
wire _guard10284 = _guard10282 & _guard10283;
wire _guard10285 = fsm_out == 1'd0;
wire _guard10286 = _guard10284 & _guard10285;
wire _guard10287 = _guard10281 | _guard10286;
wire _guard10288 = early_reset_static_par0_go_out;
wire _guard10289 = _guard10287 & _guard10288;
wire _guard10290 = fsm_out == 1'd0;
wire _guard10291 = cond_wire344_out;
wire _guard10292 = _guard10290 & _guard10291;
wire _guard10293 = fsm_out == 1'd0;
wire _guard10294 = _guard10292 & _guard10293;
wire _guard10295 = fsm_out == 1'd0;
wire _guard10296 = cond_wire346_out;
wire _guard10297 = _guard10295 & _guard10296;
wire _guard10298 = fsm_out == 1'd0;
wire _guard10299 = _guard10297 & _guard10298;
wire _guard10300 = _guard10294 | _guard10299;
wire _guard10301 = early_reset_static_par0_go_out;
wire _guard10302 = _guard10300 & _guard10301;
wire _guard10303 = cond_wire370_out;
wire _guard10304 = early_reset_static_par0_go_out;
wire _guard10305 = _guard10303 & _guard10304;
wire _guard10306 = cond_wire368_out;
wire _guard10307 = early_reset_static_par0_go_out;
wire _guard10308 = _guard10306 & _guard10307;
wire _guard10309 = fsm_out == 1'd0;
wire _guard10310 = cond_wire368_out;
wire _guard10311 = _guard10309 & _guard10310;
wire _guard10312 = fsm_out == 1'd0;
wire _guard10313 = _guard10311 & _guard10312;
wire _guard10314 = fsm_out == 1'd0;
wire _guard10315 = cond_wire370_out;
wire _guard10316 = _guard10314 & _guard10315;
wire _guard10317 = fsm_out == 1'd0;
wire _guard10318 = _guard10316 & _guard10317;
wire _guard10319 = _guard10313 | _guard10318;
wire _guard10320 = early_reset_static_par0_go_out;
wire _guard10321 = _guard10319 & _guard10320;
wire _guard10322 = fsm_out == 1'd0;
wire _guard10323 = cond_wire368_out;
wire _guard10324 = _guard10322 & _guard10323;
wire _guard10325 = fsm_out == 1'd0;
wire _guard10326 = _guard10324 & _guard10325;
wire _guard10327 = fsm_out == 1'd0;
wire _guard10328 = cond_wire370_out;
wire _guard10329 = _guard10327 & _guard10328;
wire _guard10330 = fsm_out == 1'd0;
wire _guard10331 = _guard10329 & _guard10330;
wire _guard10332 = _guard10326 | _guard10331;
wire _guard10333 = early_reset_static_par0_go_out;
wire _guard10334 = _guard10332 & _guard10333;
wire _guard10335 = fsm_out == 1'd0;
wire _guard10336 = cond_wire368_out;
wire _guard10337 = _guard10335 & _guard10336;
wire _guard10338 = fsm_out == 1'd0;
wire _guard10339 = _guard10337 & _guard10338;
wire _guard10340 = fsm_out == 1'd0;
wire _guard10341 = cond_wire370_out;
wire _guard10342 = _guard10340 & _guard10341;
wire _guard10343 = fsm_out == 1'd0;
wire _guard10344 = _guard10342 & _guard10343;
wire _guard10345 = _guard10339 | _guard10344;
wire _guard10346 = early_reset_static_par0_go_out;
wire _guard10347 = _guard10345 & _guard10346;
wire _guard10348 = cond_wire407_out;
wire _guard10349 = early_reset_static_par0_go_out;
wire _guard10350 = _guard10348 & _guard10349;
wire _guard10351 = cond_wire405_out;
wire _guard10352 = early_reset_static_par0_go_out;
wire _guard10353 = _guard10351 & _guard10352;
wire _guard10354 = fsm_out == 1'd0;
wire _guard10355 = cond_wire405_out;
wire _guard10356 = _guard10354 & _guard10355;
wire _guard10357 = fsm_out == 1'd0;
wire _guard10358 = _guard10356 & _guard10357;
wire _guard10359 = fsm_out == 1'd0;
wire _guard10360 = cond_wire407_out;
wire _guard10361 = _guard10359 & _guard10360;
wire _guard10362 = fsm_out == 1'd0;
wire _guard10363 = _guard10361 & _guard10362;
wire _guard10364 = _guard10358 | _guard10363;
wire _guard10365 = early_reset_static_par0_go_out;
wire _guard10366 = _guard10364 & _guard10365;
wire _guard10367 = fsm_out == 1'd0;
wire _guard10368 = cond_wire405_out;
wire _guard10369 = _guard10367 & _guard10368;
wire _guard10370 = fsm_out == 1'd0;
wire _guard10371 = _guard10369 & _guard10370;
wire _guard10372 = fsm_out == 1'd0;
wire _guard10373 = cond_wire407_out;
wire _guard10374 = _guard10372 & _guard10373;
wire _guard10375 = fsm_out == 1'd0;
wire _guard10376 = _guard10374 & _guard10375;
wire _guard10377 = _guard10371 | _guard10376;
wire _guard10378 = early_reset_static_par0_go_out;
wire _guard10379 = _guard10377 & _guard10378;
wire _guard10380 = fsm_out == 1'd0;
wire _guard10381 = cond_wire405_out;
wire _guard10382 = _guard10380 & _guard10381;
wire _guard10383 = fsm_out == 1'd0;
wire _guard10384 = _guard10382 & _guard10383;
wire _guard10385 = fsm_out == 1'd0;
wire _guard10386 = cond_wire407_out;
wire _guard10387 = _guard10385 & _guard10386;
wire _guard10388 = fsm_out == 1'd0;
wire _guard10389 = _guard10387 & _guard10388;
wire _guard10390 = _guard10384 | _guard10389;
wire _guard10391 = early_reset_static_par0_go_out;
wire _guard10392 = _guard10390 & _guard10391;
wire _guard10393 = cond_wire341_out;
wire _guard10394 = early_reset_static_par0_go_out;
wire _guard10395 = _guard10393 & _guard10394;
wire _guard10396 = cond_wire341_out;
wire _guard10397 = early_reset_static_par0_go_out;
wire _guard10398 = _guard10396 & _guard10397;
wire _guard10399 = cond_wire411_out;
wire _guard10400 = early_reset_static_par0_go_out;
wire _guard10401 = _guard10399 & _guard10400;
wire _guard10402 = cond_wire409_out;
wire _guard10403 = early_reset_static_par0_go_out;
wire _guard10404 = _guard10402 & _guard10403;
wire _guard10405 = fsm_out == 1'd0;
wire _guard10406 = cond_wire409_out;
wire _guard10407 = _guard10405 & _guard10406;
wire _guard10408 = fsm_out == 1'd0;
wire _guard10409 = _guard10407 & _guard10408;
wire _guard10410 = fsm_out == 1'd0;
wire _guard10411 = cond_wire411_out;
wire _guard10412 = _guard10410 & _guard10411;
wire _guard10413 = fsm_out == 1'd0;
wire _guard10414 = _guard10412 & _guard10413;
wire _guard10415 = _guard10409 | _guard10414;
wire _guard10416 = early_reset_static_par0_go_out;
wire _guard10417 = _guard10415 & _guard10416;
wire _guard10418 = fsm_out == 1'd0;
wire _guard10419 = cond_wire409_out;
wire _guard10420 = _guard10418 & _guard10419;
wire _guard10421 = fsm_out == 1'd0;
wire _guard10422 = _guard10420 & _guard10421;
wire _guard10423 = fsm_out == 1'd0;
wire _guard10424 = cond_wire411_out;
wire _guard10425 = _guard10423 & _guard10424;
wire _guard10426 = fsm_out == 1'd0;
wire _guard10427 = _guard10425 & _guard10426;
wire _guard10428 = _guard10422 | _guard10427;
wire _guard10429 = early_reset_static_par0_go_out;
wire _guard10430 = _guard10428 & _guard10429;
wire _guard10431 = fsm_out == 1'd0;
wire _guard10432 = cond_wire409_out;
wire _guard10433 = _guard10431 & _guard10432;
wire _guard10434 = fsm_out == 1'd0;
wire _guard10435 = _guard10433 & _guard10434;
wire _guard10436 = fsm_out == 1'd0;
wire _guard10437 = cond_wire411_out;
wire _guard10438 = _guard10436 & _guard10437;
wire _guard10439 = fsm_out == 1'd0;
wire _guard10440 = _guard10438 & _guard10439;
wire _guard10441 = _guard10435 | _guard10440;
wire _guard10442 = early_reset_static_par0_go_out;
wire _guard10443 = _guard10441 & _guard10442;
wire _guard10444 = cond_wire446_out;
wire _guard10445 = early_reset_static_par0_go_out;
wire _guard10446 = _guard10444 & _guard10445;
wire _guard10447 = cond_wire446_out;
wire _guard10448 = early_reset_static_par0_go_out;
wire _guard10449 = _guard10447 & _guard10448;
wire _guard10450 = cond_wire487_out;
wire _guard10451 = early_reset_static_par0_go_out;
wire _guard10452 = _guard10450 & _guard10451;
wire _guard10453 = cond_wire487_out;
wire _guard10454 = early_reset_static_par0_go_out;
wire _guard10455 = _guard10453 & _guard10454;
wire _guard10456 = cond_wire545_out;
wire _guard10457 = early_reset_static_par0_go_out;
wire _guard10458 = _guard10456 & _guard10457;
wire _guard10459 = cond_wire543_out;
wire _guard10460 = early_reset_static_par0_go_out;
wire _guard10461 = _guard10459 & _guard10460;
wire _guard10462 = fsm_out == 1'd0;
wire _guard10463 = cond_wire543_out;
wire _guard10464 = _guard10462 & _guard10463;
wire _guard10465 = fsm_out == 1'd0;
wire _guard10466 = _guard10464 & _guard10465;
wire _guard10467 = fsm_out == 1'd0;
wire _guard10468 = cond_wire545_out;
wire _guard10469 = _guard10467 & _guard10468;
wire _guard10470 = fsm_out == 1'd0;
wire _guard10471 = _guard10469 & _guard10470;
wire _guard10472 = _guard10466 | _guard10471;
wire _guard10473 = early_reset_static_par0_go_out;
wire _guard10474 = _guard10472 & _guard10473;
wire _guard10475 = fsm_out == 1'd0;
wire _guard10476 = cond_wire543_out;
wire _guard10477 = _guard10475 & _guard10476;
wire _guard10478 = fsm_out == 1'd0;
wire _guard10479 = _guard10477 & _guard10478;
wire _guard10480 = fsm_out == 1'd0;
wire _guard10481 = cond_wire545_out;
wire _guard10482 = _guard10480 & _guard10481;
wire _guard10483 = fsm_out == 1'd0;
wire _guard10484 = _guard10482 & _guard10483;
wire _guard10485 = _guard10479 | _guard10484;
wire _guard10486 = early_reset_static_par0_go_out;
wire _guard10487 = _guard10485 & _guard10486;
wire _guard10488 = fsm_out == 1'd0;
wire _guard10489 = cond_wire543_out;
wire _guard10490 = _guard10488 & _guard10489;
wire _guard10491 = fsm_out == 1'd0;
wire _guard10492 = _guard10490 & _guard10491;
wire _guard10493 = fsm_out == 1'd0;
wire _guard10494 = cond_wire545_out;
wire _guard10495 = _guard10493 & _guard10494;
wire _guard10496 = fsm_out == 1'd0;
wire _guard10497 = _guard10495 & _guard10496;
wire _guard10498 = _guard10492 | _guard10497;
wire _guard10499 = early_reset_static_par0_go_out;
wire _guard10500 = _guard10498 & _guard10499;
wire _guard10501 = cond_wire483_out;
wire _guard10502 = early_reset_static_par0_go_out;
wire _guard10503 = _guard10501 & _guard10502;
wire _guard10504 = cond_wire483_out;
wire _guard10505 = early_reset_static_par0_go_out;
wire _guard10506 = _guard10504 & _guard10505;
wire _guard10507 = cond_wire553_out;
wire _guard10508 = early_reset_static_par0_go_out;
wire _guard10509 = _guard10507 & _guard10508;
wire _guard10510 = cond_wire551_out;
wire _guard10511 = early_reset_static_par0_go_out;
wire _guard10512 = _guard10510 & _guard10511;
wire _guard10513 = fsm_out == 1'd0;
wire _guard10514 = cond_wire551_out;
wire _guard10515 = _guard10513 & _guard10514;
wire _guard10516 = fsm_out == 1'd0;
wire _guard10517 = _guard10515 & _guard10516;
wire _guard10518 = fsm_out == 1'd0;
wire _guard10519 = cond_wire553_out;
wire _guard10520 = _guard10518 & _guard10519;
wire _guard10521 = fsm_out == 1'd0;
wire _guard10522 = _guard10520 & _guard10521;
wire _guard10523 = _guard10517 | _guard10522;
wire _guard10524 = early_reset_static_par0_go_out;
wire _guard10525 = _guard10523 & _guard10524;
wire _guard10526 = fsm_out == 1'd0;
wire _guard10527 = cond_wire551_out;
wire _guard10528 = _guard10526 & _guard10527;
wire _guard10529 = fsm_out == 1'd0;
wire _guard10530 = _guard10528 & _guard10529;
wire _guard10531 = fsm_out == 1'd0;
wire _guard10532 = cond_wire553_out;
wire _guard10533 = _guard10531 & _guard10532;
wire _guard10534 = fsm_out == 1'd0;
wire _guard10535 = _guard10533 & _guard10534;
wire _guard10536 = _guard10530 | _guard10535;
wire _guard10537 = early_reset_static_par0_go_out;
wire _guard10538 = _guard10536 & _guard10537;
wire _guard10539 = fsm_out == 1'd0;
wire _guard10540 = cond_wire551_out;
wire _guard10541 = _guard10539 & _guard10540;
wire _guard10542 = fsm_out == 1'd0;
wire _guard10543 = _guard10541 & _guard10542;
wire _guard10544 = fsm_out == 1'd0;
wire _guard10545 = cond_wire553_out;
wire _guard10546 = _guard10544 & _guard10545;
wire _guard10547 = fsm_out == 1'd0;
wire _guard10548 = _guard10546 & _guard10547;
wire _guard10549 = _guard10543 | _guard10548;
wire _guard10550 = early_reset_static_par0_go_out;
wire _guard10551 = _guard10549 & _guard10550;
wire _guard10552 = cond_wire625_out;
wire _guard10553 = early_reset_static_par0_go_out;
wire _guard10554 = _guard10552 & _guard10553;
wire _guard10555 = cond_wire625_out;
wire _guard10556 = early_reset_static_par0_go_out;
wire _guard10557 = _guard10555 & _guard10556;
wire _guard10558 = cond_wire698_out;
wire _guard10559 = early_reset_static_par0_go_out;
wire _guard10560 = _guard10558 & _guard10559;
wire _guard10561 = cond_wire698_out;
wire _guard10562 = early_reset_static_par0_go_out;
wire _guard10563 = _guard10561 & _guard10562;
wire _guard10564 = cond_wire732_out;
wire _guard10565 = early_reset_static_par0_go_out;
wire _guard10566 = _guard10564 & _guard10565;
wire _guard10567 = cond_wire730_out;
wire _guard10568 = early_reset_static_par0_go_out;
wire _guard10569 = _guard10567 & _guard10568;
wire _guard10570 = fsm_out == 1'd0;
wire _guard10571 = cond_wire730_out;
wire _guard10572 = _guard10570 & _guard10571;
wire _guard10573 = fsm_out == 1'd0;
wire _guard10574 = _guard10572 & _guard10573;
wire _guard10575 = fsm_out == 1'd0;
wire _guard10576 = cond_wire732_out;
wire _guard10577 = _guard10575 & _guard10576;
wire _guard10578 = fsm_out == 1'd0;
wire _guard10579 = _guard10577 & _guard10578;
wire _guard10580 = _guard10574 | _guard10579;
wire _guard10581 = early_reset_static_par0_go_out;
wire _guard10582 = _guard10580 & _guard10581;
wire _guard10583 = fsm_out == 1'd0;
wire _guard10584 = cond_wire730_out;
wire _guard10585 = _guard10583 & _guard10584;
wire _guard10586 = fsm_out == 1'd0;
wire _guard10587 = _guard10585 & _guard10586;
wire _guard10588 = fsm_out == 1'd0;
wire _guard10589 = cond_wire732_out;
wire _guard10590 = _guard10588 & _guard10589;
wire _guard10591 = fsm_out == 1'd0;
wire _guard10592 = _guard10590 & _guard10591;
wire _guard10593 = _guard10587 | _guard10592;
wire _guard10594 = early_reset_static_par0_go_out;
wire _guard10595 = _guard10593 & _guard10594;
wire _guard10596 = fsm_out == 1'd0;
wire _guard10597 = cond_wire730_out;
wire _guard10598 = _guard10596 & _guard10597;
wire _guard10599 = fsm_out == 1'd0;
wire _guard10600 = _guard10598 & _guard10599;
wire _guard10601 = fsm_out == 1'd0;
wire _guard10602 = cond_wire732_out;
wire _guard10603 = _guard10601 & _guard10602;
wire _guard10604 = fsm_out == 1'd0;
wire _guard10605 = _guard10603 & _guard10604;
wire _guard10606 = _guard10600 | _guard10605;
wire _guard10607 = early_reset_static_par0_go_out;
wire _guard10608 = _guard10606 & _guard10607;
wire _guard10609 = cond_wire678_out;
wire _guard10610 = early_reset_static_par0_go_out;
wire _guard10611 = _guard10609 & _guard10610;
wire _guard10612 = cond_wire678_out;
wire _guard10613 = early_reset_static_par0_go_out;
wire _guard10614 = _guard10612 & _guard10613;
wire _guard10615 = cond_wire686_out;
wire _guard10616 = early_reset_static_par0_go_out;
wire _guard10617 = _guard10615 & _guard10616;
wire _guard10618 = cond_wire686_out;
wire _guard10619 = early_reset_static_par0_go_out;
wire _guard10620 = _guard10618 & _guard10619;
wire _guard10621 = cond_wire776_out;
wire _guard10622 = early_reset_static_par0_go_out;
wire _guard10623 = _guard10621 & _guard10622;
wire _guard10624 = cond_wire774_out;
wire _guard10625 = early_reset_static_par0_go_out;
wire _guard10626 = _guard10624 & _guard10625;
wire _guard10627 = fsm_out == 1'd0;
wire _guard10628 = cond_wire774_out;
wire _guard10629 = _guard10627 & _guard10628;
wire _guard10630 = fsm_out == 1'd0;
wire _guard10631 = _guard10629 & _guard10630;
wire _guard10632 = fsm_out == 1'd0;
wire _guard10633 = cond_wire776_out;
wire _guard10634 = _guard10632 & _guard10633;
wire _guard10635 = fsm_out == 1'd0;
wire _guard10636 = _guard10634 & _guard10635;
wire _guard10637 = _guard10631 | _guard10636;
wire _guard10638 = early_reset_static_par0_go_out;
wire _guard10639 = _guard10637 & _guard10638;
wire _guard10640 = fsm_out == 1'd0;
wire _guard10641 = cond_wire774_out;
wire _guard10642 = _guard10640 & _guard10641;
wire _guard10643 = fsm_out == 1'd0;
wire _guard10644 = _guard10642 & _guard10643;
wire _guard10645 = fsm_out == 1'd0;
wire _guard10646 = cond_wire776_out;
wire _guard10647 = _guard10645 & _guard10646;
wire _guard10648 = fsm_out == 1'd0;
wire _guard10649 = _guard10647 & _guard10648;
wire _guard10650 = _guard10644 | _guard10649;
wire _guard10651 = early_reset_static_par0_go_out;
wire _guard10652 = _guard10650 & _guard10651;
wire _guard10653 = fsm_out == 1'd0;
wire _guard10654 = cond_wire774_out;
wire _guard10655 = _guard10653 & _guard10654;
wire _guard10656 = fsm_out == 1'd0;
wire _guard10657 = _guard10655 & _guard10656;
wire _guard10658 = fsm_out == 1'd0;
wire _guard10659 = cond_wire776_out;
wire _guard10660 = _guard10658 & _guard10659;
wire _guard10661 = fsm_out == 1'd0;
wire _guard10662 = _guard10660 & _guard10661;
wire _guard10663 = _guard10657 | _guard10662;
wire _guard10664 = early_reset_static_par0_go_out;
wire _guard10665 = _guard10663 & _guard10664;
wire _guard10666 = cond_wire787_out;
wire _guard10667 = early_reset_static_par0_go_out;
wire _guard10668 = _guard10666 & _guard10667;
wire _guard10669 = cond_wire787_out;
wire _guard10670 = early_reset_static_par0_go_out;
wire _guard10671 = _guard10669 & _guard10670;
wire _guard10672 = cond_wire731_out;
wire _guard10673 = early_reset_static_par0_go_out;
wire _guard10674 = _guard10672 & _guard10673;
wire _guard10675 = cond_wire731_out;
wire _guard10676 = early_reset_static_par0_go_out;
wire _guard10677 = _guard10675 & _guard10676;
wire _guard10678 = cond_wire739_out;
wire _guard10679 = early_reset_static_par0_go_out;
wire _guard10680 = _guard10678 & _guard10679;
wire _guard10681 = cond_wire739_out;
wire _guard10682 = early_reset_static_par0_go_out;
wire _guard10683 = _guard10681 & _guard10682;
wire _guard10684 = cond_wire759_out;
wire _guard10685 = early_reset_static_par0_go_out;
wire _guard10686 = _guard10684 & _guard10685;
wire _guard10687 = cond_wire759_out;
wire _guard10688 = early_reset_static_par0_go_out;
wire _guard10689 = _guard10687 & _guard10688;
wire _guard10690 = cond_wire824_out;
wire _guard10691 = early_reset_static_par0_go_out;
wire _guard10692 = _guard10690 & _guard10691;
wire _guard10693 = cond_wire824_out;
wire _guard10694 = early_reset_static_par0_go_out;
wire _guard10695 = _guard10693 & _guard10694;
wire _guard10696 = cond_wire812_out;
wire _guard10697 = early_reset_static_par0_go_out;
wire _guard10698 = _guard10696 & _guard10697;
wire _guard10699 = cond_wire812_out;
wire _guard10700 = early_reset_static_par0_go_out;
wire _guard10701 = _guard10699 & _guard10700;
wire _guard10702 = cond_wire832_out;
wire _guard10703 = early_reset_static_par0_go_out;
wire _guard10704 = _guard10702 & _guard10703;
wire _guard10705 = cond_wire832_out;
wire _guard10706 = early_reset_static_par0_go_out;
wire _guard10707 = _guard10705 & _guard10706;
wire _guard10708 = cond_wire856_out;
wire _guard10709 = early_reset_static_par0_go_out;
wire _guard10710 = _guard10708 & _guard10709;
wire _guard10711 = cond_wire856_out;
wire _guard10712 = early_reset_static_par0_go_out;
wire _guard10713 = _guard10711 & _guard10712;
wire _guard10714 = cond_wire893_out;
wire _guard10715 = early_reset_static_par0_go_out;
wire _guard10716 = _guard10714 & _guard10715;
wire _guard10717 = cond_wire893_out;
wire _guard10718 = early_reset_static_par0_go_out;
wire _guard10719 = _guard10717 & _guard10718;
wire _guard10720 = cond_wire942_out;
wire _guard10721 = early_reset_static_par0_go_out;
wire _guard10722 = _guard10720 & _guard10721;
wire _guard10723 = cond_wire942_out;
wire _guard10724 = early_reset_static_par0_go_out;
wire _guard10725 = _guard10723 & _guard10724;
wire _guard10726 = cond_wire1027_out;
wire _guard10727 = early_reset_static_par0_go_out;
wire _guard10728 = _guard10726 & _guard10727;
wire _guard10729 = cond_wire1027_out;
wire _guard10730 = early_reset_static_par0_go_out;
wire _guard10731 = _guard10729 & _guard10730;
wire _guard10732 = cond_wire729_out;
wire _guard10733 = early_reset_static_par0_go_out;
wire _guard10734 = _guard10732 & _guard10733;
wire _guard10735 = cond_wire729_out;
wire _guard10736 = early_reset_static_par0_go_out;
wire _guard10737 = _guard10735 & _guard10736;
wire _guard10738 = early_reset_static_par0_go_out;
wire _guard10739 = early_reset_static_par0_go_out;
wire _guard10740 = early_reset_static_par0_go_out;
wire _guard10741 = early_reset_static_par0_go_out;
wire _guard10742 = fsm0_out == 6'd0;
wire _guard10743 = early_reset_static_seq_go_out;
wire _guard10744 = _guard10742 & _guard10743;
wire _guard10745 = early_reset_static_par0_go_out;
wire _guard10746 = _guard10744 | _guard10745;
wire _guard10747 = early_reset_static_par0_go_out;
wire _guard10748 = fsm0_out == 6'd0;
wire _guard10749 = early_reset_static_seq_go_out;
wire _guard10750 = _guard10748 & _guard10749;
wire _guard10751 = early_reset_static_par0_go_out;
wire _guard10752 = early_reset_static_par0_go_out;
wire _guard10753 = early_reset_static_par0_go_out;
wire _guard10754 = early_reset_static_par0_go_out;
wire _guard10755 = fsm0_out == 6'd0;
wire _guard10756 = early_reset_static_seq_go_out;
wire _guard10757 = _guard10755 & _guard10756;
wire _guard10758 = early_reset_static_par0_go_out;
wire _guard10759 = _guard10757 | _guard10758;
wire _guard10760 = early_reset_static_par0_go_out;
wire _guard10761 = fsm0_out == 6'd0;
wire _guard10762 = early_reset_static_seq_go_out;
wire _guard10763 = _guard10761 & _guard10762;
wire _guard10764 = fsm0_out == 6'd0;
wire _guard10765 = early_reset_static_seq_go_out;
wire _guard10766 = _guard10764 & _guard10765;
wire _guard10767 = early_reset_static_par0_go_out;
wire _guard10768 = _guard10766 | _guard10767;
wire _guard10769 = fsm0_out == 6'd0;
wire _guard10770 = early_reset_static_seq_go_out;
wire _guard10771 = _guard10769 & _guard10770;
wire _guard10772 = early_reset_static_par0_go_out;
wire _guard10773 = fsm0_out == 6'd0;
wire _guard10774 = early_reset_static_seq_go_out;
wire _guard10775 = _guard10773 & _guard10774;
wire _guard10776 = early_reset_static_par0_go_out;
wire _guard10777 = _guard10775 | _guard10776;
wire _guard10778 = early_reset_static_par0_go_out;
wire _guard10779 = fsm0_out == 6'd0;
wire _guard10780 = early_reset_static_seq_go_out;
wire _guard10781 = _guard10779 & _guard10780;
wire _guard10782 = early_reset_static_par0_go_out;
wire _guard10783 = early_reset_static_par0_go_out;
wire _guard10784 = early_reset_static_par0_go_out;
wire _guard10785 = early_reset_static_par0_go_out;
wire _guard10786 = early_reset_static_par0_go_out;
wire _guard10787 = early_reset_static_par0_go_out;
wire _guard10788 = fsm0_out == 6'd0;
wire _guard10789 = early_reset_static_seq_go_out;
wire _guard10790 = _guard10788 & _guard10789;
wire _guard10791 = early_reset_static_par0_go_out;
wire _guard10792 = _guard10790 | _guard10791;
wire _guard10793 = early_reset_static_par0_go_out;
wire _guard10794 = fsm0_out == 6'd0;
wire _guard10795 = early_reset_static_seq_go_out;
wire _guard10796 = _guard10794 & _guard10795;
wire _guard10797 = early_reset_static_par0_go_out;
wire _guard10798 = early_reset_static_par0_go_out;
wire _guard10799 = early_reset_static_par0_go_out;
wire _guard10800 = early_reset_static_par0_go_out;
wire _guard10801 = fsm0_out == 6'd0;
wire _guard10802 = early_reset_static_seq_go_out;
wire _guard10803 = _guard10801 & _guard10802;
wire _guard10804 = early_reset_static_par0_go_out;
wire _guard10805 = _guard10803 | _guard10804;
wire _guard10806 = fsm0_out == 6'd0;
wire _guard10807 = early_reset_static_seq_go_out;
wire _guard10808 = _guard10806 & _guard10807;
wire _guard10809 = early_reset_static_par0_go_out;
wire _guard10810 = early_reset_static_par0_go_out;
wire _guard10811 = early_reset_static_par0_go_out;
wire _guard10812 = early_reset_static_par0_go_out;
wire _guard10813 = early_reset_static_par0_go_out;
wire _guard10814 = fsm0_out == 6'd0;
wire _guard10815 = early_reset_static_seq_go_out;
wire _guard10816 = _guard10814 & _guard10815;
wire _guard10817 = early_reset_static_par0_go_out;
wire _guard10818 = _guard10816 | _guard10817;
wire _guard10819 = early_reset_static_par0_go_out;
wire _guard10820 = fsm0_out == 6'd0;
wire _guard10821 = early_reset_static_seq_go_out;
wire _guard10822 = _guard10820 & _guard10821;
wire _guard10823 = early_reset_static_par0_go_out;
wire _guard10824 = early_reset_static_par0_go_out;
wire _guard10825 = ~_guard0;
wire _guard10826 = early_reset_static_par0_go_out;
wire _guard10827 = _guard10825 & _guard10826;
wire _guard10828 = early_reset_static_par0_go_out;
wire _guard10829 = early_reset_static_par0_go_out;
wire _guard10830 = early_reset_static_par0_go_out;
wire _guard10831 = early_reset_static_par0_go_out;
wire _guard10832 = ~_guard0;
wire _guard10833 = early_reset_static_par0_go_out;
wire _guard10834 = _guard10832 & _guard10833;
wire _guard10835 = early_reset_static_par0_go_out;
wire _guard10836 = early_reset_static_par0_go_out;
wire _guard10837 = early_reset_static_par0_go_out;
wire _guard10838 = early_reset_static_par0_go_out;
wire _guard10839 = early_reset_static_par0_go_out;
wire _guard10840 = early_reset_static_par0_go_out;
wire _guard10841 = early_reset_static_par0_go_out;
wire _guard10842 = ~_guard0;
wire _guard10843 = early_reset_static_par0_go_out;
wire _guard10844 = _guard10842 & _guard10843;
wire _guard10845 = early_reset_static_par0_go_out;
wire _guard10846 = ~_guard0;
wire _guard10847 = early_reset_static_par0_go_out;
wire _guard10848 = _guard10846 & _guard10847;
wire _guard10849 = early_reset_static_par0_go_out;
wire _guard10850 = early_reset_static_par0_go_out;
wire _guard10851 = early_reset_static_par0_go_out;
wire _guard10852 = early_reset_static_par0_go_out;
wire _guard10853 = early_reset_static_par0_go_out;
wire _guard10854 = early_reset_static_par0_go_out;
wire _guard10855 = early_reset_static_par0_go_out;
wire _guard10856 = ~_guard0;
wire _guard10857 = early_reset_static_par0_go_out;
wire _guard10858 = _guard10856 & _guard10857;
wire _guard10859 = ~_guard0;
wire _guard10860 = early_reset_static_par0_go_out;
wire _guard10861 = _guard10859 & _guard10860;
wire _guard10862 = early_reset_static_par0_go_out;
wire _guard10863 = ~_guard0;
wire _guard10864 = early_reset_static_par0_go_out;
wire _guard10865 = _guard10863 & _guard10864;
wire _guard10866 = early_reset_static_par0_go_out;
wire _guard10867 = early_reset_static_par0_go_out;
wire _guard10868 = ~_guard0;
wire _guard10869 = early_reset_static_par0_go_out;
wire _guard10870 = _guard10868 & _guard10869;
wire _guard10871 = early_reset_static_par0_go_out;
wire _guard10872 = early_reset_static_par0_go_out;
wire _guard10873 = early_reset_static_par0_go_out;
wire _guard10874 = early_reset_static_par0_go_out;
wire _guard10875 = early_reset_static_par0_go_out;
wire _guard10876 = early_reset_static_par0_go_out;
wire _guard10877 = early_reset_static_par0_go_out;
wire _guard10878 = early_reset_static_par0_go_out;
wire _guard10879 = early_reset_static_par0_go_out;
wire _guard10880 = early_reset_static_par0_go_out;
wire _guard10881 = ~_guard0;
wire _guard10882 = early_reset_static_par0_go_out;
wire _guard10883 = _guard10881 & _guard10882;
wire _guard10884 = early_reset_static_par0_go_out;
wire _guard10885 = early_reset_static_par0_go_out;
wire _guard10886 = ~_guard0;
wire _guard10887 = early_reset_static_par0_go_out;
wire _guard10888 = _guard10886 & _guard10887;
wire _guard10889 = early_reset_static_par0_go_out;
wire _guard10890 = early_reset_static_par0_go_out;
wire _guard10891 = early_reset_static_par0_go_out;
wire _guard10892 = ~_guard0;
wire _guard10893 = early_reset_static_par0_go_out;
wire _guard10894 = _guard10892 & _guard10893;
wire _guard10895 = early_reset_static_par0_go_out;
wire _guard10896 = early_reset_static_par0_go_out;
wire _guard10897 = early_reset_static_par0_go_out;
wire _guard10898 = early_reset_static_par0_go_out;
wire _guard10899 = early_reset_static_par0_go_out;
wire _guard10900 = early_reset_static_par0_go_out;
wire _guard10901 = early_reset_static_par0_go_out;
wire _guard10902 = ~_guard0;
wire _guard10903 = early_reset_static_par0_go_out;
wire _guard10904 = _guard10902 & _guard10903;
wire _guard10905 = early_reset_static_par0_go_out;
wire _guard10906 = ~_guard0;
wire _guard10907 = early_reset_static_par0_go_out;
wire _guard10908 = _guard10906 & _guard10907;
wire _guard10909 = early_reset_static_par0_go_out;
wire _guard10910 = ~_guard0;
wire _guard10911 = early_reset_static_par0_go_out;
wire _guard10912 = _guard10910 & _guard10911;
wire _guard10913 = ~_guard0;
wire _guard10914 = early_reset_static_par0_go_out;
wire _guard10915 = _guard10913 & _guard10914;
wire _guard10916 = early_reset_static_par0_go_out;
wire _guard10917 = early_reset_static_par0_go_out;
wire _guard10918 = early_reset_static_par0_go_out;
wire _guard10919 = early_reset_static_par0_go_out;
wire _guard10920 = ~_guard0;
wire _guard10921 = early_reset_static_par0_go_out;
wire _guard10922 = _guard10920 & _guard10921;
wire _guard10923 = early_reset_static_par0_go_out;
wire _guard10924 = ~_guard0;
wire _guard10925 = early_reset_static_par0_go_out;
wire _guard10926 = _guard10924 & _guard10925;
wire _guard10927 = early_reset_static_par0_go_out;
wire _guard10928 = early_reset_static_par0_go_out;
wire _guard10929 = early_reset_static_par0_go_out;
wire _guard10930 = early_reset_static_par0_go_out;
wire _guard10931 = ~_guard0;
wire _guard10932 = early_reset_static_par0_go_out;
wire _guard10933 = _guard10931 & _guard10932;
wire _guard10934 = early_reset_static_par0_go_out;
wire _guard10935 = early_reset_static_par0_go_out;
wire _guard10936 = early_reset_static_par0_go_out;
wire _guard10937 = ~_guard0;
wire _guard10938 = early_reset_static_par0_go_out;
wire _guard10939 = _guard10937 & _guard10938;
wire _guard10940 = early_reset_static_par0_go_out;
wire _guard10941 = early_reset_static_par0_go_out;
wire _guard10942 = early_reset_static_par0_go_out;
wire _guard10943 = early_reset_static_par0_go_out;
wire _guard10944 = ~_guard0;
wire _guard10945 = early_reset_static_par0_go_out;
wire _guard10946 = _guard10944 & _guard10945;
wire _guard10947 = ~_guard0;
wire _guard10948 = early_reset_static_par0_go_out;
wire _guard10949 = _guard10947 & _guard10948;
wire _guard10950 = early_reset_static_par0_go_out;
wire _guard10951 = early_reset_static_par0_go_out;
wire _guard10952 = early_reset_static_par0_go_out;
wire _guard10953 = early_reset_static_par0_go_out;
wire _guard10954 = ~_guard0;
wire _guard10955 = early_reset_static_par0_go_out;
wire _guard10956 = _guard10954 & _guard10955;
wire _guard10957 = early_reset_static_par0_go_out;
wire _guard10958 = ~_guard0;
wire _guard10959 = early_reset_static_par0_go_out;
wire _guard10960 = _guard10958 & _guard10959;
wire _guard10961 = early_reset_static_par0_go_out;
wire _guard10962 = early_reset_static_par0_go_out;
wire _guard10963 = early_reset_static_par0_go_out;
wire _guard10964 = early_reset_static_par0_go_out;
wire _guard10965 = ~_guard0;
wire _guard10966 = early_reset_static_par0_go_out;
wire _guard10967 = _guard10965 & _guard10966;
wire _guard10968 = early_reset_static_par0_go_out;
wire _guard10969 = early_reset_static_par0_go_out;
wire _guard10970 = early_reset_static_par0_go_out;
wire _guard10971 = early_reset_static_par0_go_out;
wire _guard10972 = early_reset_static_par0_go_out;
wire _guard10973 = early_reset_static_par0_go_out;
wire _guard10974 = early_reset_static_par0_go_out;
wire _guard10975 = early_reset_static_par0_go_out;
wire _guard10976 = early_reset_static_par0_go_out;
wire _guard10977 = ~_guard0;
wire _guard10978 = early_reset_static_par0_go_out;
wire _guard10979 = _guard10977 & _guard10978;
wire _guard10980 = early_reset_static_par0_go_out;
wire _guard10981 = early_reset_static_par0_go_out;
wire _guard10982 = ~_guard0;
wire _guard10983 = early_reset_static_par0_go_out;
wire _guard10984 = _guard10982 & _guard10983;
wire _guard10985 = early_reset_static_par0_go_out;
wire _guard10986 = early_reset_static_par0_go_out;
wire _guard10987 = ~_guard0;
wire _guard10988 = early_reset_static_par0_go_out;
wire _guard10989 = _guard10987 & _guard10988;
wire _guard10990 = early_reset_static_par0_go_out;
wire _guard10991 = early_reset_static_par0_go_out;
wire _guard10992 = early_reset_static_par0_go_out;
wire _guard10993 = early_reset_static_par0_go_out;
wire _guard10994 = early_reset_static_par0_go_out;
wire _guard10995 = early_reset_static_par0_go_out;
wire _guard10996 = early_reset_static_par0_go_out;
wire _guard10997 = early_reset_static_par0_go_out;
wire _guard10998 = early_reset_static_par0_go_out;
wire _guard10999 = early_reset_static_par0_go_out;
wire _guard11000 = ~_guard0;
wire _guard11001 = early_reset_static_par0_go_out;
wire _guard11002 = _guard11000 & _guard11001;
wire _guard11003 = early_reset_static_par0_go_out;
wire _guard11004 = early_reset_static_par0_go_out;
wire _guard11005 = early_reset_static_par0_go_out;
wire _guard11006 = ~_guard0;
wire _guard11007 = early_reset_static_par0_go_out;
wire _guard11008 = _guard11006 & _guard11007;
wire _guard11009 = early_reset_static_par0_go_out;
wire _guard11010 = early_reset_static_par0_go_out;
wire _guard11011 = early_reset_static_par0_go_out;
wire _guard11012 = early_reset_static_par0_go_out;
wire _guard11013 = early_reset_static_par0_go_out;
wire _guard11014 = early_reset_static_par0_go_out;
wire _guard11015 = early_reset_static_par0_go_out;
wire _guard11016 = ~_guard0;
wire _guard11017 = early_reset_static_par0_go_out;
wire _guard11018 = _guard11016 & _guard11017;
wire _guard11019 = ~_guard0;
wire _guard11020 = early_reset_static_par0_go_out;
wire _guard11021 = _guard11019 & _guard11020;
wire _guard11022 = early_reset_static_par0_go_out;
wire _guard11023 = early_reset_static_par0_go_out;
wire _guard11024 = early_reset_static_par0_go_out;
wire _guard11025 = early_reset_static_par0_go_out;
wire _guard11026 = early_reset_static_par0_go_out;
wire _guard11027 = ~_guard0;
wire _guard11028 = early_reset_static_par0_go_out;
wire _guard11029 = _guard11027 & _guard11028;
wire _guard11030 = early_reset_static_par0_go_out;
wire _guard11031 = early_reset_static_par0_go_out;
wire _guard11032 = ~_guard0;
wire _guard11033 = early_reset_static_par0_go_out;
wire _guard11034 = _guard11032 & _guard11033;
wire _guard11035 = early_reset_static_par0_go_out;
wire _guard11036 = early_reset_static_par0_go_out;
wire _guard11037 = early_reset_static_par0_go_out;
wire _guard11038 = ~_guard0;
wire _guard11039 = early_reset_static_par0_go_out;
wire _guard11040 = _guard11038 & _guard11039;
wire _guard11041 = ~_guard0;
wire _guard11042 = early_reset_static_par0_go_out;
wire _guard11043 = _guard11041 & _guard11042;
wire _guard11044 = early_reset_static_par0_go_out;
wire _guard11045 = early_reset_static_par0_go_out;
wire _guard11046 = ~_guard0;
wire _guard11047 = early_reset_static_par0_go_out;
wire _guard11048 = _guard11046 & _guard11047;
wire _guard11049 = early_reset_static_par0_go_out;
wire _guard11050 = ~_guard0;
wire _guard11051 = early_reset_static_par0_go_out;
wire _guard11052 = _guard11050 & _guard11051;
wire _guard11053 = early_reset_static_par0_go_out;
wire _guard11054 = ~_guard0;
wire _guard11055 = early_reset_static_par0_go_out;
wire _guard11056 = _guard11054 & _guard11055;
wire _guard11057 = early_reset_static_par0_go_out;
wire _guard11058 = early_reset_static_par0_go_out;
wire _guard11059 = ~_guard0;
wire _guard11060 = early_reset_static_par0_go_out;
wire _guard11061 = _guard11059 & _guard11060;
wire _guard11062 = early_reset_static_par0_go_out;
wire _guard11063 = early_reset_static_par0_go_out;
wire _guard11064 = early_reset_static_par0_go_out;
wire _guard11065 = early_reset_static_par0_go_out;
wire _guard11066 = early_reset_static_par0_go_out;
wire _guard11067 = early_reset_static_par0_go_out;
wire _guard11068 = early_reset_static_par0_go_out;
wire _guard11069 = early_reset_static_par0_go_out;
wire _guard11070 = ~_guard0;
wire _guard11071 = early_reset_static_par0_go_out;
wire _guard11072 = _guard11070 & _guard11071;
wire _guard11073 = early_reset_static_par0_go_out;
wire _guard11074 = early_reset_static_par0_go_out;
wire _guard11075 = early_reset_static_par0_go_out;
wire _guard11076 = early_reset_static_par0_go_out;
wire _guard11077 = early_reset_static_par0_go_out;
wire _guard11078 = early_reset_static_par0_go_out;
wire _guard11079 = early_reset_static_par0_go_out;
wire _guard11080 = ~_guard0;
wire _guard11081 = early_reset_static_par0_go_out;
wire _guard11082 = _guard11080 & _guard11081;
wire _guard11083 = early_reset_static_par0_go_out;
wire _guard11084 = early_reset_static_par0_go_out;
wire _guard11085 = early_reset_static_par0_go_out;
wire _guard11086 = early_reset_static_par0_go_out;
wire _guard11087 = early_reset_static_par0_go_out;
wire _guard11088 = early_reset_static_par0_go_out;
wire _guard11089 = ~_guard0;
wire _guard11090 = early_reset_static_par0_go_out;
wire _guard11091 = _guard11089 & _guard11090;
wire _guard11092 = early_reset_static_par0_go_out;
wire _guard11093 = early_reset_static_par0_go_out;
wire _guard11094 = early_reset_static_par0_go_out;
wire _guard11095 = ~_guard0;
wire _guard11096 = early_reset_static_par0_go_out;
wire _guard11097 = _guard11095 & _guard11096;
wire _guard11098 = early_reset_static_par0_go_out;
wire _guard11099 = early_reset_static_par0_go_out;
wire _guard11100 = early_reset_static_par0_go_out;
wire _guard11101 = ~_guard0;
wire _guard11102 = early_reset_static_par0_go_out;
wire _guard11103 = _guard11101 & _guard11102;
wire _guard11104 = early_reset_static_par0_go_out;
wire _guard11105 = early_reset_static_par0_go_out;
wire _guard11106 = early_reset_static_par0_go_out;
wire _guard11107 = early_reset_static_par0_go_out;
wire _guard11108 = early_reset_static_par0_go_out;
wire _guard11109 = early_reset_static_par0_go_out;
wire _guard11110 = early_reset_static_par0_go_out;
wire _guard11111 = early_reset_static_par0_go_out;
wire _guard11112 = early_reset_static_par0_go_out;
wire _guard11113 = early_reset_static_par0_go_out;
wire _guard11114 = early_reset_static_par0_go_out;
wire _guard11115 = early_reset_static_par0_go_out;
wire _guard11116 = early_reset_static_par0_go_out;
wire _guard11117 = early_reset_static_par0_go_out;
wire _guard11118 = ~_guard0;
wire _guard11119 = early_reset_static_par0_go_out;
wire _guard11120 = _guard11118 & _guard11119;
wire _guard11121 = early_reset_static_par0_go_out;
wire _guard11122 = ~_guard0;
wire _guard11123 = early_reset_static_par0_go_out;
wire _guard11124 = _guard11122 & _guard11123;
wire _guard11125 = early_reset_static_par0_go_out;
wire _guard11126 = early_reset_static_par0_go_out;
wire _guard11127 = ~_guard0;
wire _guard11128 = early_reset_static_par0_go_out;
wire _guard11129 = _guard11127 & _guard11128;
wire _guard11130 = early_reset_static_par0_go_out;
wire _guard11131 = early_reset_static_par0_go_out;
wire _guard11132 = ~_guard0;
wire _guard11133 = early_reset_static_par0_go_out;
wire _guard11134 = _guard11132 & _guard11133;
wire _guard11135 = early_reset_static_par0_go_out;
wire _guard11136 = early_reset_static_par0_go_out;
wire _guard11137 = early_reset_static_par0_go_out;
wire _guard11138 = early_reset_static_par0_go_out;
wire _guard11139 = early_reset_static_par0_go_out;
wire _guard11140 = early_reset_static_par0_go_out;
wire _guard11141 = early_reset_static_par0_go_out;
wire _guard11142 = early_reset_static_par0_go_out;
wire _guard11143 = early_reset_static_par0_go_out;
wire _guard11144 = early_reset_static_par0_go_out;
wire _guard11145 = early_reset_static_par0_go_out;
wire _guard11146 = early_reset_static_par0_go_out;
wire _guard11147 = early_reset_static_par0_go_out;
wire _guard11148 = ~_guard0;
wire _guard11149 = early_reset_static_par0_go_out;
wire _guard11150 = _guard11148 & _guard11149;
wire _guard11151 = ~_guard0;
wire _guard11152 = early_reset_static_par0_go_out;
wire _guard11153 = _guard11151 & _guard11152;
wire _guard11154 = early_reset_static_par0_go_out;
wire _guard11155 = early_reset_static_par0_go_out;
wire _guard11156 = early_reset_static_par0_go_out;
wire _guard11157 = early_reset_static_par0_go_out;
wire _guard11158 = early_reset_static_par0_go_out;
wire _guard11159 = ~_guard0;
wire _guard11160 = early_reset_static_par0_go_out;
wire _guard11161 = _guard11159 & _guard11160;
wire _guard11162 = early_reset_static_par0_go_out;
wire _guard11163 = early_reset_static_par0_go_out;
wire _guard11164 = early_reset_static_par0_go_out;
wire _guard11165 = early_reset_static_par0_go_out;
wire _guard11166 = early_reset_static_par0_go_out;
wire _guard11167 = early_reset_static_par0_go_out;
wire _guard11168 = early_reset_static_par0_go_out;
wire _guard11169 = early_reset_static_par0_go_out;
wire _guard11170 = ~_guard0;
wire _guard11171 = early_reset_static_par0_go_out;
wire _guard11172 = _guard11170 & _guard11171;
wire _guard11173 = early_reset_static_par0_go_out;
wire _guard11174 = early_reset_static_par0_go_out;
wire _guard11175 = ~_guard0;
wire _guard11176 = early_reset_static_par0_go_out;
wire _guard11177 = _guard11175 & _guard11176;
wire _guard11178 = early_reset_static_par0_go_out;
wire _guard11179 = early_reset_static_par0_go_out;
wire _guard11180 = ~_guard0;
wire _guard11181 = early_reset_static_par0_go_out;
wire _guard11182 = _guard11180 & _guard11181;
wire _guard11183 = early_reset_static_par0_go_out;
wire _guard11184 = ~_guard0;
wire _guard11185 = early_reset_static_par0_go_out;
wire _guard11186 = _guard11184 & _guard11185;
wire _guard11187 = cond_wire12_out;
wire _guard11188 = early_reset_static_par0_go_out;
wire _guard11189 = _guard11187 & _guard11188;
wire _guard11190 = cond_wire10_out;
wire _guard11191 = early_reset_static_par0_go_out;
wire _guard11192 = _guard11190 & _guard11191;
wire _guard11193 = fsm_out == 1'd0;
wire _guard11194 = cond_wire10_out;
wire _guard11195 = _guard11193 & _guard11194;
wire _guard11196 = fsm_out == 1'd0;
wire _guard11197 = _guard11195 & _guard11196;
wire _guard11198 = fsm_out == 1'd0;
wire _guard11199 = cond_wire12_out;
wire _guard11200 = _guard11198 & _guard11199;
wire _guard11201 = fsm_out == 1'd0;
wire _guard11202 = _guard11200 & _guard11201;
wire _guard11203 = _guard11197 | _guard11202;
wire _guard11204 = early_reset_static_par0_go_out;
wire _guard11205 = _guard11203 & _guard11204;
wire _guard11206 = fsm_out == 1'd0;
wire _guard11207 = cond_wire10_out;
wire _guard11208 = _guard11206 & _guard11207;
wire _guard11209 = fsm_out == 1'd0;
wire _guard11210 = _guard11208 & _guard11209;
wire _guard11211 = fsm_out == 1'd0;
wire _guard11212 = cond_wire12_out;
wire _guard11213 = _guard11211 & _guard11212;
wire _guard11214 = fsm_out == 1'd0;
wire _guard11215 = _guard11213 & _guard11214;
wire _guard11216 = _guard11210 | _guard11215;
wire _guard11217 = early_reset_static_par0_go_out;
wire _guard11218 = _guard11216 & _guard11217;
wire _guard11219 = fsm_out == 1'd0;
wire _guard11220 = cond_wire10_out;
wire _guard11221 = _guard11219 & _guard11220;
wire _guard11222 = fsm_out == 1'd0;
wire _guard11223 = _guard11221 & _guard11222;
wire _guard11224 = fsm_out == 1'd0;
wire _guard11225 = cond_wire12_out;
wire _guard11226 = _guard11224 & _guard11225;
wire _guard11227 = fsm_out == 1'd0;
wire _guard11228 = _guard11226 & _guard11227;
wire _guard11229 = _guard11223 | _guard11228;
wire _guard11230 = early_reset_static_par0_go_out;
wire _guard11231 = _guard11229 & _guard11230;
wire _guard11232 = cond_wire62_out;
wire _guard11233 = early_reset_static_par0_go_out;
wire _guard11234 = _guard11232 & _guard11233;
wire _guard11235 = cond_wire60_out;
wire _guard11236 = early_reset_static_par0_go_out;
wire _guard11237 = _guard11235 & _guard11236;
wire _guard11238 = fsm_out == 1'd0;
wire _guard11239 = cond_wire60_out;
wire _guard11240 = _guard11238 & _guard11239;
wire _guard11241 = fsm_out == 1'd0;
wire _guard11242 = _guard11240 & _guard11241;
wire _guard11243 = fsm_out == 1'd0;
wire _guard11244 = cond_wire62_out;
wire _guard11245 = _guard11243 & _guard11244;
wire _guard11246 = fsm_out == 1'd0;
wire _guard11247 = _guard11245 & _guard11246;
wire _guard11248 = _guard11242 | _guard11247;
wire _guard11249 = early_reset_static_par0_go_out;
wire _guard11250 = _guard11248 & _guard11249;
wire _guard11251 = fsm_out == 1'd0;
wire _guard11252 = cond_wire60_out;
wire _guard11253 = _guard11251 & _guard11252;
wire _guard11254 = fsm_out == 1'd0;
wire _guard11255 = _guard11253 & _guard11254;
wire _guard11256 = fsm_out == 1'd0;
wire _guard11257 = cond_wire62_out;
wire _guard11258 = _guard11256 & _guard11257;
wire _guard11259 = fsm_out == 1'd0;
wire _guard11260 = _guard11258 & _guard11259;
wire _guard11261 = _guard11255 | _guard11260;
wire _guard11262 = early_reset_static_par0_go_out;
wire _guard11263 = _guard11261 & _guard11262;
wire _guard11264 = fsm_out == 1'd0;
wire _guard11265 = cond_wire60_out;
wire _guard11266 = _guard11264 & _guard11265;
wire _guard11267 = fsm_out == 1'd0;
wire _guard11268 = _guard11266 & _guard11267;
wire _guard11269 = fsm_out == 1'd0;
wire _guard11270 = cond_wire62_out;
wire _guard11271 = _guard11269 & _guard11270;
wire _guard11272 = fsm_out == 1'd0;
wire _guard11273 = _guard11271 & _guard11272;
wire _guard11274 = _guard11268 | _guard11273;
wire _guard11275 = early_reset_static_par0_go_out;
wire _guard11276 = _guard11274 & _guard11275;
wire _guard11277 = cond_wire77_out;
wire _guard11278 = early_reset_static_par0_go_out;
wire _guard11279 = _guard11277 & _guard11278;
wire _guard11280 = cond_wire75_out;
wire _guard11281 = early_reset_static_par0_go_out;
wire _guard11282 = _guard11280 & _guard11281;
wire _guard11283 = fsm_out == 1'd0;
wire _guard11284 = cond_wire75_out;
wire _guard11285 = _guard11283 & _guard11284;
wire _guard11286 = fsm_out == 1'd0;
wire _guard11287 = _guard11285 & _guard11286;
wire _guard11288 = fsm_out == 1'd0;
wire _guard11289 = cond_wire77_out;
wire _guard11290 = _guard11288 & _guard11289;
wire _guard11291 = fsm_out == 1'd0;
wire _guard11292 = _guard11290 & _guard11291;
wire _guard11293 = _guard11287 | _guard11292;
wire _guard11294 = early_reset_static_par0_go_out;
wire _guard11295 = _guard11293 & _guard11294;
wire _guard11296 = fsm_out == 1'd0;
wire _guard11297 = cond_wire75_out;
wire _guard11298 = _guard11296 & _guard11297;
wire _guard11299 = fsm_out == 1'd0;
wire _guard11300 = _guard11298 & _guard11299;
wire _guard11301 = fsm_out == 1'd0;
wire _guard11302 = cond_wire77_out;
wire _guard11303 = _guard11301 & _guard11302;
wire _guard11304 = fsm_out == 1'd0;
wire _guard11305 = _guard11303 & _guard11304;
wire _guard11306 = _guard11300 | _guard11305;
wire _guard11307 = early_reset_static_par0_go_out;
wire _guard11308 = _guard11306 & _guard11307;
wire _guard11309 = fsm_out == 1'd0;
wire _guard11310 = cond_wire75_out;
wire _guard11311 = _guard11309 & _guard11310;
wire _guard11312 = fsm_out == 1'd0;
wire _guard11313 = _guard11311 & _guard11312;
wire _guard11314 = fsm_out == 1'd0;
wire _guard11315 = cond_wire77_out;
wire _guard11316 = _guard11314 & _guard11315;
wire _guard11317 = fsm_out == 1'd0;
wire _guard11318 = _guard11316 & _guard11317;
wire _guard11319 = _guard11313 | _guard11318;
wire _guard11320 = early_reset_static_par0_go_out;
wire _guard11321 = _guard11319 & _guard11320;
wire _guard11322 = cond_wire106_out;
wire _guard11323 = early_reset_static_par0_go_out;
wire _guard11324 = _guard11322 & _guard11323;
wire _guard11325 = cond_wire104_out;
wire _guard11326 = early_reset_static_par0_go_out;
wire _guard11327 = _guard11325 & _guard11326;
wire _guard11328 = fsm_out == 1'd0;
wire _guard11329 = cond_wire104_out;
wire _guard11330 = _guard11328 & _guard11329;
wire _guard11331 = fsm_out == 1'd0;
wire _guard11332 = _guard11330 & _guard11331;
wire _guard11333 = fsm_out == 1'd0;
wire _guard11334 = cond_wire106_out;
wire _guard11335 = _guard11333 & _guard11334;
wire _guard11336 = fsm_out == 1'd0;
wire _guard11337 = _guard11335 & _guard11336;
wire _guard11338 = _guard11332 | _guard11337;
wire _guard11339 = early_reset_static_par0_go_out;
wire _guard11340 = _guard11338 & _guard11339;
wire _guard11341 = fsm_out == 1'd0;
wire _guard11342 = cond_wire104_out;
wire _guard11343 = _guard11341 & _guard11342;
wire _guard11344 = fsm_out == 1'd0;
wire _guard11345 = _guard11343 & _guard11344;
wire _guard11346 = fsm_out == 1'd0;
wire _guard11347 = cond_wire106_out;
wire _guard11348 = _guard11346 & _guard11347;
wire _guard11349 = fsm_out == 1'd0;
wire _guard11350 = _guard11348 & _guard11349;
wire _guard11351 = _guard11345 | _guard11350;
wire _guard11352 = early_reset_static_par0_go_out;
wire _guard11353 = _guard11351 & _guard11352;
wire _guard11354 = fsm_out == 1'd0;
wire _guard11355 = cond_wire104_out;
wire _guard11356 = _guard11354 & _guard11355;
wire _guard11357 = fsm_out == 1'd0;
wire _guard11358 = _guard11356 & _guard11357;
wire _guard11359 = fsm_out == 1'd0;
wire _guard11360 = cond_wire106_out;
wire _guard11361 = _guard11359 & _guard11360;
wire _guard11362 = fsm_out == 1'd0;
wire _guard11363 = _guard11361 & _guard11362;
wire _guard11364 = _guard11358 | _guard11363;
wire _guard11365 = early_reset_static_par0_go_out;
wire _guard11366 = _guard11364 & _guard11365;
wire _guard11367 = cond_wire227_out;
wire _guard11368 = early_reset_static_par0_go_out;
wire _guard11369 = _guard11367 & _guard11368;
wire _guard11370 = cond_wire227_out;
wire _guard11371 = early_reset_static_par0_go_out;
wire _guard11372 = _guard11370 & _guard11371;
wire _guard11373 = cond_wire264_out;
wire _guard11374 = early_reset_static_par0_go_out;
wire _guard11375 = _guard11373 & _guard11374;
wire _guard11376 = cond_wire262_out;
wire _guard11377 = early_reset_static_par0_go_out;
wire _guard11378 = _guard11376 & _guard11377;
wire _guard11379 = fsm_out == 1'd0;
wire _guard11380 = cond_wire262_out;
wire _guard11381 = _guard11379 & _guard11380;
wire _guard11382 = fsm_out == 1'd0;
wire _guard11383 = _guard11381 & _guard11382;
wire _guard11384 = fsm_out == 1'd0;
wire _guard11385 = cond_wire264_out;
wire _guard11386 = _guard11384 & _guard11385;
wire _guard11387 = fsm_out == 1'd0;
wire _guard11388 = _guard11386 & _guard11387;
wire _guard11389 = _guard11383 | _guard11388;
wire _guard11390 = early_reset_static_par0_go_out;
wire _guard11391 = _guard11389 & _guard11390;
wire _guard11392 = fsm_out == 1'd0;
wire _guard11393 = cond_wire262_out;
wire _guard11394 = _guard11392 & _guard11393;
wire _guard11395 = fsm_out == 1'd0;
wire _guard11396 = _guard11394 & _guard11395;
wire _guard11397 = fsm_out == 1'd0;
wire _guard11398 = cond_wire264_out;
wire _guard11399 = _guard11397 & _guard11398;
wire _guard11400 = fsm_out == 1'd0;
wire _guard11401 = _guard11399 & _guard11400;
wire _guard11402 = _guard11396 | _guard11401;
wire _guard11403 = early_reset_static_par0_go_out;
wire _guard11404 = _guard11402 & _guard11403;
wire _guard11405 = fsm_out == 1'd0;
wire _guard11406 = cond_wire262_out;
wire _guard11407 = _guard11405 & _guard11406;
wire _guard11408 = fsm_out == 1'd0;
wire _guard11409 = _guard11407 & _guard11408;
wire _guard11410 = fsm_out == 1'd0;
wire _guard11411 = cond_wire264_out;
wire _guard11412 = _guard11410 & _guard11411;
wire _guard11413 = fsm_out == 1'd0;
wire _guard11414 = _guard11412 & _guard11413;
wire _guard11415 = _guard11409 | _guard11414;
wire _guard11416 = early_reset_static_par0_go_out;
wire _guard11417 = _guard11415 & _guard11416;
wire _guard11418 = cond_wire268_out;
wire _guard11419 = early_reset_static_par0_go_out;
wire _guard11420 = _guard11418 & _guard11419;
wire _guard11421 = cond_wire266_out;
wire _guard11422 = early_reset_static_par0_go_out;
wire _guard11423 = _guard11421 & _guard11422;
wire _guard11424 = fsm_out == 1'd0;
wire _guard11425 = cond_wire266_out;
wire _guard11426 = _guard11424 & _guard11425;
wire _guard11427 = fsm_out == 1'd0;
wire _guard11428 = _guard11426 & _guard11427;
wire _guard11429 = fsm_out == 1'd0;
wire _guard11430 = cond_wire268_out;
wire _guard11431 = _guard11429 & _guard11430;
wire _guard11432 = fsm_out == 1'd0;
wire _guard11433 = _guard11431 & _guard11432;
wire _guard11434 = _guard11428 | _guard11433;
wire _guard11435 = early_reset_static_par0_go_out;
wire _guard11436 = _guard11434 & _guard11435;
wire _guard11437 = fsm_out == 1'd0;
wire _guard11438 = cond_wire266_out;
wire _guard11439 = _guard11437 & _guard11438;
wire _guard11440 = fsm_out == 1'd0;
wire _guard11441 = _guard11439 & _guard11440;
wire _guard11442 = fsm_out == 1'd0;
wire _guard11443 = cond_wire268_out;
wire _guard11444 = _guard11442 & _guard11443;
wire _guard11445 = fsm_out == 1'd0;
wire _guard11446 = _guard11444 & _guard11445;
wire _guard11447 = _guard11441 | _guard11446;
wire _guard11448 = early_reset_static_par0_go_out;
wire _guard11449 = _guard11447 & _guard11448;
wire _guard11450 = fsm_out == 1'd0;
wire _guard11451 = cond_wire266_out;
wire _guard11452 = _guard11450 & _guard11451;
wire _guard11453 = fsm_out == 1'd0;
wire _guard11454 = _guard11452 & _guard11453;
wire _guard11455 = fsm_out == 1'd0;
wire _guard11456 = cond_wire268_out;
wire _guard11457 = _guard11455 & _guard11456;
wire _guard11458 = fsm_out == 1'd0;
wire _guard11459 = _guard11457 & _guard11458;
wire _guard11460 = _guard11454 | _guard11459;
wire _guard11461 = early_reset_static_par0_go_out;
wire _guard11462 = _guard11460 & _guard11461;
wire _guard11463 = cond_wire304_out;
wire _guard11464 = early_reset_static_par0_go_out;
wire _guard11465 = _guard11463 & _guard11464;
wire _guard11466 = cond_wire304_out;
wire _guard11467 = early_reset_static_par0_go_out;
wire _guard11468 = _guard11466 & _guard11467;
wire _guard11469 = cond_wire325_out;
wire _guard11470 = early_reset_static_par0_go_out;
wire _guard11471 = _guard11469 & _guard11470;
wire _guard11472 = cond_wire323_out;
wire _guard11473 = early_reset_static_par0_go_out;
wire _guard11474 = _guard11472 & _guard11473;
wire _guard11475 = fsm_out == 1'd0;
wire _guard11476 = cond_wire323_out;
wire _guard11477 = _guard11475 & _guard11476;
wire _guard11478 = fsm_out == 1'd0;
wire _guard11479 = _guard11477 & _guard11478;
wire _guard11480 = fsm_out == 1'd0;
wire _guard11481 = cond_wire325_out;
wire _guard11482 = _guard11480 & _guard11481;
wire _guard11483 = fsm_out == 1'd0;
wire _guard11484 = _guard11482 & _guard11483;
wire _guard11485 = _guard11479 | _guard11484;
wire _guard11486 = early_reset_static_par0_go_out;
wire _guard11487 = _guard11485 & _guard11486;
wire _guard11488 = fsm_out == 1'd0;
wire _guard11489 = cond_wire323_out;
wire _guard11490 = _guard11488 & _guard11489;
wire _guard11491 = fsm_out == 1'd0;
wire _guard11492 = _guard11490 & _guard11491;
wire _guard11493 = fsm_out == 1'd0;
wire _guard11494 = cond_wire325_out;
wire _guard11495 = _guard11493 & _guard11494;
wire _guard11496 = fsm_out == 1'd0;
wire _guard11497 = _guard11495 & _guard11496;
wire _guard11498 = _guard11492 | _guard11497;
wire _guard11499 = early_reset_static_par0_go_out;
wire _guard11500 = _guard11498 & _guard11499;
wire _guard11501 = fsm_out == 1'd0;
wire _guard11502 = cond_wire323_out;
wire _guard11503 = _guard11501 & _guard11502;
wire _guard11504 = fsm_out == 1'd0;
wire _guard11505 = _guard11503 & _guard11504;
wire _guard11506 = fsm_out == 1'd0;
wire _guard11507 = cond_wire325_out;
wire _guard11508 = _guard11506 & _guard11507;
wire _guard11509 = fsm_out == 1'd0;
wire _guard11510 = _guard11508 & _guard11509;
wire _guard11511 = _guard11505 | _guard11510;
wire _guard11512 = early_reset_static_par0_go_out;
wire _guard11513 = _guard11511 & _guard11512;
wire _guard11514 = cond_wire296_out;
wire _guard11515 = early_reset_static_par0_go_out;
wire _guard11516 = _guard11514 & _guard11515;
wire _guard11517 = cond_wire296_out;
wire _guard11518 = early_reset_static_par0_go_out;
wire _guard11519 = _guard11517 & _guard11518;
wire _guard11520 = cond_wire378_out;
wire _guard11521 = early_reset_static_par0_go_out;
wire _guard11522 = _guard11520 & _guard11521;
wire _guard11523 = cond_wire376_out;
wire _guard11524 = early_reset_static_par0_go_out;
wire _guard11525 = _guard11523 & _guard11524;
wire _guard11526 = fsm_out == 1'd0;
wire _guard11527 = cond_wire376_out;
wire _guard11528 = _guard11526 & _guard11527;
wire _guard11529 = fsm_out == 1'd0;
wire _guard11530 = _guard11528 & _guard11529;
wire _guard11531 = fsm_out == 1'd0;
wire _guard11532 = cond_wire378_out;
wire _guard11533 = _guard11531 & _guard11532;
wire _guard11534 = fsm_out == 1'd0;
wire _guard11535 = _guard11533 & _guard11534;
wire _guard11536 = _guard11530 | _guard11535;
wire _guard11537 = early_reset_static_par0_go_out;
wire _guard11538 = _guard11536 & _guard11537;
wire _guard11539 = fsm_out == 1'd0;
wire _guard11540 = cond_wire376_out;
wire _guard11541 = _guard11539 & _guard11540;
wire _guard11542 = fsm_out == 1'd0;
wire _guard11543 = _guard11541 & _guard11542;
wire _guard11544 = fsm_out == 1'd0;
wire _guard11545 = cond_wire378_out;
wire _guard11546 = _guard11544 & _guard11545;
wire _guard11547 = fsm_out == 1'd0;
wire _guard11548 = _guard11546 & _guard11547;
wire _guard11549 = _guard11543 | _guard11548;
wire _guard11550 = early_reset_static_par0_go_out;
wire _guard11551 = _guard11549 & _guard11550;
wire _guard11552 = fsm_out == 1'd0;
wire _guard11553 = cond_wire376_out;
wire _guard11554 = _guard11552 & _guard11553;
wire _guard11555 = fsm_out == 1'd0;
wire _guard11556 = _guard11554 & _guard11555;
wire _guard11557 = fsm_out == 1'd0;
wire _guard11558 = cond_wire378_out;
wire _guard11559 = _guard11557 & _guard11558;
wire _guard11560 = fsm_out == 1'd0;
wire _guard11561 = _guard11559 & _guard11560;
wire _guard11562 = _guard11556 | _guard11561;
wire _guard11563 = early_reset_static_par0_go_out;
wire _guard11564 = _guard11562 & _guard11563;
wire _guard11565 = cond_wire382_out;
wire _guard11566 = early_reset_static_par0_go_out;
wire _guard11567 = _guard11565 & _guard11566;
wire _guard11568 = cond_wire380_out;
wire _guard11569 = early_reset_static_par0_go_out;
wire _guard11570 = _guard11568 & _guard11569;
wire _guard11571 = fsm_out == 1'd0;
wire _guard11572 = cond_wire380_out;
wire _guard11573 = _guard11571 & _guard11572;
wire _guard11574 = fsm_out == 1'd0;
wire _guard11575 = _guard11573 & _guard11574;
wire _guard11576 = fsm_out == 1'd0;
wire _guard11577 = cond_wire382_out;
wire _guard11578 = _guard11576 & _guard11577;
wire _guard11579 = fsm_out == 1'd0;
wire _guard11580 = _guard11578 & _guard11579;
wire _guard11581 = _guard11575 | _guard11580;
wire _guard11582 = early_reset_static_par0_go_out;
wire _guard11583 = _guard11581 & _guard11582;
wire _guard11584 = fsm_out == 1'd0;
wire _guard11585 = cond_wire380_out;
wire _guard11586 = _guard11584 & _guard11585;
wire _guard11587 = fsm_out == 1'd0;
wire _guard11588 = _guard11586 & _guard11587;
wire _guard11589 = fsm_out == 1'd0;
wire _guard11590 = cond_wire382_out;
wire _guard11591 = _guard11589 & _guard11590;
wire _guard11592 = fsm_out == 1'd0;
wire _guard11593 = _guard11591 & _guard11592;
wire _guard11594 = _guard11588 | _guard11593;
wire _guard11595 = early_reset_static_par0_go_out;
wire _guard11596 = _guard11594 & _guard11595;
wire _guard11597 = fsm_out == 1'd0;
wire _guard11598 = cond_wire380_out;
wire _guard11599 = _guard11597 & _guard11598;
wire _guard11600 = fsm_out == 1'd0;
wire _guard11601 = _guard11599 & _guard11600;
wire _guard11602 = fsm_out == 1'd0;
wire _guard11603 = cond_wire382_out;
wire _guard11604 = _guard11602 & _guard11603;
wire _guard11605 = fsm_out == 1'd0;
wire _guard11606 = _guard11604 & _guard11605;
wire _guard11607 = _guard11601 | _guard11606;
wire _guard11608 = early_reset_static_par0_go_out;
wire _guard11609 = _guard11607 & _guard11608;
wire _guard11610 = cond_wire381_out;
wire _guard11611 = early_reset_static_par0_go_out;
wire _guard11612 = _guard11610 & _guard11611;
wire _guard11613 = cond_wire381_out;
wire _guard11614 = early_reset_static_par0_go_out;
wire _guard11615 = _guard11613 & _guard11614;
wire _guard11616 = cond_wire406_out;
wire _guard11617 = early_reset_static_par0_go_out;
wire _guard11618 = _guard11616 & _guard11617;
wire _guard11619 = cond_wire406_out;
wire _guard11620 = early_reset_static_par0_go_out;
wire _guard11621 = _guard11619 & _guard11620;
wire _guard11622 = cond_wire427_out;
wire _guard11623 = early_reset_static_par0_go_out;
wire _guard11624 = _guard11622 & _guard11623;
wire _guard11625 = cond_wire425_out;
wire _guard11626 = early_reset_static_par0_go_out;
wire _guard11627 = _guard11625 & _guard11626;
wire _guard11628 = fsm_out == 1'd0;
wire _guard11629 = cond_wire425_out;
wire _guard11630 = _guard11628 & _guard11629;
wire _guard11631 = fsm_out == 1'd0;
wire _guard11632 = _guard11630 & _guard11631;
wire _guard11633 = fsm_out == 1'd0;
wire _guard11634 = cond_wire427_out;
wire _guard11635 = _guard11633 & _guard11634;
wire _guard11636 = fsm_out == 1'd0;
wire _guard11637 = _guard11635 & _guard11636;
wire _guard11638 = _guard11632 | _guard11637;
wire _guard11639 = early_reset_static_par0_go_out;
wire _guard11640 = _guard11638 & _guard11639;
wire _guard11641 = fsm_out == 1'd0;
wire _guard11642 = cond_wire425_out;
wire _guard11643 = _guard11641 & _guard11642;
wire _guard11644 = fsm_out == 1'd0;
wire _guard11645 = _guard11643 & _guard11644;
wire _guard11646 = fsm_out == 1'd0;
wire _guard11647 = cond_wire427_out;
wire _guard11648 = _guard11646 & _guard11647;
wire _guard11649 = fsm_out == 1'd0;
wire _guard11650 = _guard11648 & _guard11649;
wire _guard11651 = _guard11645 | _guard11650;
wire _guard11652 = early_reset_static_par0_go_out;
wire _guard11653 = _guard11651 & _guard11652;
wire _guard11654 = fsm_out == 1'd0;
wire _guard11655 = cond_wire425_out;
wire _guard11656 = _guard11654 & _guard11655;
wire _guard11657 = fsm_out == 1'd0;
wire _guard11658 = _guard11656 & _guard11657;
wire _guard11659 = fsm_out == 1'd0;
wire _guard11660 = cond_wire427_out;
wire _guard11661 = _guard11659 & _guard11660;
wire _guard11662 = fsm_out == 1'd0;
wire _guard11663 = _guard11661 & _guard11662;
wire _guard11664 = _guard11658 | _guard11663;
wire _guard11665 = early_reset_static_par0_go_out;
wire _guard11666 = _guard11664 & _guard11665;
wire _guard11667 = cond_wire430_out;
wire _guard11668 = early_reset_static_par0_go_out;
wire _guard11669 = _guard11667 & _guard11668;
wire _guard11670 = cond_wire430_out;
wire _guard11671 = early_reset_static_par0_go_out;
wire _guard11672 = _guard11670 & _guard11671;
wire _guard11673 = cond_wire455_out;
wire _guard11674 = early_reset_static_par0_go_out;
wire _guard11675 = _guard11673 & _guard11674;
wire _guard11676 = cond_wire453_out;
wire _guard11677 = early_reset_static_par0_go_out;
wire _guard11678 = _guard11676 & _guard11677;
wire _guard11679 = fsm_out == 1'd0;
wire _guard11680 = cond_wire453_out;
wire _guard11681 = _guard11679 & _guard11680;
wire _guard11682 = fsm_out == 1'd0;
wire _guard11683 = _guard11681 & _guard11682;
wire _guard11684 = fsm_out == 1'd0;
wire _guard11685 = cond_wire455_out;
wire _guard11686 = _guard11684 & _guard11685;
wire _guard11687 = fsm_out == 1'd0;
wire _guard11688 = _guard11686 & _guard11687;
wire _guard11689 = _guard11683 | _guard11688;
wire _guard11690 = early_reset_static_par0_go_out;
wire _guard11691 = _guard11689 & _guard11690;
wire _guard11692 = fsm_out == 1'd0;
wire _guard11693 = cond_wire453_out;
wire _guard11694 = _guard11692 & _guard11693;
wire _guard11695 = fsm_out == 1'd0;
wire _guard11696 = _guard11694 & _guard11695;
wire _guard11697 = fsm_out == 1'd0;
wire _guard11698 = cond_wire455_out;
wire _guard11699 = _guard11697 & _guard11698;
wire _guard11700 = fsm_out == 1'd0;
wire _guard11701 = _guard11699 & _guard11700;
wire _guard11702 = _guard11696 | _guard11701;
wire _guard11703 = early_reset_static_par0_go_out;
wire _guard11704 = _guard11702 & _guard11703;
wire _guard11705 = fsm_out == 1'd0;
wire _guard11706 = cond_wire453_out;
wire _guard11707 = _guard11705 & _guard11706;
wire _guard11708 = fsm_out == 1'd0;
wire _guard11709 = _guard11707 & _guard11708;
wire _guard11710 = fsm_out == 1'd0;
wire _guard11711 = cond_wire455_out;
wire _guard11712 = _guard11710 & _guard11711;
wire _guard11713 = fsm_out == 1'd0;
wire _guard11714 = _guard11712 & _guard11713;
wire _guard11715 = _guard11709 | _guard11714;
wire _guard11716 = early_reset_static_par0_go_out;
wire _guard11717 = _guard11715 & _guard11716;
wire _guard11718 = cond_wire389_out;
wire _guard11719 = early_reset_static_par0_go_out;
wire _guard11720 = _guard11718 & _guard11719;
wire _guard11721 = cond_wire389_out;
wire _guard11722 = early_reset_static_par0_go_out;
wire _guard11723 = _guard11721 & _guard11722;
wire _guard11724 = cond_wire472_out;
wire _guard11725 = early_reset_static_par0_go_out;
wire _guard11726 = _guard11724 & _guard11725;
wire _guard11727 = cond_wire470_out;
wire _guard11728 = early_reset_static_par0_go_out;
wire _guard11729 = _guard11727 & _guard11728;
wire _guard11730 = fsm_out == 1'd0;
wire _guard11731 = cond_wire470_out;
wire _guard11732 = _guard11730 & _guard11731;
wire _guard11733 = fsm_out == 1'd0;
wire _guard11734 = _guard11732 & _guard11733;
wire _guard11735 = fsm_out == 1'd0;
wire _guard11736 = cond_wire472_out;
wire _guard11737 = _guard11735 & _guard11736;
wire _guard11738 = fsm_out == 1'd0;
wire _guard11739 = _guard11737 & _guard11738;
wire _guard11740 = _guard11734 | _guard11739;
wire _guard11741 = early_reset_static_par0_go_out;
wire _guard11742 = _guard11740 & _guard11741;
wire _guard11743 = fsm_out == 1'd0;
wire _guard11744 = cond_wire470_out;
wire _guard11745 = _guard11743 & _guard11744;
wire _guard11746 = fsm_out == 1'd0;
wire _guard11747 = _guard11745 & _guard11746;
wire _guard11748 = fsm_out == 1'd0;
wire _guard11749 = cond_wire472_out;
wire _guard11750 = _guard11748 & _guard11749;
wire _guard11751 = fsm_out == 1'd0;
wire _guard11752 = _guard11750 & _guard11751;
wire _guard11753 = _guard11747 | _guard11752;
wire _guard11754 = early_reset_static_par0_go_out;
wire _guard11755 = _guard11753 & _guard11754;
wire _guard11756 = fsm_out == 1'd0;
wire _guard11757 = cond_wire470_out;
wire _guard11758 = _guard11756 & _guard11757;
wire _guard11759 = fsm_out == 1'd0;
wire _guard11760 = _guard11758 & _guard11759;
wire _guard11761 = fsm_out == 1'd0;
wire _guard11762 = cond_wire472_out;
wire _guard11763 = _guard11761 & _guard11762;
wire _guard11764 = fsm_out == 1'd0;
wire _guard11765 = _guard11763 & _guard11764;
wire _guard11766 = _guard11760 | _guard11765;
wire _guard11767 = early_reset_static_par0_go_out;
wire _guard11768 = _guard11766 & _guard11767;
wire _guard11769 = cond_wire422_out;
wire _guard11770 = early_reset_static_par0_go_out;
wire _guard11771 = _guard11769 & _guard11770;
wire _guard11772 = cond_wire422_out;
wire _guard11773 = early_reset_static_par0_go_out;
wire _guard11774 = _guard11772 & _guard11773;
wire _guard11775 = cond_wire512_out;
wire _guard11776 = early_reset_static_par0_go_out;
wire _guard11777 = _guard11775 & _guard11776;
wire _guard11778 = cond_wire510_out;
wire _guard11779 = early_reset_static_par0_go_out;
wire _guard11780 = _guard11778 & _guard11779;
wire _guard11781 = fsm_out == 1'd0;
wire _guard11782 = cond_wire510_out;
wire _guard11783 = _guard11781 & _guard11782;
wire _guard11784 = fsm_out == 1'd0;
wire _guard11785 = _guard11783 & _guard11784;
wire _guard11786 = fsm_out == 1'd0;
wire _guard11787 = cond_wire512_out;
wire _guard11788 = _guard11786 & _guard11787;
wire _guard11789 = fsm_out == 1'd0;
wire _guard11790 = _guard11788 & _guard11789;
wire _guard11791 = _guard11785 | _guard11790;
wire _guard11792 = early_reset_static_par0_go_out;
wire _guard11793 = _guard11791 & _guard11792;
wire _guard11794 = fsm_out == 1'd0;
wire _guard11795 = cond_wire510_out;
wire _guard11796 = _guard11794 & _guard11795;
wire _guard11797 = fsm_out == 1'd0;
wire _guard11798 = _guard11796 & _guard11797;
wire _guard11799 = fsm_out == 1'd0;
wire _guard11800 = cond_wire512_out;
wire _guard11801 = _guard11799 & _guard11800;
wire _guard11802 = fsm_out == 1'd0;
wire _guard11803 = _guard11801 & _guard11802;
wire _guard11804 = _guard11798 | _guard11803;
wire _guard11805 = early_reset_static_par0_go_out;
wire _guard11806 = _guard11804 & _guard11805;
wire _guard11807 = fsm_out == 1'd0;
wire _guard11808 = cond_wire510_out;
wire _guard11809 = _guard11807 & _guard11808;
wire _guard11810 = fsm_out == 1'd0;
wire _guard11811 = _guard11809 & _guard11810;
wire _guard11812 = fsm_out == 1'd0;
wire _guard11813 = cond_wire512_out;
wire _guard11814 = _guard11812 & _guard11813;
wire _guard11815 = fsm_out == 1'd0;
wire _guard11816 = _guard11814 & _guard11815;
wire _guard11817 = _guard11811 | _guard11816;
wire _guard11818 = early_reset_static_par0_go_out;
wire _guard11819 = _guard11817 & _guard11818;
wire _guard11820 = cond_wire537_out;
wire _guard11821 = early_reset_static_par0_go_out;
wire _guard11822 = _guard11820 & _guard11821;
wire _guard11823 = cond_wire535_out;
wire _guard11824 = early_reset_static_par0_go_out;
wire _guard11825 = _guard11823 & _guard11824;
wire _guard11826 = fsm_out == 1'd0;
wire _guard11827 = cond_wire535_out;
wire _guard11828 = _guard11826 & _guard11827;
wire _guard11829 = fsm_out == 1'd0;
wire _guard11830 = _guard11828 & _guard11829;
wire _guard11831 = fsm_out == 1'd0;
wire _guard11832 = cond_wire537_out;
wire _guard11833 = _guard11831 & _guard11832;
wire _guard11834 = fsm_out == 1'd0;
wire _guard11835 = _guard11833 & _guard11834;
wire _guard11836 = _guard11830 | _guard11835;
wire _guard11837 = early_reset_static_par0_go_out;
wire _guard11838 = _guard11836 & _guard11837;
wire _guard11839 = fsm_out == 1'd0;
wire _guard11840 = cond_wire535_out;
wire _guard11841 = _guard11839 & _guard11840;
wire _guard11842 = fsm_out == 1'd0;
wire _guard11843 = _guard11841 & _guard11842;
wire _guard11844 = fsm_out == 1'd0;
wire _guard11845 = cond_wire537_out;
wire _guard11846 = _guard11844 & _guard11845;
wire _guard11847 = fsm_out == 1'd0;
wire _guard11848 = _guard11846 & _guard11847;
wire _guard11849 = _guard11843 | _guard11848;
wire _guard11850 = early_reset_static_par0_go_out;
wire _guard11851 = _guard11849 & _guard11850;
wire _guard11852 = fsm_out == 1'd0;
wire _guard11853 = cond_wire535_out;
wire _guard11854 = _guard11852 & _guard11853;
wire _guard11855 = fsm_out == 1'd0;
wire _guard11856 = _guard11854 & _guard11855;
wire _guard11857 = fsm_out == 1'd0;
wire _guard11858 = cond_wire537_out;
wire _guard11859 = _guard11857 & _guard11858;
wire _guard11860 = fsm_out == 1'd0;
wire _guard11861 = _guard11859 & _guard11860;
wire _guard11862 = _guard11856 | _guard11861;
wire _guard11863 = early_reset_static_par0_go_out;
wire _guard11864 = _guard11862 & _guard11863;
wire _guard11865 = cond_wire548_out;
wire _guard11866 = early_reset_static_par0_go_out;
wire _guard11867 = _guard11865 & _guard11866;
wire _guard11868 = cond_wire548_out;
wire _guard11869 = early_reset_static_par0_go_out;
wire _guard11870 = _guard11868 & _guard11869;
wire _guard11871 = cond_wire557_out;
wire _guard11872 = early_reset_static_par0_go_out;
wire _guard11873 = _guard11871 & _guard11872;
wire _guard11874 = cond_wire555_out;
wire _guard11875 = early_reset_static_par0_go_out;
wire _guard11876 = _guard11874 & _guard11875;
wire _guard11877 = fsm_out == 1'd0;
wire _guard11878 = cond_wire555_out;
wire _guard11879 = _guard11877 & _guard11878;
wire _guard11880 = fsm_out == 1'd0;
wire _guard11881 = _guard11879 & _guard11880;
wire _guard11882 = fsm_out == 1'd0;
wire _guard11883 = cond_wire557_out;
wire _guard11884 = _guard11882 & _guard11883;
wire _guard11885 = fsm_out == 1'd0;
wire _guard11886 = _guard11884 & _guard11885;
wire _guard11887 = _guard11881 | _guard11886;
wire _guard11888 = early_reset_static_par0_go_out;
wire _guard11889 = _guard11887 & _guard11888;
wire _guard11890 = fsm_out == 1'd0;
wire _guard11891 = cond_wire555_out;
wire _guard11892 = _guard11890 & _guard11891;
wire _guard11893 = fsm_out == 1'd0;
wire _guard11894 = _guard11892 & _guard11893;
wire _guard11895 = fsm_out == 1'd0;
wire _guard11896 = cond_wire557_out;
wire _guard11897 = _guard11895 & _guard11896;
wire _guard11898 = fsm_out == 1'd0;
wire _guard11899 = _guard11897 & _guard11898;
wire _guard11900 = _guard11894 | _guard11899;
wire _guard11901 = early_reset_static_par0_go_out;
wire _guard11902 = _guard11900 & _guard11901;
wire _guard11903 = fsm_out == 1'd0;
wire _guard11904 = cond_wire555_out;
wire _guard11905 = _guard11903 & _guard11904;
wire _guard11906 = fsm_out == 1'd0;
wire _guard11907 = _guard11905 & _guard11906;
wire _guard11908 = fsm_out == 1'd0;
wire _guard11909 = cond_wire557_out;
wire _guard11910 = _guard11908 & _guard11909;
wire _guard11911 = fsm_out == 1'd0;
wire _guard11912 = _guard11910 & _guard11911;
wire _guard11913 = _guard11907 | _guard11912;
wire _guard11914 = early_reset_static_par0_go_out;
wire _guard11915 = _guard11913 & _guard11914;
wire _guard11916 = cond_wire503_out;
wire _guard11917 = early_reset_static_par0_go_out;
wire _guard11918 = _guard11916 & _guard11917;
wire _guard11919 = cond_wire503_out;
wire _guard11920 = early_reset_static_par0_go_out;
wire _guard11921 = _guard11919 & _guard11920;
wire _guard11922 = cond_wire564_out;
wire _guard11923 = early_reset_static_par0_go_out;
wire _guard11924 = _guard11922 & _guard11923;
wire _guard11925 = cond_wire564_out;
wire _guard11926 = early_reset_static_par0_go_out;
wire _guard11927 = _guard11925 & _guard11926;
wire _guard11928 = cond_wire527_out;
wire _guard11929 = early_reset_static_par0_go_out;
wire _guard11930 = _guard11928 & _guard11929;
wire _guard11931 = cond_wire527_out;
wire _guard11932 = early_reset_static_par0_go_out;
wire _guard11933 = _guard11931 & _guard11932;
wire _guard11934 = cond_wire540_out;
wire _guard11935 = early_reset_static_par0_go_out;
wire _guard11936 = _guard11934 & _guard11935;
wire _guard11937 = cond_wire540_out;
wire _guard11938 = early_reset_static_par0_go_out;
wire _guard11939 = _guard11937 & _guard11938;
wire _guard11940 = cond_wire626_out;
wire _guard11941 = early_reset_static_par0_go_out;
wire _guard11942 = _guard11940 & _guard11941;
wire _guard11943 = cond_wire624_out;
wire _guard11944 = early_reset_static_par0_go_out;
wire _guard11945 = _guard11943 & _guard11944;
wire _guard11946 = fsm_out == 1'd0;
wire _guard11947 = cond_wire624_out;
wire _guard11948 = _guard11946 & _guard11947;
wire _guard11949 = fsm_out == 1'd0;
wire _guard11950 = _guard11948 & _guard11949;
wire _guard11951 = fsm_out == 1'd0;
wire _guard11952 = cond_wire626_out;
wire _guard11953 = _guard11951 & _guard11952;
wire _guard11954 = fsm_out == 1'd0;
wire _guard11955 = _guard11953 & _guard11954;
wire _guard11956 = _guard11950 | _guard11955;
wire _guard11957 = early_reset_static_par0_go_out;
wire _guard11958 = _guard11956 & _guard11957;
wire _guard11959 = fsm_out == 1'd0;
wire _guard11960 = cond_wire624_out;
wire _guard11961 = _guard11959 & _guard11960;
wire _guard11962 = fsm_out == 1'd0;
wire _guard11963 = _guard11961 & _guard11962;
wire _guard11964 = fsm_out == 1'd0;
wire _guard11965 = cond_wire626_out;
wire _guard11966 = _guard11964 & _guard11965;
wire _guard11967 = fsm_out == 1'd0;
wire _guard11968 = _guard11966 & _guard11967;
wire _guard11969 = _guard11963 | _guard11968;
wire _guard11970 = early_reset_static_par0_go_out;
wire _guard11971 = _guard11969 & _guard11970;
wire _guard11972 = fsm_out == 1'd0;
wire _guard11973 = cond_wire624_out;
wire _guard11974 = _guard11972 & _guard11973;
wire _guard11975 = fsm_out == 1'd0;
wire _guard11976 = _guard11974 & _guard11975;
wire _guard11977 = fsm_out == 1'd0;
wire _guard11978 = cond_wire626_out;
wire _guard11979 = _guard11977 & _guard11978;
wire _guard11980 = fsm_out == 1'd0;
wire _guard11981 = _guard11979 & _guard11980;
wire _guard11982 = _guard11976 | _guard11981;
wire _guard11983 = early_reset_static_par0_go_out;
wire _guard11984 = _guard11982 & _guard11983;
wire _guard11985 = cond_wire633_out;
wire _guard11986 = early_reset_static_par0_go_out;
wire _guard11987 = _guard11985 & _guard11986;
wire _guard11988 = cond_wire633_out;
wire _guard11989 = early_reset_static_par0_go_out;
wire _guard11990 = _guard11988 & _guard11989;
wire _guard11991 = cond_wire637_out;
wire _guard11992 = early_reset_static_par0_go_out;
wire _guard11993 = _guard11991 & _guard11992;
wire _guard11994 = cond_wire637_out;
wire _guard11995 = early_reset_static_par0_go_out;
wire _guard11996 = _guard11994 & _guard11995;
wire _guard11997 = cond_wire596_out;
wire _guard11998 = early_reset_static_par0_go_out;
wire _guard11999 = _guard11997 & _guard11998;
wire _guard12000 = cond_wire596_out;
wire _guard12001 = early_reset_static_par0_go_out;
wire _guard12002 = _guard12000 & _guard12001;
wire _guard12003 = cond_wire601_out;
wire _guard12004 = early_reset_static_par0_go_out;
wire _guard12005 = _guard12003 & _guard12004;
wire _guard12006 = cond_wire601_out;
wire _guard12007 = early_reset_static_par0_go_out;
wire _guard12008 = _guard12006 & _guard12007;
wire _guard12009 = cond_wire621_out;
wire _guard12010 = early_reset_static_par0_go_out;
wire _guard12011 = _guard12009 & _guard12010;
wire _guard12012 = cond_wire621_out;
wire _guard12013 = early_reset_static_par0_go_out;
wire _guard12014 = _guard12012 & _guard12013;
wire _guard12015 = cond_wire702_out;
wire _guard12016 = early_reset_static_par0_go_out;
wire _guard12017 = _guard12015 & _guard12016;
wire _guard12018 = cond_wire702_out;
wire _guard12019 = early_reset_static_par0_go_out;
wire _guard12020 = _guard12018 & _guard12019;
wire _guard12021 = cond_wire715_out;
wire _guard12022 = early_reset_static_par0_go_out;
wire _guard12023 = _guard12021 & _guard12022;
wire _guard12024 = cond_wire713_out;
wire _guard12025 = early_reset_static_par0_go_out;
wire _guard12026 = _guard12024 & _guard12025;
wire _guard12027 = fsm_out == 1'd0;
wire _guard12028 = cond_wire713_out;
wire _guard12029 = _guard12027 & _guard12028;
wire _guard12030 = fsm_out == 1'd0;
wire _guard12031 = _guard12029 & _guard12030;
wire _guard12032 = fsm_out == 1'd0;
wire _guard12033 = cond_wire715_out;
wire _guard12034 = _guard12032 & _guard12033;
wire _guard12035 = fsm_out == 1'd0;
wire _guard12036 = _guard12034 & _guard12035;
wire _guard12037 = _guard12031 | _guard12036;
wire _guard12038 = early_reset_static_par0_go_out;
wire _guard12039 = _guard12037 & _guard12038;
wire _guard12040 = fsm_out == 1'd0;
wire _guard12041 = cond_wire713_out;
wire _guard12042 = _guard12040 & _guard12041;
wire _guard12043 = fsm_out == 1'd0;
wire _guard12044 = _guard12042 & _guard12043;
wire _guard12045 = fsm_out == 1'd0;
wire _guard12046 = cond_wire715_out;
wire _guard12047 = _guard12045 & _guard12046;
wire _guard12048 = fsm_out == 1'd0;
wire _guard12049 = _guard12047 & _guard12048;
wire _guard12050 = _guard12044 | _guard12049;
wire _guard12051 = early_reset_static_par0_go_out;
wire _guard12052 = _guard12050 & _guard12051;
wire _guard12053 = fsm_out == 1'd0;
wire _guard12054 = cond_wire713_out;
wire _guard12055 = _guard12053 & _guard12054;
wire _guard12056 = fsm_out == 1'd0;
wire _guard12057 = _guard12055 & _guard12056;
wire _guard12058 = fsm_out == 1'd0;
wire _guard12059 = cond_wire715_out;
wire _guard12060 = _guard12058 & _guard12059;
wire _guard12061 = fsm_out == 1'd0;
wire _guard12062 = _guard12060 & _guard12061;
wire _guard12063 = _guard12057 | _guard12062;
wire _guard12064 = early_reset_static_par0_go_out;
wire _guard12065 = _guard12063 & _guard12064;
wire _guard12066 = cond_wire670_out;
wire _guard12067 = early_reset_static_par0_go_out;
wire _guard12068 = _guard12066 & _guard12067;
wire _guard12069 = cond_wire670_out;
wire _guard12070 = early_reset_static_par0_go_out;
wire _guard12071 = _guard12069 & _guard12070;
wire _guard12072 = cond_wire756_out;
wire _guard12073 = early_reset_static_par0_go_out;
wire _guard12074 = _guard12072 & _guard12073;
wire _guard12075 = cond_wire754_out;
wire _guard12076 = early_reset_static_par0_go_out;
wire _guard12077 = _guard12075 & _guard12076;
wire _guard12078 = fsm_out == 1'd0;
wire _guard12079 = cond_wire754_out;
wire _guard12080 = _guard12078 & _guard12079;
wire _guard12081 = fsm_out == 1'd0;
wire _guard12082 = _guard12080 & _guard12081;
wire _guard12083 = fsm_out == 1'd0;
wire _guard12084 = cond_wire756_out;
wire _guard12085 = _guard12083 & _guard12084;
wire _guard12086 = fsm_out == 1'd0;
wire _guard12087 = _guard12085 & _guard12086;
wire _guard12088 = _guard12082 | _guard12087;
wire _guard12089 = early_reset_static_par0_go_out;
wire _guard12090 = _guard12088 & _guard12089;
wire _guard12091 = fsm_out == 1'd0;
wire _guard12092 = cond_wire754_out;
wire _guard12093 = _guard12091 & _guard12092;
wire _guard12094 = fsm_out == 1'd0;
wire _guard12095 = _guard12093 & _guard12094;
wire _guard12096 = fsm_out == 1'd0;
wire _guard12097 = cond_wire756_out;
wire _guard12098 = _guard12096 & _guard12097;
wire _guard12099 = fsm_out == 1'd0;
wire _guard12100 = _guard12098 & _guard12099;
wire _guard12101 = _guard12095 | _guard12100;
wire _guard12102 = early_reset_static_par0_go_out;
wire _guard12103 = _guard12101 & _guard12102;
wire _guard12104 = fsm_out == 1'd0;
wire _guard12105 = cond_wire754_out;
wire _guard12106 = _guard12104 & _guard12105;
wire _guard12107 = fsm_out == 1'd0;
wire _guard12108 = _guard12106 & _guard12107;
wire _guard12109 = fsm_out == 1'd0;
wire _guard12110 = cond_wire756_out;
wire _guard12111 = _guard12109 & _guard12110;
wire _guard12112 = fsm_out == 1'd0;
wire _guard12113 = _guard12111 & _guard12112;
wire _guard12114 = _guard12108 | _guard12113;
wire _guard12115 = early_reset_static_par0_go_out;
wire _guard12116 = _guard12114 & _guard12115;
wire _guard12117 = cond_wire760_out;
wire _guard12118 = early_reset_static_par0_go_out;
wire _guard12119 = _guard12117 & _guard12118;
wire _guard12120 = cond_wire758_out;
wire _guard12121 = early_reset_static_par0_go_out;
wire _guard12122 = _guard12120 & _guard12121;
wire _guard12123 = fsm_out == 1'd0;
wire _guard12124 = cond_wire758_out;
wire _guard12125 = _guard12123 & _guard12124;
wire _guard12126 = fsm_out == 1'd0;
wire _guard12127 = _guard12125 & _guard12126;
wire _guard12128 = fsm_out == 1'd0;
wire _guard12129 = cond_wire760_out;
wire _guard12130 = _guard12128 & _guard12129;
wire _guard12131 = fsm_out == 1'd0;
wire _guard12132 = _guard12130 & _guard12131;
wire _guard12133 = _guard12127 | _guard12132;
wire _guard12134 = early_reset_static_par0_go_out;
wire _guard12135 = _guard12133 & _guard12134;
wire _guard12136 = fsm_out == 1'd0;
wire _guard12137 = cond_wire758_out;
wire _guard12138 = _guard12136 & _guard12137;
wire _guard12139 = fsm_out == 1'd0;
wire _guard12140 = _guard12138 & _guard12139;
wire _guard12141 = fsm_out == 1'd0;
wire _guard12142 = cond_wire760_out;
wire _guard12143 = _guard12141 & _guard12142;
wire _guard12144 = fsm_out == 1'd0;
wire _guard12145 = _guard12143 & _guard12144;
wire _guard12146 = _guard12140 | _guard12145;
wire _guard12147 = early_reset_static_par0_go_out;
wire _guard12148 = _guard12146 & _guard12147;
wire _guard12149 = fsm_out == 1'd0;
wire _guard12150 = cond_wire758_out;
wire _guard12151 = _guard12149 & _guard12150;
wire _guard12152 = fsm_out == 1'd0;
wire _guard12153 = _guard12151 & _guard12152;
wire _guard12154 = fsm_out == 1'd0;
wire _guard12155 = cond_wire760_out;
wire _guard12156 = _guard12154 & _guard12155;
wire _guard12157 = fsm_out == 1'd0;
wire _guard12158 = _guard12156 & _guard12157;
wire _guard12159 = _guard12153 | _guard12158;
wire _guard12160 = early_reset_static_par0_go_out;
wire _guard12161 = _guard12159 & _guard12160;
wire _guard12162 = cond_wire735_out;
wire _guard12163 = early_reset_static_par0_go_out;
wire _guard12164 = _guard12162 & _guard12163;
wire _guard12165 = cond_wire735_out;
wire _guard12166 = early_reset_static_par0_go_out;
wire _guard12167 = _guard12165 & _guard12166;
wire _guard12168 = cond_wire809_out;
wire _guard12169 = early_reset_static_par0_go_out;
wire _guard12170 = _guard12168 & _guard12169;
wire _guard12171 = cond_wire807_out;
wire _guard12172 = early_reset_static_par0_go_out;
wire _guard12173 = _guard12171 & _guard12172;
wire _guard12174 = fsm_out == 1'd0;
wire _guard12175 = cond_wire807_out;
wire _guard12176 = _guard12174 & _guard12175;
wire _guard12177 = fsm_out == 1'd0;
wire _guard12178 = _guard12176 & _guard12177;
wire _guard12179 = fsm_out == 1'd0;
wire _guard12180 = cond_wire809_out;
wire _guard12181 = _guard12179 & _guard12180;
wire _guard12182 = fsm_out == 1'd0;
wire _guard12183 = _guard12181 & _guard12182;
wire _guard12184 = _guard12178 | _guard12183;
wire _guard12185 = early_reset_static_par0_go_out;
wire _guard12186 = _guard12184 & _guard12185;
wire _guard12187 = fsm_out == 1'd0;
wire _guard12188 = cond_wire807_out;
wire _guard12189 = _guard12187 & _guard12188;
wire _guard12190 = fsm_out == 1'd0;
wire _guard12191 = _guard12189 & _guard12190;
wire _guard12192 = fsm_out == 1'd0;
wire _guard12193 = cond_wire809_out;
wire _guard12194 = _guard12192 & _guard12193;
wire _guard12195 = fsm_out == 1'd0;
wire _guard12196 = _guard12194 & _guard12195;
wire _guard12197 = _guard12191 | _guard12196;
wire _guard12198 = early_reset_static_par0_go_out;
wire _guard12199 = _guard12197 & _guard12198;
wire _guard12200 = fsm_out == 1'd0;
wire _guard12201 = cond_wire807_out;
wire _guard12202 = _guard12200 & _guard12201;
wire _guard12203 = fsm_out == 1'd0;
wire _guard12204 = _guard12202 & _guard12203;
wire _guard12205 = fsm_out == 1'd0;
wire _guard12206 = cond_wire809_out;
wire _guard12207 = _guard12205 & _guard12206;
wire _guard12208 = fsm_out == 1'd0;
wire _guard12209 = _guard12207 & _guard12208;
wire _guard12210 = _guard12204 | _guard12209;
wire _guard12211 = early_reset_static_par0_go_out;
wire _guard12212 = _guard12210 & _guard12211;
wire _guard12213 = cond_wire813_out;
wire _guard12214 = early_reset_static_par0_go_out;
wire _guard12215 = _guard12213 & _guard12214;
wire _guard12216 = cond_wire811_out;
wire _guard12217 = early_reset_static_par0_go_out;
wire _guard12218 = _guard12216 & _guard12217;
wire _guard12219 = fsm_out == 1'd0;
wire _guard12220 = cond_wire811_out;
wire _guard12221 = _guard12219 & _guard12220;
wire _guard12222 = fsm_out == 1'd0;
wire _guard12223 = _guard12221 & _guard12222;
wire _guard12224 = fsm_out == 1'd0;
wire _guard12225 = cond_wire813_out;
wire _guard12226 = _guard12224 & _guard12225;
wire _guard12227 = fsm_out == 1'd0;
wire _guard12228 = _guard12226 & _guard12227;
wire _guard12229 = _guard12223 | _guard12228;
wire _guard12230 = early_reset_static_par0_go_out;
wire _guard12231 = _guard12229 & _guard12230;
wire _guard12232 = fsm_out == 1'd0;
wire _guard12233 = cond_wire811_out;
wire _guard12234 = _guard12232 & _guard12233;
wire _guard12235 = fsm_out == 1'd0;
wire _guard12236 = _guard12234 & _guard12235;
wire _guard12237 = fsm_out == 1'd0;
wire _guard12238 = cond_wire813_out;
wire _guard12239 = _guard12237 & _guard12238;
wire _guard12240 = fsm_out == 1'd0;
wire _guard12241 = _guard12239 & _guard12240;
wire _guard12242 = _guard12236 | _guard12241;
wire _guard12243 = early_reset_static_par0_go_out;
wire _guard12244 = _guard12242 & _guard12243;
wire _guard12245 = fsm_out == 1'd0;
wire _guard12246 = cond_wire811_out;
wire _guard12247 = _guard12245 & _guard12246;
wire _guard12248 = fsm_out == 1'd0;
wire _guard12249 = _guard12247 & _guard12248;
wire _guard12250 = fsm_out == 1'd0;
wire _guard12251 = cond_wire813_out;
wire _guard12252 = _guard12250 & _guard12251;
wire _guard12253 = fsm_out == 1'd0;
wire _guard12254 = _guard12252 & _guard12253;
wire _guard12255 = _guard12249 | _guard12254;
wire _guard12256 = early_reset_static_par0_go_out;
wire _guard12257 = _guard12255 & _guard12256;
wire _guard12258 = cond_wire828_out;
wire _guard12259 = early_reset_static_par0_go_out;
wire _guard12260 = _guard12258 & _guard12259;
wire _guard12261 = cond_wire828_out;
wire _guard12262 = early_reset_static_par0_go_out;
wire _guard12263 = _guard12261 & _guard12262;
wire _guard12264 = cond_wire775_out;
wire _guard12265 = early_reset_static_par0_go_out;
wire _guard12266 = _guard12264 & _guard12265;
wire _guard12267 = cond_wire775_out;
wire _guard12268 = early_reset_static_par0_go_out;
wire _guard12269 = _guard12267 & _guard12268;
wire _guard12270 = cond_wire779_out;
wire _guard12271 = early_reset_static_par0_go_out;
wire _guard12272 = _guard12270 & _guard12271;
wire _guard12273 = cond_wire779_out;
wire _guard12274 = early_reset_static_par0_go_out;
wire _guard12275 = _guard12273 & _guard12274;
wire _guard12276 = cond_wire862_out;
wire _guard12277 = early_reset_static_par0_go_out;
wire _guard12278 = _guard12276 & _guard12277;
wire _guard12279 = cond_wire860_out;
wire _guard12280 = early_reset_static_par0_go_out;
wire _guard12281 = _guard12279 & _guard12280;
wire _guard12282 = fsm_out == 1'd0;
wire _guard12283 = cond_wire860_out;
wire _guard12284 = _guard12282 & _guard12283;
wire _guard12285 = fsm_out == 1'd0;
wire _guard12286 = _guard12284 & _guard12285;
wire _guard12287 = fsm_out == 1'd0;
wire _guard12288 = cond_wire862_out;
wire _guard12289 = _guard12287 & _guard12288;
wire _guard12290 = fsm_out == 1'd0;
wire _guard12291 = _guard12289 & _guard12290;
wire _guard12292 = _guard12286 | _guard12291;
wire _guard12293 = early_reset_static_par0_go_out;
wire _guard12294 = _guard12292 & _guard12293;
wire _guard12295 = fsm_out == 1'd0;
wire _guard12296 = cond_wire860_out;
wire _guard12297 = _guard12295 & _guard12296;
wire _guard12298 = fsm_out == 1'd0;
wire _guard12299 = _guard12297 & _guard12298;
wire _guard12300 = fsm_out == 1'd0;
wire _guard12301 = cond_wire862_out;
wire _guard12302 = _guard12300 & _guard12301;
wire _guard12303 = fsm_out == 1'd0;
wire _guard12304 = _guard12302 & _guard12303;
wire _guard12305 = _guard12299 | _guard12304;
wire _guard12306 = early_reset_static_par0_go_out;
wire _guard12307 = _guard12305 & _guard12306;
wire _guard12308 = fsm_out == 1'd0;
wire _guard12309 = cond_wire860_out;
wire _guard12310 = _guard12308 & _guard12309;
wire _guard12311 = fsm_out == 1'd0;
wire _guard12312 = _guard12310 & _guard12311;
wire _guard12313 = fsm_out == 1'd0;
wire _guard12314 = cond_wire862_out;
wire _guard12315 = _guard12313 & _guard12314;
wire _guard12316 = fsm_out == 1'd0;
wire _guard12317 = _guard12315 & _guard12316;
wire _guard12318 = _guard12312 | _guard12317;
wire _guard12319 = early_reset_static_par0_go_out;
wire _guard12320 = _guard12318 & _guard12319;
wire _guard12321 = cond_wire874_out;
wire _guard12322 = early_reset_static_par0_go_out;
wire _guard12323 = _guard12321 & _guard12322;
wire _guard12324 = cond_wire872_out;
wire _guard12325 = early_reset_static_par0_go_out;
wire _guard12326 = _guard12324 & _guard12325;
wire _guard12327 = fsm_out == 1'd0;
wire _guard12328 = cond_wire872_out;
wire _guard12329 = _guard12327 & _guard12328;
wire _guard12330 = fsm_out == 1'd0;
wire _guard12331 = _guard12329 & _guard12330;
wire _guard12332 = fsm_out == 1'd0;
wire _guard12333 = cond_wire874_out;
wire _guard12334 = _guard12332 & _guard12333;
wire _guard12335 = fsm_out == 1'd0;
wire _guard12336 = _guard12334 & _guard12335;
wire _guard12337 = _guard12331 | _guard12336;
wire _guard12338 = early_reset_static_par0_go_out;
wire _guard12339 = _guard12337 & _guard12338;
wire _guard12340 = fsm_out == 1'd0;
wire _guard12341 = cond_wire872_out;
wire _guard12342 = _guard12340 & _guard12341;
wire _guard12343 = fsm_out == 1'd0;
wire _guard12344 = _guard12342 & _guard12343;
wire _guard12345 = fsm_out == 1'd0;
wire _guard12346 = cond_wire874_out;
wire _guard12347 = _guard12345 & _guard12346;
wire _guard12348 = fsm_out == 1'd0;
wire _guard12349 = _guard12347 & _guard12348;
wire _guard12350 = _guard12344 | _guard12349;
wire _guard12351 = early_reset_static_par0_go_out;
wire _guard12352 = _guard12350 & _guard12351;
wire _guard12353 = fsm_out == 1'd0;
wire _guard12354 = cond_wire872_out;
wire _guard12355 = _guard12353 & _guard12354;
wire _guard12356 = fsm_out == 1'd0;
wire _guard12357 = _guard12355 & _guard12356;
wire _guard12358 = fsm_out == 1'd0;
wire _guard12359 = cond_wire874_out;
wire _guard12360 = _guard12358 & _guard12359;
wire _guard12361 = fsm_out == 1'd0;
wire _guard12362 = _guard12360 & _guard12361;
wire _guard12363 = _guard12357 | _guard12362;
wire _guard12364 = early_reset_static_par0_go_out;
wire _guard12365 = _guard12363 & _guard12364;
wire _guard12366 = cond_wire885_out;
wire _guard12367 = early_reset_static_par0_go_out;
wire _guard12368 = _guard12366 & _guard12367;
wire _guard12369 = cond_wire885_out;
wire _guard12370 = early_reset_static_par0_go_out;
wire _guard12371 = _guard12369 & _guard12370;
wire _guard12372 = cond_wire889_out;
wire _guard12373 = early_reset_static_par0_go_out;
wire _guard12374 = _guard12372 & _guard12373;
wire _guard12375 = cond_wire889_out;
wire _guard12376 = early_reset_static_par0_go_out;
wire _guard12377 = _guard12375 & _guard12376;
wire _guard12378 = cond_wire914_out;
wire _guard12379 = early_reset_static_par0_go_out;
wire _guard12380 = _guard12378 & _guard12379;
wire _guard12381 = cond_wire912_out;
wire _guard12382 = early_reset_static_par0_go_out;
wire _guard12383 = _guard12381 & _guard12382;
wire _guard12384 = fsm_out == 1'd0;
wire _guard12385 = cond_wire912_out;
wire _guard12386 = _guard12384 & _guard12385;
wire _guard12387 = fsm_out == 1'd0;
wire _guard12388 = _guard12386 & _guard12387;
wire _guard12389 = fsm_out == 1'd0;
wire _guard12390 = cond_wire914_out;
wire _guard12391 = _guard12389 & _guard12390;
wire _guard12392 = fsm_out == 1'd0;
wire _guard12393 = _guard12391 & _guard12392;
wire _guard12394 = _guard12388 | _guard12393;
wire _guard12395 = early_reset_static_par0_go_out;
wire _guard12396 = _guard12394 & _guard12395;
wire _guard12397 = fsm_out == 1'd0;
wire _guard12398 = cond_wire912_out;
wire _guard12399 = _guard12397 & _guard12398;
wire _guard12400 = fsm_out == 1'd0;
wire _guard12401 = _guard12399 & _guard12400;
wire _guard12402 = fsm_out == 1'd0;
wire _guard12403 = cond_wire914_out;
wire _guard12404 = _guard12402 & _guard12403;
wire _guard12405 = fsm_out == 1'd0;
wire _guard12406 = _guard12404 & _guard12405;
wire _guard12407 = _guard12401 | _guard12406;
wire _guard12408 = early_reset_static_par0_go_out;
wire _guard12409 = _guard12407 & _guard12408;
wire _guard12410 = fsm_out == 1'd0;
wire _guard12411 = cond_wire912_out;
wire _guard12412 = _guard12410 & _guard12411;
wire _guard12413 = fsm_out == 1'd0;
wire _guard12414 = _guard12412 & _guard12413;
wire _guard12415 = fsm_out == 1'd0;
wire _guard12416 = cond_wire914_out;
wire _guard12417 = _guard12415 & _guard12416;
wire _guard12418 = fsm_out == 1'd0;
wire _guard12419 = _guard12417 & _guard12418;
wire _guard12420 = _guard12414 | _guard12419;
wire _guard12421 = early_reset_static_par0_go_out;
wire _guard12422 = _guard12420 & _guard12421;
wire _guard12423 = cond_wire909_out;
wire _guard12424 = early_reset_static_par0_go_out;
wire _guard12425 = _guard12423 & _guard12424;
wire _guard12426 = cond_wire909_out;
wire _guard12427 = early_reset_static_par0_go_out;
wire _guard12428 = _guard12426 & _guard12427;
wire _guard12429 = cond_wire934_out;
wire _guard12430 = early_reset_static_par0_go_out;
wire _guard12431 = _guard12429 & _guard12430;
wire _guard12432 = cond_wire934_out;
wire _guard12433 = early_reset_static_par0_go_out;
wire _guard12434 = _guard12432 & _guard12433;
wire _guard12435 = cond_wire946_out;
wire _guard12436 = early_reset_static_par0_go_out;
wire _guard12437 = _guard12435 & _guard12436;
wire _guard12438 = cond_wire946_out;
wire _guard12439 = early_reset_static_par0_go_out;
wire _guard12440 = _guard12438 & _guard12439;
wire _guard12441 = cond_wire1015_out;
wire _guard12442 = early_reset_static_par0_go_out;
wire _guard12443 = _guard12441 & _guard12442;
wire _guard12444 = cond_wire1015_out;
wire _guard12445 = early_reset_static_par0_go_out;
wire _guard12446 = _guard12444 & _guard12445;
wire _guard12447 = cond_wire1044_out;
wire _guard12448 = early_reset_static_par0_go_out;
wire _guard12449 = _guard12447 & _guard12448;
wire _guard12450 = cond_wire1042_out;
wire _guard12451 = early_reset_static_par0_go_out;
wire _guard12452 = _guard12450 & _guard12451;
wire _guard12453 = fsm_out == 1'd0;
wire _guard12454 = cond_wire1042_out;
wire _guard12455 = _guard12453 & _guard12454;
wire _guard12456 = fsm_out == 1'd0;
wire _guard12457 = _guard12455 & _guard12456;
wire _guard12458 = fsm_out == 1'd0;
wire _guard12459 = cond_wire1044_out;
wire _guard12460 = _guard12458 & _guard12459;
wire _guard12461 = fsm_out == 1'd0;
wire _guard12462 = _guard12460 & _guard12461;
wire _guard12463 = _guard12457 | _guard12462;
wire _guard12464 = early_reset_static_par0_go_out;
wire _guard12465 = _guard12463 & _guard12464;
wire _guard12466 = fsm_out == 1'd0;
wire _guard12467 = cond_wire1042_out;
wire _guard12468 = _guard12466 & _guard12467;
wire _guard12469 = fsm_out == 1'd0;
wire _guard12470 = _guard12468 & _guard12469;
wire _guard12471 = fsm_out == 1'd0;
wire _guard12472 = cond_wire1044_out;
wire _guard12473 = _guard12471 & _guard12472;
wire _guard12474 = fsm_out == 1'd0;
wire _guard12475 = _guard12473 & _guard12474;
wire _guard12476 = _guard12470 | _guard12475;
wire _guard12477 = early_reset_static_par0_go_out;
wire _guard12478 = _guard12476 & _guard12477;
wire _guard12479 = fsm_out == 1'd0;
wire _guard12480 = cond_wire1042_out;
wire _guard12481 = _guard12479 & _guard12480;
wire _guard12482 = fsm_out == 1'd0;
wire _guard12483 = _guard12481 & _guard12482;
wire _guard12484 = fsm_out == 1'd0;
wire _guard12485 = cond_wire1044_out;
wire _guard12486 = _guard12484 & _guard12485;
wire _guard12487 = fsm_out == 1'd0;
wire _guard12488 = _guard12486 & _guard12487;
wire _guard12489 = _guard12483 | _guard12488;
wire _guard12490 = early_reset_static_par0_go_out;
wire _guard12491 = _guard12489 & _guard12490;
wire _guard12492 = fsm0_out == 6'd0;
wire _guard12493 = early_reset_static_seq_go_out;
wire _guard12494 = _guard12492 & _guard12493;
wire _guard12495 = cond_wire_out;
wire _guard12496 = early_reset_static_par0_go_out;
wire _guard12497 = _guard12495 & _guard12496;
wire _guard12498 = _guard12494 | _guard12497;
wire _guard12499 = fsm0_out == 6'd0;
wire _guard12500 = early_reset_static_seq_go_out;
wire _guard12501 = _guard12499 & _guard12500;
wire _guard12502 = cond_wire_out;
wire _guard12503 = early_reset_static_par0_go_out;
wire _guard12504 = _guard12502 & _guard12503;
wire _guard12505 = fsm0_out == 6'd0;
wire _guard12506 = early_reset_static_seq_go_out;
wire _guard12507 = _guard12505 & _guard12506;
wire _guard12508 = cond_wire19_out;
wire _guard12509 = early_reset_static_par0_go_out;
wire _guard12510 = _guard12508 & _guard12509;
wire _guard12511 = _guard12507 | _guard12510;
wire _guard12512 = fsm0_out == 6'd0;
wire _guard12513 = early_reset_static_seq_go_out;
wire _guard12514 = _guard12512 & _guard12513;
wire _guard12515 = cond_wire19_out;
wire _guard12516 = early_reset_static_par0_go_out;
wire _guard12517 = _guard12515 & _guard12516;
wire _guard12518 = fsm0_out == 6'd0;
wire _guard12519 = early_reset_static_seq_go_out;
wire _guard12520 = _guard12518 & _guard12519;
wire _guard12521 = cond_wire29_out;
wire _guard12522 = early_reset_static_par0_go_out;
wire _guard12523 = _guard12521 & _guard12522;
wire _guard12524 = _guard12520 | _guard12523;
wire _guard12525 = fsm0_out == 6'd0;
wire _guard12526 = early_reset_static_seq_go_out;
wire _guard12527 = _guard12525 & _guard12526;
wire _guard12528 = cond_wire29_out;
wire _guard12529 = early_reset_static_par0_go_out;
wire _guard12530 = _guard12528 & _guard12529;
wire _guard12531 = fsm0_out == 6'd0;
wire _guard12532 = early_reset_static_seq_go_out;
wire _guard12533 = _guard12531 & _guard12532;
wire _guard12534 = cond_wire59_out;
wire _guard12535 = early_reset_static_par0_go_out;
wire _guard12536 = _guard12534 & _guard12535;
wire _guard12537 = _guard12533 | _guard12536;
wire _guard12538 = fsm0_out == 6'd0;
wire _guard12539 = early_reset_static_seq_go_out;
wire _guard12540 = _guard12538 & _guard12539;
wire _guard12541 = cond_wire59_out;
wire _guard12542 = early_reset_static_par0_go_out;
wire _guard12543 = _guard12541 & _guard12542;
wire _guard12544 = fsm0_out == 6'd0;
wire _guard12545 = early_reset_static_seq_go_out;
wire _guard12546 = _guard12544 & _guard12545;
wire _guard12547 = cond_wire69_out;
wire _guard12548 = early_reset_static_par0_go_out;
wire _guard12549 = _guard12547 & _guard12548;
wire _guard12550 = _guard12546 | _guard12549;
wire _guard12551 = fsm0_out == 6'd0;
wire _guard12552 = early_reset_static_seq_go_out;
wire _guard12553 = _guard12551 & _guard12552;
wire _guard12554 = cond_wire69_out;
wire _guard12555 = early_reset_static_par0_go_out;
wire _guard12556 = _guard12554 & _guard12555;
wire _guard12557 = fsm0_out == 6'd0;
wire _guard12558 = early_reset_static_seq_go_out;
wire _guard12559 = _guard12557 & _guard12558;
wire _guard12560 = cond_wire79_out;
wire _guard12561 = early_reset_static_par0_go_out;
wire _guard12562 = _guard12560 & _guard12561;
wire _guard12563 = _guard12559 | _guard12562;
wire _guard12564 = cond_wire79_out;
wire _guard12565 = early_reset_static_par0_go_out;
wire _guard12566 = _guard12564 & _guard12565;
wire _guard12567 = fsm0_out == 6'd0;
wire _guard12568 = early_reset_static_seq_go_out;
wire _guard12569 = _guard12567 & _guard12568;
wire _guard12570 = cond_wire339_out;
wire _guard12571 = early_reset_static_par0_go_out;
wire _guard12572 = _guard12570 & _guard12571;
wire _guard12573 = cond_wire339_out;
wire _guard12574 = early_reset_static_par0_go_out;
wire _guard12575 = _guard12573 & _guard12574;
wire _guard12576 = early_reset_static_par0_go_out;
wire _guard12577 = early_reset_static_par0_go_out;
wire _guard12578 = early_reset_static_par0_go_out;
wire _guard12579 = early_reset_static_par0_go_out;
wire _guard12580 = early_reset_static_par0_go_out;
wire _guard12581 = early_reset_static_par0_go_out;
wire _guard12582 = fsm0_out == 6'd0;
wire _guard12583 = early_reset_static_seq_go_out;
wire _guard12584 = _guard12582 & _guard12583;
wire _guard12585 = early_reset_static_par0_go_out;
wire _guard12586 = _guard12584 | _guard12585;
wire _guard12587 = early_reset_static_par0_go_out;
wire _guard12588 = fsm0_out == 6'd0;
wire _guard12589 = early_reset_static_seq_go_out;
wire _guard12590 = _guard12588 & _guard12589;
wire _guard12591 = early_reset_static_par0_go_out;
wire _guard12592 = early_reset_static_par0_go_out;
wire _guard12593 = early_reset_static_par0_go_out;
wire _guard12594 = early_reset_static_par0_go_out;
wire _guard12595 = early_reset_static_par0_go_out;
wire _guard12596 = early_reset_static_par0_go_out;
wire _guard12597 = early_reset_static_par0_go_out;
wire _guard12598 = early_reset_static_par0_go_out;
wire _guard12599 = early_reset_static_par0_go_out;
wire _guard12600 = early_reset_static_par0_go_out;
wire _guard12601 = early_reset_static_par0_go_out;
wire _guard12602 = early_reset_static_par0_go_out;
wire _guard12603 = fsm0_out == 6'd0;
wire _guard12604 = early_reset_static_seq_go_out;
wire _guard12605 = _guard12603 & _guard12604;
wire _guard12606 = early_reset_static_par0_go_out;
wire _guard12607 = _guard12605 | _guard12606;
wire _guard12608 = early_reset_static_par0_go_out;
wire _guard12609 = fsm0_out == 6'd0;
wire _guard12610 = early_reset_static_seq_go_out;
wire _guard12611 = _guard12609 & _guard12610;
wire _guard12612 = early_reset_static_par0_go_out;
wire _guard12613 = early_reset_static_par0_go_out;
wire _guard12614 = early_reset_static_par0_go_out;
wire _guard12615 = early_reset_static_par0_go_out;
wire _guard12616 = early_reset_static_par0_go_out;
wire _guard12617 = early_reset_static_par0_go_out;
wire _guard12618 = fsm0_out == 6'd0;
wire _guard12619 = early_reset_static_seq_go_out;
wire _guard12620 = _guard12618 & _guard12619;
wire _guard12621 = early_reset_static_par0_go_out;
wire _guard12622 = _guard12620 | _guard12621;
wire _guard12623 = early_reset_static_par0_go_out;
wire _guard12624 = fsm0_out == 6'd0;
wire _guard12625 = early_reset_static_seq_go_out;
wire _guard12626 = _guard12624 & _guard12625;
wire _guard12627 = early_reset_static_par0_go_out;
wire _guard12628 = early_reset_static_par0_go_out;
wire _guard12629 = fsm0_out == 6'd0;
wire _guard12630 = early_reset_static_seq_go_out;
wire _guard12631 = _guard12629 & _guard12630;
wire _guard12632 = early_reset_static_par0_go_out;
wire _guard12633 = _guard12631 | _guard12632;
wire _guard12634 = early_reset_static_par0_go_out;
wire _guard12635 = fsm0_out == 6'd0;
wire _guard12636 = early_reset_static_seq_go_out;
wire _guard12637 = _guard12635 & _guard12636;
wire _guard12638 = early_reset_static_par0_go_out;
wire _guard12639 = early_reset_static_par0_go_out;
wire _guard12640 = fsm0_out == 6'd0;
wire _guard12641 = early_reset_static_seq_go_out;
wire _guard12642 = _guard12640 & _guard12641;
wire _guard12643 = early_reset_static_par0_go_out;
wire _guard12644 = _guard12642 | _guard12643;
wire _guard12645 = fsm0_out == 6'd0;
wire _guard12646 = early_reset_static_seq_go_out;
wire _guard12647 = _guard12645 & _guard12646;
wire _guard12648 = early_reset_static_par0_go_out;
wire _guard12649 = early_reset_static_par0_go_out;
wire _guard12650 = early_reset_static_par0_go_out;
wire _guard12651 = early_reset_static_par0_go_out;
wire _guard12652 = early_reset_static_par0_go_out;
wire _guard12653 = early_reset_static_par0_go_out;
wire _guard12654 = early_reset_static_par0_go_out;
wire _guard12655 = early_reset_static_par0_go_out;
wire _guard12656 = early_reset_static_par0_go_out;
wire _guard12657 = early_reset_static_par0_go_out;
wire _guard12658 = early_reset_static_par0_go_out;
wire _guard12659 = early_reset_static_par0_go_out;
wire _guard12660 = early_reset_static_par0_go_out;
wire _guard12661 = early_reset_static_par0_go_out;
wire _guard12662 = early_reset_static_par0_go_out;
wire _guard12663 = early_reset_static_par0_go_out;
wire _guard12664 = early_reset_static_par0_go_out;
wire _guard12665 = early_reset_static_par0_go_out;
wire _guard12666 = early_reset_static_par0_go_out;
wire _guard12667 = early_reset_static_par0_go_out;
wire _guard12668 = early_reset_static_par0_go_out;
wire _guard12669 = early_reset_static_par0_go_out;
wire _guard12670 = early_reset_static_par0_go_out;
wire _guard12671 = early_reset_static_par0_go_out;
wire _guard12672 = early_reset_static_par0_go_out;
wire _guard12673 = early_reset_static_par0_go_out;
wire _guard12674 = ~_guard0;
wire _guard12675 = early_reset_static_par0_go_out;
wire _guard12676 = _guard12674 & _guard12675;
wire _guard12677 = early_reset_static_par0_go_out;
wire _guard12678 = early_reset_static_par0_go_out;
wire _guard12679 = early_reset_static_par0_go_out;
wire _guard12680 = early_reset_static_par0_go_out;
wire _guard12681 = early_reset_static_par0_go_out;
wire _guard12682 = early_reset_static_par0_go_out;
wire _guard12683 = early_reset_static_par0_go_out;
wire _guard12684 = ~_guard0;
wire _guard12685 = early_reset_static_par0_go_out;
wire _guard12686 = _guard12684 & _guard12685;
wire _guard12687 = early_reset_static_par0_go_out;
wire _guard12688 = early_reset_static_par0_go_out;
wire _guard12689 = early_reset_static_par0_go_out;
wire _guard12690 = early_reset_static_par0_go_out;
wire _guard12691 = early_reset_static_par0_go_out;
wire _guard12692 = early_reset_static_par0_go_out;
wire _guard12693 = early_reset_static_par0_go_out;
wire _guard12694 = early_reset_static_par0_go_out;
wire _guard12695 = early_reset_static_par0_go_out;
wire _guard12696 = ~_guard0;
wire _guard12697 = early_reset_static_par0_go_out;
wire _guard12698 = _guard12696 & _guard12697;
wire _guard12699 = early_reset_static_par0_go_out;
wire _guard12700 = ~_guard0;
wire _guard12701 = early_reset_static_par0_go_out;
wire _guard12702 = _guard12700 & _guard12701;
wire _guard12703 = ~_guard0;
wire _guard12704 = early_reset_static_par0_go_out;
wire _guard12705 = _guard12703 & _guard12704;
wire _guard12706 = early_reset_static_par0_go_out;
wire _guard12707 = early_reset_static_par0_go_out;
wire _guard12708 = ~_guard0;
wire _guard12709 = early_reset_static_par0_go_out;
wire _guard12710 = _guard12708 & _guard12709;
wire _guard12711 = early_reset_static_par0_go_out;
wire _guard12712 = ~_guard0;
wire _guard12713 = early_reset_static_par0_go_out;
wire _guard12714 = _guard12712 & _guard12713;
wire _guard12715 = early_reset_static_par0_go_out;
wire _guard12716 = ~_guard0;
wire _guard12717 = early_reset_static_par0_go_out;
wire _guard12718 = _guard12716 & _guard12717;
wire _guard12719 = early_reset_static_par0_go_out;
wire _guard12720 = ~_guard0;
wire _guard12721 = early_reset_static_par0_go_out;
wire _guard12722 = _guard12720 & _guard12721;
wire _guard12723 = early_reset_static_par0_go_out;
wire _guard12724 = early_reset_static_par0_go_out;
wire _guard12725 = ~_guard0;
wire _guard12726 = early_reset_static_par0_go_out;
wire _guard12727 = _guard12725 & _guard12726;
wire _guard12728 = early_reset_static_par0_go_out;
wire _guard12729 = early_reset_static_par0_go_out;
wire _guard12730 = early_reset_static_par0_go_out;
wire _guard12731 = early_reset_static_par0_go_out;
wire _guard12732 = early_reset_static_par0_go_out;
wire _guard12733 = early_reset_static_par0_go_out;
wire _guard12734 = early_reset_static_par0_go_out;
wire _guard12735 = early_reset_static_par0_go_out;
wire _guard12736 = early_reset_static_par0_go_out;
wire _guard12737 = early_reset_static_par0_go_out;
wire _guard12738 = early_reset_static_par0_go_out;
wire _guard12739 = early_reset_static_par0_go_out;
wire _guard12740 = early_reset_static_par0_go_out;
wire _guard12741 = early_reset_static_par0_go_out;
wire _guard12742 = early_reset_static_par0_go_out;
wire _guard12743 = early_reset_static_par0_go_out;
wire _guard12744 = ~_guard0;
wire _guard12745 = early_reset_static_par0_go_out;
wire _guard12746 = _guard12744 & _guard12745;
wire _guard12747 = early_reset_static_par0_go_out;
wire _guard12748 = ~_guard0;
wire _guard12749 = early_reset_static_par0_go_out;
wire _guard12750 = _guard12748 & _guard12749;
wire _guard12751 = ~_guard0;
wire _guard12752 = early_reset_static_par0_go_out;
wire _guard12753 = _guard12751 & _guard12752;
wire _guard12754 = early_reset_static_par0_go_out;
wire _guard12755 = early_reset_static_par0_go_out;
wire _guard12756 = early_reset_static_par0_go_out;
wire _guard12757 = early_reset_static_par0_go_out;
wire _guard12758 = ~_guard0;
wire _guard12759 = early_reset_static_par0_go_out;
wire _guard12760 = _guard12758 & _guard12759;
wire _guard12761 = early_reset_static_par0_go_out;
wire _guard12762 = early_reset_static_par0_go_out;
wire _guard12763 = ~_guard0;
wire _guard12764 = early_reset_static_par0_go_out;
wire _guard12765 = _guard12763 & _guard12764;
wire _guard12766 = early_reset_static_par0_go_out;
wire _guard12767 = early_reset_static_par0_go_out;
wire _guard12768 = early_reset_static_par0_go_out;
wire _guard12769 = early_reset_static_par0_go_out;
wire _guard12770 = early_reset_static_par0_go_out;
wire _guard12771 = early_reset_static_par0_go_out;
wire _guard12772 = early_reset_static_par0_go_out;
wire _guard12773 = early_reset_static_par0_go_out;
wire _guard12774 = ~_guard0;
wire _guard12775 = early_reset_static_par0_go_out;
wire _guard12776 = _guard12774 & _guard12775;
wire _guard12777 = early_reset_static_par0_go_out;
wire _guard12778 = early_reset_static_par0_go_out;
wire _guard12779 = early_reset_static_par0_go_out;
wire _guard12780 = early_reset_static_par0_go_out;
wire _guard12781 = early_reset_static_par0_go_out;
wire _guard12782 = early_reset_static_par0_go_out;
wire _guard12783 = early_reset_static_par0_go_out;
wire _guard12784 = early_reset_static_par0_go_out;
wire _guard12785 = early_reset_static_par0_go_out;
wire _guard12786 = early_reset_static_par0_go_out;
wire _guard12787 = early_reset_static_par0_go_out;
wire _guard12788 = early_reset_static_par0_go_out;
wire _guard12789 = early_reset_static_par0_go_out;
wire _guard12790 = early_reset_static_par0_go_out;
wire _guard12791 = ~_guard0;
wire _guard12792 = early_reset_static_par0_go_out;
wire _guard12793 = _guard12791 & _guard12792;
wire _guard12794 = early_reset_static_par0_go_out;
wire _guard12795 = early_reset_static_par0_go_out;
wire _guard12796 = early_reset_static_par0_go_out;
wire _guard12797 = early_reset_static_par0_go_out;
wire _guard12798 = early_reset_static_par0_go_out;
wire _guard12799 = early_reset_static_par0_go_out;
wire _guard12800 = early_reset_static_par0_go_out;
wire _guard12801 = early_reset_static_par0_go_out;
wire _guard12802 = early_reset_static_par0_go_out;
wire _guard12803 = ~_guard0;
wire _guard12804 = early_reset_static_par0_go_out;
wire _guard12805 = _guard12803 & _guard12804;
wire _guard12806 = early_reset_static_par0_go_out;
wire _guard12807 = early_reset_static_par0_go_out;
wire _guard12808 = ~_guard0;
wire _guard12809 = early_reset_static_par0_go_out;
wire _guard12810 = _guard12808 & _guard12809;
wire _guard12811 = ~_guard0;
wire _guard12812 = early_reset_static_par0_go_out;
wire _guard12813 = _guard12811 & _guard12812;
wire _guard12814 = early_reset_static_par0_go_out;
wire _guard12815 = ~_guard0;
wire _guard12816 = early_reset_static_par0_go_out;
wire _guard12817 = _guard12815 & _guard12816;
wire _guard12818 = early_reset_static_par0_go_out;
wire _guard12819 = ~_guard0;
wire _guard12820 = early_reset_static_par0_go_out;
wire _guard12821 = _guard12819 & _guard12820;
wire _guard12822 = early_reset_static_par0_go_out;
wire _guard12823 = early_reset_static_par0_go_out;
wire _guard12824 = ~_guard0;
wire _guard12825 = early_reset_static_par0_go_out;
wire _guard12826 = _guard12824 & _guard12825;
wire _guard12827 = early_reset_static_par0_go_out;
wire _guard12828 = ~_guard0;
wire _guard12829 = early_reset_static_par0_go_out;
wire _guard12830 = _guard12828 & _guard12829;
wire _guard12831 = early_reset_static_par0_go_out;
wire _guard12832 = early_reset_static_par0_go_out;
wire _guard12833 = early_reset_static_par0_go_out;
wire _guard12834 = ~_guard0;
wire _guard12835 = early_reset_static_par0_go_out;
wire _guard12836 = _guard12834 & _guard12835;
wire _guard12837 = early_reset_static_par0_go_out;
wire _guard12838 = early_reset_static_par0_go_out;
wire _guard12839 = early_reset_static_par0_go_out;
wire _guard12840 = ~_guard0;
wire _guard12841 = early_reset_static_par0_go_out;
wire _guard12842 = _guard12840 & _guard12841;
wire _guard12843 = early_reset_static_par0_go_out;
wire _guard12844 = early_reset_static_par0_go_out;
wire _guard12845 = early_reset_static_par0_go_out;
wire _guard12846 = ~_guard0;
wire _guard12847 = early_reset_static_par0_go_out;
wire _guard12848 = _guard12846 & _guard12847;
wire _guard12849 = early_reset_static_par0_go_out;
wire _guard12850 = ~_guard0;
wire _guard12851 = early_reset_static_par0_go_out;
wire _guard12852 = _guard12850 & _guard12851;
wire _guard12853 = early_reset_static_par0_go_out;
wire _guard12854 = early_reset_static_par0_go_out;
wire _guard12855 = early_reset_static_par0_go_out;
wire _guard12856 = ~_guard0;
wire _guard12857 = early_reset_static_par0_go_out;
wire _guard12858 = _guard12856 & _guard12857;
wire _guard12859 = early_reset_static_par0_go_out;
wire _guard12860 = ~_guard0;
wire _guard12861 = early_reset_static_par0_go_out;
wire _guard12862 = _guard12860 & _guard12861;
wire _guard12863 = early_reset_static_par0_go_out;
wire _guard12864 = early_reset_static_par0_go_out;
wire _guard12865 = early_reset_static_par0_go_out;
wire _guard12866 = early_reset_static_par0_go_out;
wire _guard12867 = ~_guard0;
wire _guard12868 = early_reset_static_par0_go_out;
wire _guard12869 = _guard12867 & _guard12868;
wire _guard12870 = early_reset_static_par0_go_out;
wire _guard12871 = early_reset_static_par0_go_out;
wire _guard12872 = early_reset_static_par0_go_out;
wire _guard12873 = early_reset_static_par0_go_out;
wire _guard12874 = early_reset_static_par0_go_out;
wire _guard12875 = early_reset_static_par0_go_out;
wire _guard12876 = early_reset_static_par0_go_out;
wire _guard12877 = early_reset_static_par0_go_out;
wire _guard12878 = ~_guard0;
wire _guard12879 = early_reset_static_par0_go_out;
wire _guard12880 = _guard12878 & _guard12879;
wire _guard12881 = early_reset_static_par0_go_out;
wire _guard12882 = early_reset_static_par0_go_out;
wire _guard12883 = ~_guard0;
wire _guard12884 = early_reset_static_par0_go_out;
wire _guard12885 = _guard12883 & _guard12884;
wire _guard12886 = early_reset_static_par0_go_out;
wire _guard12887 = early_reset_static_par0_go_out;
wire _guard12888 = early_reset_static_par0_go_out;
wire _guard12889 = early_reset_static_par0_go_out;
wire _guard12890 = early_reset_static_par0_go_out;
wire _guard12891 = early_reset_static_par0_go_out;
wire _guard12892 = early_reset_static_par0_go_out;
wire _guard12893 = early_reset_static_par0_go_out;
wire _guard12894 = early_reset_static_par0_go_out;
wire _guard12895 = early_reset_static_par0_go_out;
wire _guard12896 = ~_guard0;
wire _guard12897 = early_reset_static_par0_go_out;
wire _guard12898 = _guard12896 & _guard12897;
wire _guard12899 = early_reset_static_par0_go_out;
wire _guard12900 = early_reset_static_par0_go_out;
wire _guard12901 = early_reset_static_par0_go_out;
wire _guard12902 = early_reset_static_par0_go_out;
wire _guard12903 = early_reset_static_par0_go_out;
wire _guard12904 = ~_guard0;
wire _guard12905 = early_reset_static_par0_go_out;
wire _guard12906 = _guard12904 & _guard12905;
wire _guard12907 = early_reset_static_par0_go_out;
wire _guard12908 = early_reset_static_par0_go_out;
wire _guard12909 = early_reset_static_par0_go_out;
wire _guard12910 = ~_guard0;
wire _guard12911 = early_reset_static_par0_go_out;
wire _guard12912 = _guard12910 & _guard12911;
wire _guard12913 = early_reset_static_par0_go_out;
wire _guard12914 = early_reset_static_par0_go_out;
wire _guard12915 = early_reset_static_par0_go_out;
wire _guard12916 = early_reset_static_par0_go_out;
wire _guard12917 = ~_guard0;
wire _guard12918 = early_reset_static_par0_go_out;
wire _guard12919 = _guard12917 & _guard12918;
wire _guard12920 = early_reset_static_par0_go_out;
wire _guard12921 = early_reset_static_par0_go_out;
wire _guard12922 = early_reset_static_par0_go_out;
wire _guard12923 = early_reset_static_par0_go_out;
wire _guard12924 = early_reset_static_par0_go_out;
wire _guard12925 = early_reset_static_par0_go_out;
wire _guard12926 = early_reset_static_par0_go_out;
wire _guard12927 = early_reset_static_par0_go_out;
wire _guard12928 = early_reset_static_par0_go_out;
wire _guard12929 = ~_guard0;
wire _guard12930 = early_reset_static_par0_go_out;
wire _guard12931 = _guard12929 & _guard12930;
wire _guard12932 = early_reset_static_par0_go_out;
wire _guard12933 = early_reset_static_par0_go_out;
wire _guard12934 = early_reset_static_par0_go_out;
wire _guard12935 = early_reset_static_par0_go_out;
wire _guard12936 = ~_guard0;
wire _guard12937 = early_reset_static_par0_go_out;
wire _guard12938 = _guard12936 & _guard12937;
wire _guard12939 = early_reset_static_par0_go_out;
wire _guard12940 = early_reset_static_par0_go_out;
wire _guard12941 = ~_guard0;
wire _guard12942 = early_reset_static_par0_go_out;
wire _guard12943 = _guard12941 & _guard12942;
wire _guard12944 = early_reset_static_par0_go_out;
wire _guard12945 = early_reset_static_par0_go_out;
wire _guard12946 = early_reset_static_par0_go_out;
wire _guard12947 = ~_guard0;
wire _guard12948 = early_reset_static_par0_go_out;
wire _guard12949 = _guard12947 & _guard12948;
wire _guard12950 = early_reset_static_par0_go_out;
wire _guard12951 = early_reset_static_par0_go_out;
wire _guard12952 = early_reset_static_par0_go_out;
wire _guard12953 = early_reset_static_par0_go_out;
wire _guard12954 = ~_guard0;
wire _guard12955 = early_reset_static_par0_go_out;
wire _guard12956 = _guard12954 & _guard12955;
wire _guard12957 = early_reset_static_par0_go_out;
wire _guard12958 = early_reset_static_par0_go_out;
wire _guard12959 = early_reset_static_par0_go_out;
wire _guard12960 = early_reset_static_par0_go_out;
wire _guard12961 = early_reset_static_par0_go_out;
wire _guard12962 = early_reset_static_par0_go_out;
wire _guard12963 = early_reset_static_par0_go_out;
wire _guard12964 = ~_guard0;
wire _guard12965 = early_reset_static_par0_go_out;
wire _guard12966 = _guard12964 & _guard12965;
wire _guard12967 = early_reset_static_par0_go_out;
wire _guard12968 = early_reset_static_par0_go_out;
wire _guard12969 = early_reset_static_par0_go_out;
wire _guard12970 = early_reset_static_par0_go_out;
wire _guard12971 = early_reset_static_par0_go_out;
wire _guard12972 = ~_guard0;
wire _guard12973 = early_reset_static_par0_go_out;
wire _guard12974 = _guard12972 & _guard12973;
wire _guard12975 = early_reset_static_par0_go_out;
wire _guard12976 = early_reset_static_par0_go_out;
wire _guard12977 = early_reset_static_par0_go_out;
wire _guard12978 = early_reset_static_par0_go_out;
wire _guard12979 = early_reset_static_par0_go_out;
wire _guard12980 = early_reset_static_par0_go_out;
wire _guard12981 = early_reset_static_par0_go_out;
wire _guard12982 = early_reset_static_par0_go_out;
wire _guard12983 = early_reset_static_par0_go_out;
wire _guard12984 = ~_guard0;
wire _guard12985 = early_reset_static_par0_go_out;
wire _guard12986 = _guard12984 & _guard12985;
wire _guard12987 = early_reset_static_par0_go_out;
wire _guard12988 = early_reset_static_par0_go_out;
wire _guard12989 = ~_guard0;
wire _guard12990 = early_reset_static_par0_go_out;
wire _guard12991 = _guard12989 & _guard12990;
wire _guard12992 = early_reset_static_par0_go_out;
wire _guard12993 = early_reset_static_par0_go_out;
wire _guard12994 = ~_guard0;
wire _guard12995 = early_reset_static_par0_go_out;
wire _guard12996 = _guard12994 & _guard12995;
wire _guard12997 = ~_guard0;
wire _guard12998 = early_reset_static_par0_go_out;
wire _guard12999 = _guard12997 & _guard12998;
wire _guard13000 = early_reset_static_par0_go_out;
wire _guard13001 = early_reset_static_par0_go_out;
wire _guard13002 = early_reset_static_par0_go_out;
wire _guard13003 = ~_guard0;
wire _guard13004 = early_reset_static_par0_go_out;
wire _guard13005 = _guard13003 & _guard13004;
wire _guard13006 = early_reset_static_par0_go_out;
wire _guard13007 = cond_wire31_out;
wire _guard13008 = early_reset_static_par0_go_out;
wire _guard13009 = _guard13007 & _guard13008;
wire _guard13010 = cond_wire31_out;
wire _guard13011 = early_reset_static_par0_go_out;
wire _guard13012 = _guard13010 & _guard13011;
wire _guard13013 = cond_wire69_out;
wire _guard13014 = early_reset_static_par0_go_out;
wire _guard13015 = _guard13013 & _guard13014;
wire _guard13016 = cond_wire69_out;
wire _guard13017 = early_reset_static_par0_go_out;
wire _guard13018 = _guard13016 & _guard13017;
wire _guard13019 = cond_wire130_out;
wire _guard13020 = early_reset_static_par0_go_out;
wire _guard13021 = _guard13019 & _guard13020;
wire _guard13022 = cond_wire128_out;
wire _guard13023 = early_reset_static_par0_go_out;
wire _guard13024 = _guard13022 & _guard13023;
wire _guard13025 = fsm_out == 1'd0;
wire _guard13026 = cond_wire128_out;
wire _guard13027 = _guard13025 & _guard13026;
wire _guard13028 = fsm_out == 1'd0;
wire _guard13029 = _guard13027 & _guard13028;
wire _guard13030 = fsm_out == 1'd0;
wire _guard13031 = cond_wire130_out;
wire _guard13032 = _guard13030 & _guard13031;
wire _guard13033 = fsm_out == 1'd0;
wire _guard13034 = _guard13032 & _guard13033;
wire _guard13035 = _guard13029 | _guard13034;
wire _guard13036 = early_reset_static_par0_go_out;
wire _guard13037 = _guard13035 & _guard13036;
wire _guard13038 = fsm_out == 1'd0;
wire _guard13039 = cond_wire128_out;
wire _guard13040 = _guard13038 & _guard13039;
wire _guard13041 = fsm_out == 1'd0;
wire _guard13042 = _guard13040 & _guard13041;
wire _guard13043 = fsm_out == 1'd0;
wire _guard13044 = cond_wire130_out;
wire _guard13045 = _guard13043 & _guard13044;
wire _guard13046 = fsm_out == 1'd0;
wire _guard13047 = _guard13045 & _guard13046;
wire _guard13048 = _guard13042 | _guard13047;
wire _guard13049 = early_reset_static_par0_go_out;
wire _guard13050 = _guard13048 & _guard13049;
wire _guard13051 = fsm_out == 1'd0;
wire _guard13052 = cond_wire128_out;
wire _guard13053 = _guard13051 & _guard13052;
wire _guard13054 = fsm_out == 1'd0;
wire _guard13055 = _guard13053 & _guard13054;
wire _guard13056 = fsm_out == 1'd0;
wire _guard13057 = cond_wire130_out;
wire _guard13058 = _guard13056 & _guard13057;
wire _guard13059 = fsm_out == 1'd0;
wire _guard13060 = _guard13058 & _guard13059;
wire _guard13061 = _guard13055 | _guard13060;
wire _guard13062 = early_reset_static_par0_go_out;
wire _guard13063 = _guard13061 & _guard13062;
wire _guard13064 = cond_wire151_out;
wire _guard13065 = early_reset_static_par0_go_out;
wire _guard13066 = _guard13064 & _guard13065;
wire _guard13067 = cond_wire149_out;
wire _guard13068 = early_reset_static_par0_go_out;
wire _guard13069 = _guard13067 & _guard13068;
wire _guard13070 = fsm_out == 1'd0;
wire _guard13071 = cond_wire149_out;
wire _guard13072 = _guard13070 & _guard13071;
wire _guard13073 = fsm_out == 1'd0;
wire _guard13074 = _guard13072 & _guard13073;
wire _guard13075 = fsm_out == 1'd0;
wire _guard13076 = cond_wire151_out;
wire _guard13077 = _guard13075 & _guard13076;
wire _guard13078 = fsm_out == 1'd0;
wire _guard13079 = _guard13077 & _guard13078;
wire _guard13080 = _guard13074 | _guard13079;
wire _guard13081 = early_reset_static_par0_go_out;
wire _guard13082 = _guard13080 & _guard13081;
wire _guard13083 = fsm_out == 1'd0;
wire _guard13084 = cond_wire149_out;
wire _guard13085 = _guard13083 & _guard13084;
wire _guard13086 = fsm_out == 1'd0;
wire _guard13087 = _guard13085 & _guard13086;
wire _guard13088 = fsm_out == 1'd0;
wire _guard13089 = cond_wire151_out;
wire _guard13090 = _guard13088 & _guard13089;
wire _guard13091 = fsm_out == 1'd0;
wire _guard13092 = _guard13090 & _guard13091;
wire _guard13093 = _guard13087 | _guard13092;
wire _guard13094 = early_reset_static_par0_go_out;
wire _guard13095 = _guard13093 & _guard13094;
wire _guard13096 = fsm_out == 1'd0;
wire _guard13097 = cond_wire149_out;
wire _guard13098 = _guard13096 & _guard13097;
wire _guard13099 = fsm_out == 1'd0;
wire _guard13100 = _guard13098 & _guard13099;
wire _guard13101 = fsm_out == 1'd0;
wire _guard13102 = cond_wire151_out;
wire _guard13103 = _guard13101 & _guard13102;
wire _guard13104 = fsm_out == 1'd0;
wire _guard13105 = _guard13103 & _guard13104;
wire _guard13106 = _guard13100 | _guard13105;
wire _guard13107 = early_reset_static_par0_go_out;
wire _guard13108 = _guard13106 & _guard13107;
wire _guard13109 = cond_wire159_out;
wire _guard13110 = early_reset_static_par0_go_out;
wire _guard13111 = _guard13109 & _guard13110;
wire _guard13112 = cond_wire157_out;
wire _guard13113 = early_reset_static_par0_go_out;
wire _guard13114 = _guard13112 & _guard13113;
wire _guard13115 = fsm_out == 1'd0;
wire _guard13116 = cond_wire157_out;
wire _guard13117 = _guard13115 & _guard13116;
wire _guard13118 = fsm_out == 1'd0;
wire _guard13119 = _guard13117 & _guard13118;
wire _guard13120 = fsm_out == 1'd0;
wire _guard13121 = cond_wire159_out;
wire _guard13122 = _guard13120 & _guard13121;
wire _guard13123 = fsm_out == 1'd0;
wire _guard13124 = _guard13122 & _guard13123;
wire _guard13125 = _guard13119 | _guard13124;
wire _guard13126 = early_reset_static_par0_go_out;
wire _guard13127 = _guard13125 & _guard13126;
wire _guard13128 = fsm_out == 1'd0;
wire _guard13129 = cond_wire157_out;
wire _guard13130 = _guard13128 & _guard13129;
wire _guard13131 = fsm_out == 1'd0;
wire _guard13132 = _guard13130 & _guard13131;
wire _guard13133 = fsm_out == 1'd0;
wire _guard13134 = cond_wire159_out;
wire _guard13135 = _guard13133 & _guard13134;
wire _guard13136 = fsm_out == 1'd0;
wire _guard13137 = _guard13135 & _guard13136;
wire _guard13138 = _guard13132 | _guard13137;
wire _guard13139 = early_reset_static_par0_go_out;
wire _guard13140 = _guard13138 & _guard13139;
wire _guard13141 = fsm_out == 1'd0;
wire _guard13142 = cond_wire157_out;
wire _guard13143 = _guard13141 & _guard13142;
wire _guard13144 = fsm_out == 1'd0;
wire _guard13145 = _guard13143 & _guard13144;
wire _guard13146 = fsm_out == 1'd0;
wire _guard13147 = cond_wire159_out;
wire _guard13148 = _guard13146 & _guard13147;
wire _guard13149 = fsm_out == 1'd0;
wire _guard13150 = _guard13148 & _guard13149;
wire _guard13151 = _guard13145 | _guard13150;
wire _guard13152 = early_reset_static_par0_go_out;
wire _guard13153 = _guard13151 & _guard13152;
wire _guard13154 = cond_wire167_out;
wire _guard13155 = early_reset_static_par0_go_out;
wire _guard13156 = _guard13154 & _guard13155;
wire _guard13157 = cond_wire165_out;
wire _guard13158 = early_reset_static_par0_go_out;
wire _guard13159 = _guard13157 & _guard13158;
wire _guard13160 = fsm_out == 1'd0;
wire _guard13161 = cond_wire165_out;
wire _guard13162 = _guard13160 & _guard13161;
wire _guard13163 = fsm_out == 1'd0;
wire _guard13164 = _guard13162 & _guard13163;
wire _guard13165 = fsm_out == 1'd0;
wire _guard13166 = cond_wire167_out;
wire _guard13167 = _guard13165 & _guard13166;
wire _guard13168 = fsm_out == 1'd0;
wire _guard13169 = _guard13167 & _guard13168;
wire _guard13170 = _guard13164 | _guard13169;
wire _guard13171 = early_reset_static_par0_go_out;
wire _guard13172 = _guard13170 & _guard13171;
wire _guard13173 = fsm_out == 1'd0;
wire _guard13174 = cond_wire165_out;
wire _guard13175 = _guard13173 & _guard13174;
wire _guard13176 = fsm_out == 1'd0;
wire _guard13177 = _guard13175 & _guard13176;
wire _guard13178 = fsm_out == 1'd0;
wire _guard13179 = cond_wire167_out;
wire _guard13180 = _guard13178 & _guard13179;
wire _guard13181 = fsm_out == 1'd0;
wire _guard13182 = _guard13180 & _guard13181;
wire _guard13183 = _guard13177 | _guard13182;
wire _guard13184 = early_reset_static_par0_go_out;
wire _guard13185 = _guard13183 & _guard13184;
wire _guard13186 = fsm_out == 1'd0;
wire _guard13187 = cond_wire165_out;
wire _guard13188 = _guard13186 & _guard13187;
wire _guard13189 = fsm_out == 1'd0;
wire _guard13190 = _guard13188 & _guard13189;
wire _guard13191 = fsm_out == 1'd0;
wire _guard13192 = cond_wire167_out;
wire _guard13193 = _guard13191 & _guard13192;
wire _guard13194 = fsm_out == 1'd0;
wire _guard13195 = _guard13193 & _guard13194;
wire _guard13196 = _guard13190 | _guard13195;
wire _guard13197 = early_reset_static_par0_go_out;
wire _guard13198 = _guard13196 & _guard13197;
wire _guard13199 = cond_wire216_out;
wire _guard13200 = early_reset_static_par0_go_out;
wire _guard13201 = _guard13199 & _guard13200;
wire _guard13202 = cond_wire214_out;
wire _guard13203 = early_reset_static_par0_go_out;
wire _guard13204 = _guard13202 & _guard13203;
wire _guard13205 = fsm_out == 1'd0;
wire _guard13206 = cond_wire214_out;
wire _guard13207 = _guard13205 & _guard13206;
wire _guard13208 = fsm_out == 1'd0;
wire _guard13209 = _guard13207 & _guard13208;
wire _guard13210 = fsm_out == 1'd0;
wire _guard13211 = cond_wire216_out;
wire _guard13212 = _guard13210 & _guard13211;
wire _guard13213 = fsm_out == 1'd0;
wire _guard13214 = _guard13212 & _guard13213;
wire _guard13215 = _guard13209 | _guard13214;
wire _guard13216 = early_reset_static_par0_go_out;
wire _guard13217 = _guard13215 & _guard13216;
wire _guard13218 = fsm_out == 1'd0;
wire _guard13219 = cond_wire214_out;
wire _guard13220 = _guard13218 & _guard13219;
wire _guard13221 = fsm_out == 1'd0;
wire _guard13222 = _guard13220 & _guard13221;
wire _guard13223 = fsm_out == 1'd0;
wire _guard13224 = cond_wire216_out;
wire _guard13225 = _guard13223 & _guard13224;
wire _guard13226 = fsm_out == 1'd0;
wire _guard13227 = _guard13225 & _guard13226;
wire _guard13228 = _guard13222 | _guard13227;
wire _guard13229 = early_reset_static_par0_go_out;
wire _guard13230 = _guard13228 & _guard13229;
wire _guard13231 = fsm_out == 1'd0;
wire _guard13232 = cond_wire214_out;
wire _guard13233 = _guard13231 & _guard13232;
wire _guard13234 = fsm_out == 1'd0;
wire _guard13235 = _guard13233 & _guard13234;
wire _guard13236 = fsm_out == 1'd0;
wire _guard13237 = cond_wire216_out;
wire _guard13238 = _guard13236 & _guard13237;
wire _guard13239 = fsm_out == 1'd0;
wire _guard13240 = _guard13238 & _guard13239;
wire _guard13241 = _guard13235 | _guard13240;
wire _guard13242 = early_reset_static_par0_go_out;
wire _guard13243 = _guard13241 & _guard13242;
wire _guard13244 = cond_wire162_out;
wire _guard13245 = early_reset_static_par0_go_out;
wire _guard13246 = _guard13244 & _guard13245;
wire _guard13247 = cond_wire162_out;
wire _guard13248 = early_reset_static_par0_go_out;
wire _guard13249 = _guard13247 & _guard13248;
wire _guard13250 = cond_wire252_out;
wire _guard13251 = early_reset_static_par0_go_out;
wire _guard13252 = _guard13250 & _guard13251;
wire _guard13253 = cond_wire250_out;
wire _guard13254 = early_reset_static_par0_go_out;
wire _guard13255 = _guard13253 & _guard13254;
wire _guard13256 = fsm_out == 1'd0;
wire _guard13257 = cond_wire250_out;
wire _guard13258 = _guard13256 & _guard13257;
wire _guard13259 = fsm_out == 1'd0;
wire _guard13260 = _guard13258 & _guard13259;
wire _guard13261 = fsm_out == 1'd0;
wire _guard13262 = cond_wire252_out;
wire _guard13263 = _guard13261 & _guard13262;
wire _guard13264 = fsm_out == 1'd0;
wire _guard13265 = _guard13263 & _guard13264;
wire _guard13266 = _guard13260 | _guard13265;
wire _guard13267 = early_reset_static_par0_go_out;
wire _guard13268 = _guard13266 & _guard13267;
wire _guard13269 = fsm_out == 1'd0;
wire _guard13270 = cond_wire250_out;
wire _guard13271 = _guard13269 & _guard13270;
wire _guard13272 = fsm_out == 1'd0;
wire _guard13273 = _guard13271 & _guard13272;
wire _guard13274 = fsm_out == 1'd0;
wire _guard13275 = cond_wire252_out;
wire _guard13276 = _guard13274 & _guard13275;
wire _guard13277 = fsm_out == 1'd0;
wire _guard13278 = _guard13276 & _guard13277;
wire _guard13279 = _guard13273 | _guard13278;
wire _guard13280 = early_reset_static_par0_go_out;
wire _guard13281 = _guard13279 & _guard13280;
wire _guard13282 = fsm_out == 1'd0;
wire _guard13283 = cond_wire250_out;
wire _guard13284 = _guard13282 & _guard13283;
wire _guard13285 = fsm_out == 1'd0;
wire _guard13286 = _guard13284 & _guard13285;
wire _guard13287 = fsm_out == 1'd0;
wire _guard13288 = cond_wire252_out;
wire _guard13289 = _guard13287 & _guard13288;
wire _guard13290 = fsm_out == 1'd0;
wire _guard13291 = _guard13289 & _guard13290;
wire _guard13292 = _guard13286 | _guard13291;
wire _guard13293 = early_reset_static_par0_go_out;
wire _guard13294 = _guard13292 & _guard13293;
wire _guard13295 = cond_wire263_out;
wire _guard13296 = early_reset_static_par0_go_out;
wire _guard13297 = _guard13295 & _guard13296;
wire _guard13298 = cond_wire263_out;
wire _guard13299 = early_reset_static_par0_go_out;
wire _guard13300 = _guard13298 & _guard13299;
wire _guard13301 = cond_wire333_out;
wire _guard13302 = early_reset_static_par0_go_out;
wire _guard13303 = _guard13301 & _guard13302;
wire _guard13304 = cond_wire331_out;
wire _guard13305 = early_reset_static_par0_go_out;
wire _guard13306 = _guard13304 & _guard13305;
wire _guard13307 = fsm_out == 1'd0;
wire _guard13308 = cond_wire331_out;
wire _guard13309 = _guard13307 & _guard13308;
wire _guard13310 = fsm_out == 1'd0;
wire _guard13311 = _guard13309 & _guard13310;
wire _guard13312 = fsm_out == 1'd0;
wire _guard13313 = cond_wire333_out;
wire _guard13314 = _guard13312 & _guard13313;
wire _guard13315 = fsm_out == 1'd0;
wire _guard13316 = _guard13314 & _guard13315;
wire _guard13317 = _guard13311 | _guard13316;
wire _guard13318 = early_reset_static_par0_go_out;
wire _guard13319 = _guard13317 & _guard13318;
wire _guard13320 = fsm_out == 1'd0;
wire _guard13321 = cond_wire331_out;
wire _guard13322 = _guard13320 & _guard13321;
wire _guard13323 = fsm_out == 1'd0;
wire _guard13324 = _guard13322 & _guard13323;
wire _guard13325 = fsm_out == 1'd0;
wire _guard13326 = cond_wire333_out;
wire _guard13327 = _guard13325 & _guard13326;
wire _guard13328 = fsm_out == 1'd0;
wire _guard13329 = _guard13327 & _guard13328;
wire _guard13330 = _guard13324 | _guard13329;
wire _guard13331 = early_reset_static_par0_go_out;
wire _guard13332 = _guard13330 & _guard13331;
wire _guard13333 = fsm_out == 1'd0;
wire _guard13334 = cond_wire331_out;
wire _guard13335 = _guard13333 & _guard13334;
wire _guard13336 = fsm_out == 1'd0;
wire _guard13337 = _guard13335 & _guard13336;
wire _guard13338 = fsm_out == 1'd0;
wire _guard13339 = cond_wire333_out;
wire _guard13340 = _guard13338 & _guard13339;
wire _guard13341 = fsm_out == 1'd0;
wire _guard13342 = _guard13340 & _guard13341;
wire _guard13343 = _guard13337 | _guard13342;
wire _guard13344 = early_reset_static_par0_go_out;
wire _guard13345 = _guard13343 & _guard13344;
wire _guard13346 = cond_wire337_out;
wire _guard13347 = early_reset_static_par0_go_out;
wire _guard13348 = _guard13346 & _guard13347;
wire _guard13349 = cond_wire335_out;
wire _guard13350 = early_reset_static_par0_go_out;
wire _guard13351 = _guard13349 & _guard13350;
wire _guard13352 = fsm_out == 1'd0;
wire _guard13353 = cond_wire335_out;
wire _guard13354 = _guard13352 & _guard13353;
wire _guard13355 = fsm_out == 1'd0;
wire _guard13356 = _guard13354 & _guard13355;
wire _guard13357 = fsm_out == 1'd0;
wire _guard13358 = cond_wire337_out;
wire _guard13359 = _guard13357 & _guard13358;
wire _guard13360 = fsm_out == 1'd0;
wire _guard13361 = _guard13359 & _guard13360;
wire _guard13362 = _guard13356 | _guard13361;
wire _guard13363 = early_reset_static_par0_go_out;
wire _guard13364 = _guard13362 & _guard13363;
wire _guard13365 = fsm_out == 1'd0;
wire _guard13366 = cond_wire335_out;
wire _guard13367 = _guard13365 & _guard13366;
wire _guard13368 = fsm_out == 1'd0;
wire _guard13369 = _guard13367 & _guard13368;
wire _guard13370 = fsm_out == 1'd0;
wire _guard13371 = cond_wire337_out;
wire _guard13372 = _guard13370 & _guard13371;
wire _guard13373 = fsm_out == 1'd0;
wire _guard13374 = _guard13372 & _guard13373;
wire _guard13375 = _guard13369 | _guard13374;
wire _guard13376 = early_reset_static_par0_go_out;
wire _guard13377 = _guard13375 & _guard13376;
wire _guard13378 = fsm_out == 1'd0;
wire _guard13379 = cond_wire335_out;
wire _guard13380 = _guard13378 & _guard13379;
wire _guard13381 = fsm_out == 1'd0;
wire _guard13382 = _guard13380 & _guard13381;
wire _guard13383 = fsm_out == 1'd0;
wire _guard13384 = cond_wire337_out;
wire _guard13385 = _guard13383 & _guard13384;
wire _guard13386 = fsm_out == 1'd0;
wire _guard13387 = _guard13385 & _guard13386;
wire _guard13388 = _guard13382 | _guard13387;
wire _guard13389 = early_reset_static_par0_go_out;
wire _guard13390 = _guard13388 & _guard13389;
wire _guard13391 = cond_wire354_out;
wire _guard13392 = early_reset_static_par0_go_out;
wire _guard13393 = _guard13391 & _guard13392;
wire _guard13394 = cond_wire352_out;
wire _guard13395 = early_reset_static_par0_go_out;
wire _guard13396 = _guard13394 & _guard13395;
wire _guard13397 = fsm_out == 1'd0;
wire _guard13398 = cond_wire352_out;
wire _guard13399 = _guard13397 & _guard13398;
wire _guard13400 = fsm_out == 1'd0;
wire _guard13401 = _guard13399 & _guard13400;
wire _guard13402 = fsm_out == 1'd0;
wire _guard13403 = cond_wire354_out;
wire _guard13404 = _guard13402 & _guard13403;
wire _guard13405 = fsm_out == 1'd0;
wire _guard13406 = _guard13404 & _guard13405;
wire _guard13407 = _guard13401 | _guard13406;
wire _guard13408 = early_reset_static_par0_go_out;
wire _guard13409 = _guard13407 & _guard13408;
wire _guard13410 = fsm_out == 1'd0;
wire _guard13411 = cond_wire352_out;
wire _guard13412 = _guard13410 & _guard13411;
wire _guard13413 = fsm_out == 1'd0;
wire _guard13414 = _guard13412 & _guard13413;
wire _guard13415 = fsm_out == 1'd0;
wire _guard13416 = cond_wire354_out;
wire _guard13417 = _guard13415 & _guard13416;
wire _guard13418 = fsm_out == 1'd0;
wire _guard13419 = _guard13417 & _guard13418;
wire _guard13420 = _guard13414 | _guard13419;
wire _guard13421 = early_reset_static_par0_go_out;
wire _guard13422 = _guard13420 & _guard13421;
wire _guard13423 = fsm_out == 1'd0;
wire _guard13424 = cond_wire352_out;
wire _guard13425 = _guard13423 & _guard13424;
wire _guard13426 = fsm_out == 1'd0;
wire _guard13427 = _guard13425 & _guard13426;
wire _guard13428 = fsm_out == 1'd0;
wire _guard13429 = cond_wire354_out;
wire _guard13430 = _guard13428 & _guard13429;
wire _guard13431 = fsm_out == 1'd0;
wire _guard13432 = _guard13430 & _guard13431;
wire _guard13433 = _guard13427 | _guard13432;
wire _guard13434 = early_reset_static_par0_go_out;
wire _guard13435 = _guard13433 & _guard13434;
wire _guard13436 = cond_wire362_out;
wire _guard13437 = early_reset_static_par0_go_out;
wire _guard13438 = _guard13436 & _guard13437;
wire _guard13439 = cond_wire360_out;
wire _guard13440 = early_reset_static_par0_go_out;
wire _guard13441 = _guard13439 & _guard13440;
wire _guard13442 = fsm_out == 1'd0;
wire _guard13443 = cond_wire360_out;
wire _guard13444 = _guard13442 & _guard13443;
wire _guard13445 = fsm_out == 1'd0;
wire _guard13446 = _guard13444 & _guard13445;
wire _guard13447 = fsm_out == 1'd0;
wire _guard13448 = cond_wire362_out;
wire _guard13449 = _guard13447 & _guard13448;
wire _guard13450 = fsm_out == 1'd0;
wire _guard13451 = _guard13449 & _guard13450;
wire _guard13452 = _guard13446 | _guard13451;
wire _guard13453 = early_reset_static_par0_go_out;
wire _guard13454 = _guard13452 & _guard13453;
wire _guard13455 = fsm_out == 1'd0;
wire _guard13456 = cond_wire360_out;
wire _guard13457 = _guard13455 & _guard13456;
wire _guard13458 = fsm_out == 1'd0;
wire _guard13459 = _guard13457 & _guard13458;
wire _guard13460 = fsm_out == 1'd0;
wire _guard13461 = cond_wire362_out;
wire _guard13462 = _guard13460 & _guard13461;
wire _guard13463 = fsm_out == 1'd0;
wire _guard13464 = _guard13462 & _guard13463;
wire _guard13465 = _guard13459 | _guard13464;
wire _guard13466 = early_reset_static_par0_go_out;
wire _guard13467 = _guard13465 & _guard13466;
wire _guard13468 = fsm_out == 1'd0;
wire _guard13469 = cond_wire360_out;
wire _guard13470 = _guard13468 & _guard13469;
wire _guard13471 = fsm_out == 1'd0;
wire _guard13472 = _guard13470 & _guard13471;
wire _guard13473 = fsm_out == 1'd0;
wire _guard13474 = cond_wire362_out;
wire _guard13475 = _guard13473 & _guard13474;
wire _guard13476 = fsm_out == 1'd0;
wire _guard13477 = _guard13475 & _guard13476;
wire _guard13478 = _guard13472 | _guard13477;
wire _guard13479 = early_reset_static_par0_go_out;
wire _guard13480 = _guard13478 & _guard13479;
wire _guard13481 = cond_wire369_out;
wire _guard13482 = early_reset_static_par0_go_out;
wire _guard13483 = _guard13481 & _guard13482;
wire _guard13484 = cond_wire369_out;
wire _guard13485 = early_reset_static_par0_go_out;
wire _guard13486 = _guard13484 & _guard13485;
wire _guard13487 = cond_wire389_out;
wire _guard13488 = early_reset_static_par0_go_out;
wire _guard13489 = _guard13487 & _guard13488;
wire _guard13490 = cond_wire389_out;
wire _guard13491 = early_reset_static_par0_go_out;
wire _guard13492 = _guard13490 & _guard13491;
wire _guard13493 = cond_wire415_out;
wire _guard13494 = early_reset_static_par0_go_out;
wire _guard13495 = _guard13493 & _guard13494;
wire _guard13496 = cond_wire413_out;
wire _guard13497 = early_reset_static_par0_go_out;
wire _guard13498 = _guard13496 & _guard13497;
wire _guard13499 = fsm_out == 1'd0;
wire _guard13500 = cond_wire413_out;
wire _guard13501 = _guard13499 & _guard13500;
wire _guard13502 = fsm_out == 1'd0;
wire _guard13503 = _guard13501 & _guard13502;
wire _guard13504 = fsm_out == 1'd0;
wire _guard13505 = cond_wire415_out;
wire _guard13506 = _guard13504 & _guard13505;
wire _guard13507 = fsm_out == 1'd0;
wire _guard13508 = _guard13506 & _guard13507;
wire _guard13509 = _guard13503 | _guard13508;
wire _guard13510 = early_reset_static_par0_go_out;
wire _guard13511 = _guard13509 & _guard13510;
wire _guard13512 = fsm_out == 1'd0;
wire _guard13513 = cond_wire413_out;
wire _guard13514 = _guard13512 & _guard13513;
wire _guard13515 = fsm_out == 1'd0;
wire _guard13516 = _guard13514 & _guard13515;
wire _guard13517 = fsm_out == 1'd0;
wire _guard13518 = cond_wire415_out;
wire _guard13519 = _guard13517 & _guard13518;
wire _guard13520 = fsm_out == 1'd0;
wire _guard13521 = _guard13519 & _guard13520;
wire _guard13522 = _guard13516 | _guard13521;
wire _guard13523 = early_reset_static_par0_go_out;
wire _guard13524 = _guard13522 & _guard13523;
wire _guard13525 = fsm_out == 1'd0;
wire _guard13526 = cond_wire413_out;
wire _guard13527 = _guard13525 & _guard13526;
wire _guard13528 = fsm_out == 1'd0;
wire _guard13529 = _guard13527 & _guard13528;
wire _guard13530 = fsm_out == 1'd0;
wire _guard13531 = cond_wire415_out;
wire _guard13532 = _guard13530 & _guard13531;
wire _guard13533 = fsm_out == 1'd0;
wire _guard13534 = _guard13532 & _guard13533;
wire _guard13535 = _guard13529 | _guard13534;
wire _guard13536 = early_reset_static_par0_go_out;
wire _guard13537 = _guard13535 & _guard13536;
wire _guard13538 = cond_wire419_out;
wire _guard13539 = early_reset_static_par0_go_out;
wire _guard13540 = _guard13538 & _guard13539;
wire _guard13541 = cond_wire417_out;
wire _guard13542 = early_reset_static_par0_go_out;
wire _guard13543 = _guard13541 & _guard13542;
wire _guard13544 = fsm_out == 1'd0;
wire _guard13545 = cond_wire417_out;
wire _guard13546 = _guard13544 & _guard13545;
wire _guard13547 = fsm_out == 1'd0;
wire _guard13548 = _guard13546 & _guard13547;
wire _guard13549 = fsm_out == 1'd0;
wire _guard13550 = cond_wire419_out;
wire _guard13551 = _guard13549 & _guard13550;
wire _guard13552 = fsm_out == 1'd0;
wire _guard13553 = _guard13551 & _guard13552;
wire _guard13554 = _guard13548 | _guard13553;
wire _guard13555 = early_reset_static_par0_go_out;
wire _guard13556 = _guard13554 & _guard13555;
wire _guard13557 = fsm_out == 1'd0;
wire _guard13558 = cond_wire417_out;
wire _guard13559 = _guard13557 & _guard13558;
wire _guard13560 = fsm_out == 1'd0;
wire _guard13561 = _guard13559 & _guard13560;
wire _guard13562 = fsm_out == 1'd0;
wire _guard13563 = cond_wire419_out;
wire _guard13564 = _guard13562 & _guard13563;
wire _guard13565 = fsm_out == 1'd0;
wire _guard13566 = _guard13564 & _guard13565;
wire _guard13567 = _guard13561 | _guard13566;
wire _guard13568 = early_reset_static_par0_go_out;
wire _guard13569 = _guard13567 & _guard13568;
wire _guard13570 = fsm_out == 1'd0;
wire _guard13571 = cond_wire417_out;
wire _guard13572 = _guard13570 & _guard13571;
wire _guard13573 = fsm_out == 1'd0;
wire _guard13574 = _guard13572 & _guard13573;
wire _guard13575 = fsm_out == 1'd0;
wire _guard13576 = cond_wire419_out;
wire _guard13577 = _guard13575 & _guard13576;
wire _guard13578 = fsm_out == 1'd0;
wire _guard13579 = _guard13577 & _guard13578;
wire _guard13580 = _guard13574 | _guard13579;
wire _guard13581 = early_reset_static_par0_go_out;
wire _guard13582 = _guard13580 & _guard13581;
wire _guard13583 = cond_wire373_out;
wire _guard13584 = early_reset_static_par0_go_out;
wire _guard13585 = _guard13583 & _guard13584;
wire _guard13586 = cond_wire373_out;
wire _guard13587 = early_reset_static_par0_go_out;
wire _guard13588 = _guard13586 & _guard13587;
wire _guard13589 = cond_wire447_out;
wire _guard13590 = early_reset_static_par0_go_out;
wire _guard13591 = _guard13589 & _guard13590;
wire _guard13592 = cond_wire445_out;
wire _guard13593 = early_reset_static_par0_go_out;
wire _guard13594 = _guard13592 & _guard13593;
wire _guard13595 = fsm_out == 1'd0;
wire _guard13596 = cond_wire445_out;
wire _guard13597 = _guard13595 & _guard13596;
wire _guard13598 = fsm_out == 1'd0;
wire _guard13599 = _guard13597 & _guard13598;
wire _guard13600 = fsm_out == 1'd0;
wire _guard13601 = cond_wire447_out;
wire _guard13602 = _guard13600 & _guard13601;
wire _guard13603 = fsm_out == 1'd0;
wire _guard13604 = _guard13602 & _guard13603;
wire _guard13605 = _guard13599 | _guard13604;
wire _guard13606 = early_reset_static_par0_go_out;
wire _guard13607 = _guard13605 & _guard13606;
wire _guard13608 = fsm_out == 1'd0;
wire _guard13609 = cond_wire445_out;
wire _guard13610 = _guard13608 & _guard13609;
wire _guard13611 = fsm_out == 1'd0;
wire _guard13612 = _guard13610 & _guard13611;
wire _guard13613 = fsm_out == 1'd0;
wire _guard13614 = cond_wire447_out;
wire _guard13615 = _guard13613 & _guard13614;
wire _guard13616 = fsm_out == 1'd0;
wire _guard13617 = _guard13615 & _guard13616;
wire _guard13618 = _guard13612 | _guard13617;
wire _guard13619 = early_reset_static_par0_go_out;
wire _guard13620 = _guard13618 & _guard13619;
wire _guard13621 = fsm_out == 1'd0;
wire _guard13622 = cond_wire445_out;
wire _guard13623 = _guard13621 & _guard13622;
wire _guard13624 = fsm_out == 1'd0;
wire _guard13625 = _guard13623 & _guard13624;
wire _guard13626 = fsm_out == 1'd0;
wire _guard13627 = cond_wire447_out;
wire _guard13628 = _guard13626 & _guard13627;
wire _guard13629 = fsm_out == 1'd0;
wire _guard13630 = _guard13628 & _guard13629;
wire _guard13631 = _guard13625 | _guard13630;
wire _guard13632 = early_reset_static_par0_go_out;
wire _guard13633 = _guard13631 & _guard13632;
wire _guard13634 = cond_wire454_out;
wire _guard13635 = early_reset_static_par0_go_out;
wire _guard13636 = _guard13634 & _guard13635;
wire _guard13637 = cond_wire454_out;
wire _guard13638 = early_reset_static_par0_go_out;
wire _guard13639 = _guard13637 & _guard13638;
wire _guard13640 = cond_wire471_out;
wire _guard13641 = early_reset_static_par0_go_out;
wire _guard13642 = _guard13640 & _guard13641;
wire _guard13643 = cond_wire471_out;
wire _guard13644 = early_reset_static_par0_go_out;
wire _guard13645 = _guard13643 & _guard13644;
wire _guard13646 = cond_wire479_out;
wire _guard13647 = early_reset_static_par0_go_out;
wire _guard13648 = _guard13646 & _guard13647;
wire _guard13649 = cond_wire479_out;
wire _guard13650 = early_reset_static_par0_go_out;
wire _guard13651 = _guard13649 & _guard13650;
wire _guard13652 = cond_wire426_out;
wire _guard13653 = early_reset_static_par0_go_out;
wire _guard13654 = _guard13652 & _guard13653;
wire _guard13655 = cond_wire426_out;
wire _guard13656 = early_reset_static_par0_go_out;
wire _guard13657 = _guard13655 & _guard13656;
wire _guard13658 = cond_wire573_out;
wire _guard13659 = early_reset_static_par0_go_out;
wire _guard13660 = _guard13658 & _guard13659;
wire _guard13661 = cond_wire571_out;
wire _guard13662 = early_reset_static_par0_go_out;
wire _guard13663 = _guard13661 & _guard13662;
wire _guard13664 = fsm_out == 1'd0;
wire _guard13665 = cond_wire571_out;
wire _guard13666 = _guard13664 & _guard13665;
wire _guard13667 = fsm_out == 1'd0;
wire _guard13668 = _guard13666 & _guard13667;
wire _guard13669 = fsm_out == 1'd0;
wire _guard13670 = cond_wire573_out;
wire _guard13671 = _guard13669 & _guard13670;
wire _guard13672 = fsm_out == 1'd0;
wire _guard13673 = _guard13671 & _guard13672;
wire _guard13674 = _guard13668 | _guard13673;
wire _guard13675 = early_reset_static_par0_go_out;
wire _guard13676 = _guard13674 & _guard13675;
wire _guard13677 = fsm_out == 1'd0;
wire _guard13678 = cond_wire571_out;
wire _guard13679 = _guard13677 & _guard13678;
wire _guard13680 = fsm_out == 1'd0;
wire _guard13681 = _guard13679 & _guard13680;
wire _guard13682 = fsm_out == 1'd0;
wire _guard13683 = cond_wire573_out;
wire _guard13684 = _guard13682 & _guard13683;
wire _guard13685 = fsm_out == 1'd0;
wire _guard13686 = _guard13684 & _guard13685;
wire _guard13687 = _guard13681 | _guard13686;
wire _guard13688 = early_reset_static_par0_go_out;
wire _guard13689 = _guard13687 & _guard13688;
wire _guard13690 = fsm_out == 1'd0;
wire _guard13691 = cond_wire571_out;
wire _guard13692 = _guard13690 & _guard13691;
wire _guard13693 = fsm_out == 1'd0;
wire _guard13694 = _guard13692 & _guard13693;
wire _guard13695 = fsm_out == 1'd0;
wire _guard13696 = cond_wire573_out;
wire _guard13697 = _guard13695 & _guard13696;
wire _guard13698 = fsm_out == 1'd0;
wire _guard13699 = _guard13697 & _guard13698;
wire _guard13700 = _guard13694 | _guard13699;
wire _guard13701 = early_reset_static_par0_go_out;
wire _guard13702 = _guard13700 & _guard13701;
wire _guard13703 = cond_wire519_out;
wire _guard13704 = early_reset_static_par0_go_out;
wire _guard13705 = _guard13703 & _guard13704;
wire _guard13706 = cond_wire519_out;
wire _guard13707 = early_reset_static_par0_go_out;
wire _guard13708 = _guard13706 & _guard13707;
wire _guard13709 = cond_wire597_out;
wire _guard13710 = early_reset_static_par0_go_out;
wire _guard13711 = _guard13709 & _guard13710;
wire _guard13712 = cond_wire595_out;
wire _guard13713 = early_reset_static_par0_go_out;
wire _guard13714 = _guard13712 & _guard13713;
wire _guard13715 = fsm_out == 1'd0;
wire _guard13716 = cond_wire595_out;
wire _guard13717 = _guard13715 & _guard13716;
wire _guard13718 = fsm_out == 1'd0;
wire _guard13719 = _guard13717 & _guard13718;
wire _guard13720 = fsm_out == 1'd0;
wire _guard13721 = cond_wire597_out;
wire _guard13722 = _guard13720 & _guard13721;
wire _guard13723 = fsm_out == 1'd0;
wire _guard13724 = _guard13722 & _guard13723;
wire _guard13725 = _guard13719 | _guard13724;
wire _guard13726 = early_reset_static_par0_go_out;
wire _guard13727 = _guard13725 & _guard13726;
wire _guard13728 = fsm_out == 1'd0;
wire _guard13729 = cond_wire595_out;
wire _guard13730 = _guard13728 & _guard13729;
wire _guard13731 = fsm_out == 1'd0;
wire _guard13732 = _guard13730 & _guard13731;
wire _guard13733 = fsm_out == 1'd0;
wire _guard13734 = cond_wire597_out;
wire _guard13735 = _guard13733 & _guard13734;
wire _guard13736 = fsm_out == 1'd0;
wire _guard13737 = _guard13735 & _guard13736;
wire _guard13738 = _guard13732 | _guard13737;
wire _guard13739 = early_reset_static_par0_go_out;
wire _guard13740 = _guard13738 & _guard13739;
wire _guard13741 = fsm_out == 1'd0;
wire _guard13742 = cond_wire595_out;
wire _guard13743 = _guard13741 & _guard13742;
wire _guard13744 = fsm_out == 1'd0;
wire _guard13745 = _guard13743 & _guard13744;
wire _guard13746 = fsm_out == 1'd0;
wire _guard13747 = cond_wire597_out;
wire _guard13748 = _guard13746 & _guard13747;
wire _guard13749 = fsm_out == 1'd0;
wire _guard13750 = _guard13748 & _guard13749;
wire _guard13751 = _guard13745 | _guard13750;
wire _guard13752 = early_reset_static_par0_go_out;
wire _guard13753 = _guard13751 & _guard13752;
wire _guard13754 = cond_wire560_out;
wire _guard13755 = early_reset_static_par0_go_out;
wire _guard13756 = _guard13754 & _guard13755;
wire _guard13757 = cond_wire560_out;
wire _guard13758 = early_reset_static_par0_go_out;
wire _guard13759 = _guard13757 & _guard13758;
wire _guard13760 = cond_wire572_out;
wire _guard13761 = early_reset_static_par0_go_out;
wire _guard13762 = _guard13760 & _guard13761;
wire _guard13763 = cond_wire572_out;
wire _guard13764 = early_reset_static_par0_go_out;
wire _guard13765 = _guard13763 & _guard13764;
wire _guard13766 = cond_wire667_out;
wire _guard13767 = early_reset_static_par0_go_out;
wire _guard13768 = _guard13766 & _guard13767;
wire _guard13769 = cond_wire665_out;
wire _guard13770 = early_reset_static_par0_go_out;
wire _guard13771 = _guard13769 & _guard13770;
wire _guard13772 = fsm_out == 1'd0;
wire _guard13773 = cond_wire665_out;
wire _guard13774 = _guard13772 & _guard13773;
wire _guard13775 = fsm_out == 1'd0;
wire _guard13776 = _guard13774 & _guard13775;
wire _guard13777 = fsm_out == 1'd0;
wire _guard13778 = cond_wire667_out;
wire _guard13779 = _guard13777 & _guard13778;
wire _guard13780 = fsm_out == 1'd0;
wire _guard13781 = _guard13779 & _guard13780;
wire _guard13782 = _guard13776 | _guard13781;
wire _guard13783 = early_reset_static_par0_go_out;
wire _guard13784 = _guard13782 & _guard13783;
wire _guard13785 = fsm_out == 1'd0;
wire _guard13786 = cond_wire665_out;
wire _guard13787 = _guard13785 & _guard13786;
wire _guard13788 = fsm_out == 1'd0;
wire _guard13789 = _guard13787 & _guard13788;
wire _guard13790 = fsm_out == 1'd0;
wire _guard13791 = cond_wire667_out;
wire _guard13792 = _guard13790 & _guard13791;
wire _guard13793 = fsm_out == 1'd0;
wire _guard13794 = _guard13792 & _guard13793;
wire _guard13795 = _guard13789 | _guard13794;
wire _guard13796 = early_reset_static_par0_go_out;
wire _guard13797 = _guard13795 & _guard13796;
wire _guard13798 = fsm_out == 1'd0;
wire _guard13799 = cond_wire665_out;
wire _guard13800 = _guard13798 & _guard13799;
wire _guard13801 = fsm_out == 1'd0;
wire _guard13802 = _guard13800 & _guard13801;
wire _guard13803 = fsm_out == 1'd0;
wire _guard13804 = cond_wire667_out;
wire _guard13805 = _guard13803 & _guard13804;
wire _guard13806 = fsm_out == 1'd0;
wire _guard13807 = _guard13805 & _guard13806;
wire _guard13808 = _guard13802 | _guard13807;
wire _guard13809 = early_reset_static_par0_go_out;
wire _guard13810 = _guard13808 & _guard13809;
wire _guard13811 = cond_wire706_out;
wire _guard13812 = early_reset_static_par0_go_out;
wire _guard13813 = _guard13811 & _guard13812;
wire _guard13814 = cond_wire706_out;
wire _guard13815 = early_reset_static_par0_go_out;
wire _guard13816 = _guard13814 & _guard13815;
wire _guard13817 = cond_wire714_out;
wire _guard13818 = early_reset_static_par0_go_out;
wire _guard13819 = _guard13817 & _guard13818;
wire _guard13820 = cond_wire714_out;
wire _guard13821 = early_reset_static_par0_go_out;
wire _guard13822 = _guard13820 & _guard13821;
wire _guard13823 = cond_wire657_out;
wire _guard13824 = early_reset_static_par0_go_out;
wire _guard13825 = _guard13823 & _guard13824;
wire _guard13826 = cond_wire657_out;
wire _guard13827 = early_reset_static_par0_go_out;
wire _guard13828 = _guard13826 & _guard13827;
wire _guard13829 = cond_wire718_out;
wire _guard13830 = early_reset_static_par0_go_out;
wire _guard13831 = _guard13829 & _guard13830;
wire _guard13832 = cond_wire718_out;
wire _guard13833 = early_reset_static_par0_go_out;
wire _guard13834 = _guard13832 & _guard13833;
wire _guard13835 = cond_wire743_out;
wire _guard13836 = early_reset_static_par0_go_out;
wire _guard13837 = _guard13835 & _guard13836;
wire _guard13838 = cond_wire743_out;
wire _guard13839 = early_reset_static_par0_go_out;
wire _guard13840 = _guard13838 & _guard13839;
wire _guard13841 = cond_wire768_out;
wire _guard13842 = early_reset_static_par0_go_out;
wire _guard13843 = _guard13841 & _guard13842;
wire _guard13844 = cond_wire766_out;
wire _guard13845 = early_reset_static_par0_go_out;
wire _guard13846 = _guard13844 & _guard13845;
wire _guard13847 = fsm_out == 1'd0;
wire _guard13848 = cond_wire766_out;
wire _guard13849 = _guard13847 & _guard13848;
wire _guard13850 = fsm_out == 1'd0;
wire _guard13851 = _guard13849 & _guard13850;
wire _guard13852 = fsm_out == 1'd0;
wire _guard13853 = cond_wire768_out;
wire _guard13854 = _guard13852 & _guard13853;
wire _guard13855 = fsm_out == 1'd0;
wire _guard13856 = _guard13854 & _guard13855;
wire _guard13857 = _guard13851 | _guard13856;
wire _guard13858 = early_reset_static_par0_go_out;
wire _guard13859 = _guard13857 & _guard13858;
wire _guard13860 = fsm_out == 1'd0;
wire _guard13861 = cond_wire766_out;
wire _guard13862 = _guard13860 & _guard13861;
wire _guard13863 = fsm_out == 1'd0;
wire _guard13864 = _guard13862 & _guard13863;
wire _guard13865 = fsm_out == 1'd0;
wire _guard13866 = cond_wire768_out;
wire _guard13867 = _guard13865 & _guard13866;
wire _guard13868 = fsm_out == 1'd0;
wire _guard13869 = _guard13867 & _guard13868;
wire _guard13870 = _guard13864 | _guard13869;
wire _guard13871 = early_reset_static_par0_go_out;
wire _guard13872 = _guard13870 & _guard13871;
wire _guard13873 = fsm_out == 1'd0;
wire _guard13874 = cond_wire766_out;
wire _guard13875 = _guard13873 & _guard13874;
wire _guard13876 = fsm_out == 1'd0;
wire _guard13877 = _guard13875 & _guard13876;
wire _guard13878 = fsm_out == 1'd0;
wire _guard13879 = cond_wire768_out;
wire _guard13880 = _guard13878 & _guard13879;
wire _guard13881 = fsm_out == 1'd0;
wire _guard13882 = _guard13880 & _guard13881;
wire _guard13883 = _guard13877 | _guard13882;
wire _guard13884 = early_reset_static_par0_go_out;
wire _guard13885 = _guard13883 & _guard13884;
wire _guard13886 = cond_wire763_out;
wire _guard13887 = early_reset_static_par0_go_out;
wire _guard13888 = _guard13886 & _guard13887;
wire _guard13889 = cond_wire763_out;
wire _guard13890 = early_reset_static_par0_go_out;
wire _guard13891 = _guard13889 & _guard13890;
wire _guard13892 = cond_wire771_out;
wire _guard13893 = early_reset_static_par0_go_out;
wire _guard13894 = _guard13892 & _guard13893;
wire _guard13895 = cond_wire771_out;
wire _guard13896 = early_reset_static_par0_go_out;
wire _guard13897 = _guard13895 & _guard13896;
wire _guard13898 = cond_wire775_out;
wire _guard13899 = early_reset_static_par0_go_out;
wire _guard13900 = _guard13898 & _guard13899;
wire _guard13901 = cond_wire775_out;
wire _guard13902 = early_reset_static_par0_go_out;
wire _guard13903 = _guard13901 & _guard13902;
wire _guard13904 = cond_wire836_out;
wire _guard13905 = early_reset_static_par0_go_out;
wire _guard13906 = _guard13904 & _guard13905;
wire _guard13907 = cond_wire836_out;
wire _guard13908 = early_reset_static_par0_go_out;
wire _guard13909 = _guard13907 & _guard13908;
wire _guard13910 = cond_wire859_out;
wire _guard13911 = early_reset_static_par0_go_out;
wire _guard13912 = _guard13910 & _guard13911;
wire _guard13913 = cond_wire859_out;
wire _guard13914 = early_reset_static_par0_go_out;
wire _guard13915 = _guard13913 & _guard13914;
wire _guard13916 = cond_wire861_out;
wire _guard13917 = early_reset_static_par0_go_out;
wire _guard13918 = _guard13916 & _guard13917;
wire _guard13919 = cond_wire861_out;
wire _guard13920 = early_reset_static_par0_go_out;
wire _guard13921 = _guard13919 & _guard13920;
wire _guard13922 = cond_wire882_out;
wire _guard13923 = early_reset_static_par0_go_out;
wire _guard13924 = _guard13922 & _guard13923;
wire _guard13925 = cond_wire880_out;
wire _guard13926 = early_reset_static_par0_go_out;
wire _guard13927 = _guard13925 & _guard13926;
wire _guard13928 = fsm_out == 1'd0;
wire _guard13929 = cond_wire880_out;
wire _guard13930 = _guard13928 & _guard13929;
wire _guard13931 = fsm_out == 1'd0;
wire _guard13932 = _guard13930 & _guard13931;
wire _guard13933 = fsm_out == 1'd0;
wire _guard13934 = cond_wire882_out;
wire _guard13935 = _guard13933 & _guard13934;
wire _guard13936 = fsm_out == 1'd0;
wire _guard13937 = _guard13935 & _guard13936;
wire _guard13938 = _guard13932 | _guard13937;
wire _guard13939 = early_reset_static_par0_go_out;
wire _guard13940 = _guard13938 & _guard13939;
wire _guard13941 = fsm_out == 1'd0;
wire _guard13942 = cond_wire880_out;
wire _guard13943 = _guard13941 & _guard13942;
wire _guard13944 = fsm_out == 1'd0;
wire _guard13945 = _guard13943 & _guard13944;
wire _guard13946 = fsm_out == 1'd0;
wire _guard13947 = cond_wire882_out;
wire _guard13948 = _guard13946 & _guard13947;
wire _guard13949 = fsm_out == 1'd0;
wire _guard13950 = _guard13948 & _guard13949;
wire _guard13951 = _guard13945 | _guard13950;
wire _guard13952 = early_reset_static_par0_go_out;
wire _guard13953 = _guard13951 & _guard13952;
wire _guard13954 = fsm_out == 1'd0;
wire _guard13955 = cond_wire880_out;
wire _guard13956 = _guard13954 & _guard13955;
wire _guard13957 = fsm_out == 1'd0;
wire _guard13958 = _guard13956 & _guard13957;
wire _guard13959 = fsm_out == 1'd0;
wire _guard13960 = cond_wire882_out;
wire _guard13961 = _guard13959 & _guard13960;
wire _guard13962 = fsm_out == 1'd0;
wire _guard13963 = _guard13961 & _guard13962;
wire _guard13964 = _guard13958 | _guard13963;
wire _guard13965 = early_reset_static_par0_go_out;
wire _guard13966 = _guard13964 & _guard13965;
wire _guard13967 = cond_wire886_out;
wire _guard13968 = early_reset_static_par0_go_out;
wire _guard13969 = _guard13967 & _guard13968;
wire _guard13970 = cond_wire884_out;
wire _guard13971 = early_reset_static_par0_go_out;
wire _guard13972 = _guard13970 & _guard13971;
wire _guard13973 = fsm_out == 1'd0;
wire _guard13974 = cond_wire884_out;
wire _guard13975 = _guard13973 & _guard13974;
wire _guard13976 = fsm_out == 1'd0;
wire _guard13977 = _guard13975 & _guard13976;
wire _guard13978 = fsm_out == 1'd0;
wire _guard13979 = cond_wire886_out;
wire _guard13980 = _guard13978 & _guard13979;
wire _guard13981 = fsm_out == 1'd0;
wire _guard13982 = _guard13980 & _guard13981;
wire _guard13983 = _guard13977 | _guard13982;
wire _guard13984 = early_reset_static_par0_go_out;
wire _guard13985 = _guard13983 & _guard13984;
wire _guard13986 = fsm_out == 1'd0;
wire _guard13987 = cond_wire884_out;
wire _guard13988 = _guard13986 & _guard13987;
wire _guard13989 = fsm_out == 1'd0;
wire _guard13990 = _guard13988 & _guard13989;
wire _guard13991 = fsm_out == 1'd0;
wire _guard13992 = cond_wire886_out;
wire _guard13993 = _guard13991 & _guard13992;
wire _guard13994 = fsm_out == 1'd0;
wire _guard13995 = _guard13993 & _guard13994;
wire _guard13996 = _guard13990 | _guard13995;
wire _guard13997 = early_reset_static_par0_go_out;
wire _guard13998 = _guard13996 & _guard13997;
wire _guard13999 = fsm_out == 1'd0;
wire _guard14000 = cond_wire884_out;
wire _guard14001 = _guard13999 & _guard14000;
wire _guard14002 = fsm_out == 1'd0;
wire _guard14003 = _guard14001 & _guard14002;
wire _guard14004 = fsm_out == 1'd0;
wire _guard14005 = cond_wire886_out;
wire _guard14006 = _guard14004 & _guard14005;
wire _guard14007 = fsm_out == 1'd0;
wire _guard14008 = _guard14006 & _guard14007;
wire _guard14009 = _guard14003 | _guard14008;
wire _guard14010 = early_reset_static_par0_go_out;
wire _guard14011 = _guard14009 & _guard14010;
wire _guard14012 = cond_wire881_out;
wire _guard14013 = early_reset_static_par0_go_out;
wire _guard14014 = _guard14012 & _guard14013;
wire _guard14015 = cond_wire881_out;
wire _guard14016 = early_reset_static_par0_go_out;
wire _guard14017 = _guard14015 & _guard14016;
wire _guard14018 = cond_wire894_out;
wire _guard14019 = early_reset_static_par0_go_out;
wire _guard14020 = _guard14018 & _guard14019;
wire _guard14021 = cond_wire892_out;
wire _guard14022 = early_reset_static_par0_go_out;
wire _guard14023 = _guard14021 & _guard14022;
wire _guard14024 = fsm_out == 1'd0;
wire _guard14025 = cond_wire892_out;
wire _guard14026 = _guard14024 & _guard14025;
wire _guard14027 = fsm_out == 1'd0;
wire _guard14028 = _guard14026 & _guard14027;
wire _guard14029 = fsm_out == 1'd0;
wire _guard14030 = cond_wire894_out;
wire _guard14031 = _guard14029 & _guard14030;
wire _guard14032 = fsm_out == 1'd0;
wire _guard14033 = _guard14031 & _guard14032;
wire _guard14034 = _guard14028 | _guard14033;
wire _guard14035 = early_reset_static_par0_go_out;
wire _guard14036 = _guard14034 & _guard14035;
wire _guard14037 = fsm_out == 1'd0;
wire _guard14038 = cond_wire892_out;
wire _guard14039 = _guard14037 & _guard14038;
wire _guard14040 = fsm_out == 1'd0;
wire _guard14041 = _guard14039 & _guard14040;
wire _guard14042 = fsm_out == 1'd0;
wire _guard14043 = cond_wire894_out;
wire _guard14044 = _guard14042 & _guard14043;
wire _guard14045 = fsm_out == 1'd0;
wire _guard14046 = _guard14044 & _guard14045;
wire _guard14047 = _guard14041 | _guard14046;
wire _guard14048 = early_reset_static_par0_go_out;
wire _guard14049 = _guard14047 & _guard14048;
wire _guard14050 = fsm_out == 1'd0;
wire _guard14051 = cond_wire892_out;
wire _guard14052 = _guard14050 & _guard14051;
wire _guard14053 = fsm_out == 1'd0;
wire _guard14054 = _guard14052 & _guard14053;
wire _guard14055 = fsm_out == 1'd0;
wire _guard14056 = cond_wire894_out;
wire _guard14057 = _guard14055 & _guard14056;
wire _guard14058 = fsm_out == 1'd0;
wire _guard14059 = _guard14057 & _guard14058;
wire _guard14060 = _guard14054 | _guard14059;
wire _guard14061 = early_reset_static_par0_go_out;
wire _guard14062 = _guard14060 & _guard14061;
wire _guard14063 = cond_wire910_out;
wire _guard14064 = early_reset_static_par0_go_out;
wire _guard14065 = _guard14063 & _guard14064;
wire _guard14066 = cond_wire908_out;
wire _guard14067 = early_reset_static_par0_go_out;
wire _guard14068 = _guard14066 & _guard14067;
wire _guard14069 = fsm_out == 1'd0;
wire _guard14070 = cond_wire908_out;
wire _guard14071 = _guard14069 & _guard14070;
wire _guard14072 = fsm_out == 1'd0;
wire _guard14073 = _guard14071 & _guard14072;
wire _guard14074 = fsm_out == 1'd0;
wire _guard14075 = cond_wire910_out;
wire _guard14076 = _guard14074 & _guard14075;
wire _guard14077 = fsm_out == 1'd0;
wire _guard14078 = _guard14076 & _guard14077;
wire _guard14079 = _guard14073 | _guard14078;
wire _guard14080 = early_reset_static_par0_go_out;
wire _guard14081 = _guard14079 & _guard14080;
wire _guard14082 = fsm_out == 1'd0;
wire _guard14083 = cond_wire908_out;
wire _guard14084 = _guard14082 & _guard14083;
wire _guard14085 = fsm_out == 1'd0;
wire _guard14086 = _guard14084 & _guard14085;
wire _guard14087 = fsm_out == 1'd0;
wire _guard14088 = cond_wire910_out;
wire _guard14089 = _guard14087 & _guard14088;
wire _guard14090 = fsm_out == 1'd0;
wire _guard14091 = _guard14089 & _guard14090;
wire _guard14092 = _guard14086 | _guard14091;
wire _guard14093 = early_reset_static_par0_go_out;
wire _guard14094 = _guard14092 & _guard14093;
wire _guard14095 = fsm_out == 1'd0;
wire _guard14096 = cond_wire908_out;
wire _guard14097 = _guard14095 & _guard14096;
wire _guard14098 = fsm_out == 1'd0;
wire _guard14099 = _guard14097 & _guard14098;
wire _guard14100 = fsm_out == 1'd0;
wire _guard14101 = cond_wire910_out;
wire _guard14102 = _guard14100 & _guard14101;
wire _guard14103 = fsm_out == 1'd0;
wire _guard14104 = _guard14102 & _guard14103;
wire _guard14105 = _guard14099 | _guard14104;
wire _guard14106 = early_reset_static_par0_go_out;
wire _guard14107 = _guard14105 & _guard14106;
wire _guard14108 = cond_wire943_out;
wire _guard14109 = early_reset_static_par0_go_out;
wire _guard14110 = _guard14108 & _guard14109;
wire _guard14111 = cond_wire941_out;
wire _guard14112 = early_reset_static_par0_go_out;
wire _guard14113 = _guard14111 & _guard14112;
wire _guard14114 = fsm_out == 1'd0;
wire _guard14115 = cond_wire941_out;
wire _guard14116 = _guard14114 & _guard14115;
wire _guard14117 = fsm_out == 1'd0;
wire _guard14118 = _guard14116 & _guard14117;
wire _guard14119 = fsm_out == 1'd0;
wire _guard14120 = cond_wire943_out;
wire _guard14121 = _guard14119 & _guard14120;
wire _guard14122 = fsm_out == 1'd0;
wire _guard14123 = _guard14121 & _guard14122;
wire _guard14124 = _guard14118 | _guard14123;
wire _guard14125 = early_reset_static_par0_go_out;
wire _guard14126 = _guard14124 & _guard14125;
wire _guard14127 = fsm_out == 1'd0;
wire _guard14128 = cond_wire941_out;
wire _guard14129 = _guard14127 & _guard14128;
wire _guard14130 = fsm_out == 1'd0;
wire _guard14131 = _guard14129 & _guard14130;
wire _guard14132 = fsm_out == 1'd0;
wire _guard14133 = cond_wire943_out;
wire _guard14134 = _guard14132 & _guard14133;
wire _guard14135 = fsm_out == 1'd0;
wire _guard14136 = _guard14134 & _guard14135;
wire _guard14137 = _guard14131 | _guard14136;
wire _guard14138 = early_reset_static_par0_go_out;
wire _guard14139 = _guard14137 & _guard14138;
wire _guard14140 = fsm_out == 1'd0;
wire _guard14141 = cond_wire941_out;
wire _guard14142 = _guard14140 & _guard14141;
wire _guard14143 = fsm_out == 1'd0;
wire _guard14144 = _guard14142 & _guard14143;
wire _guard14145 = fsm_out == 1'd0;
wire _guard14146 = cond_wire943_out;
wire _guard14147 = _guard14145 & _guard14146;
wire _guard14148 = fsm_out == 1'd0;
wire _guard14149 = _guard14147 & _guard14148;
wire _guard14150 = _guard14144 | _guard14149;
wire _guard14151 = early_reset_static_par0_go_out;
wire _guard14152 = _guard14150 & _guard14151;
wire _guard14153 = cond_wire946_out;
wire _guard14154 = early_reset_static_par0_go_out;
wire _guard14155 = _guard14153 & _guard14154;
wire _guard14156 = cond_wire946_out;
wire _guard14157 = early_reset_static_par0_go_out;
wire _guard14158 = _guard14156 & _guard14157;
wire _guard14159 = cond_wire975_out;
wire _guard14160 = early_reset_static_par0_go_out;
wire _guard14161 = _guard14159 & _guard14160;
wire _guard14162 = cond_wire973_out;
wire _guard14163 = early_reset_static_par0_go_out;
wire _guard14164 = _guard14162 & _guard14163;
wire _guard14165 = fsm_out == 1'd0;
wire _guard14166 = cond_wire973_out;
wire _guard14167 = _guard14165 & _guard14166;
wire _guard14168 = fsm_out == 1'd0;
wire _guard14169 = _guard14167 & _guard14168;
wire _guard14170 = fsm_out == 1'd0;
wire _guard14171 = cond_wire975_out;
wire _guard14172 = _guard14170 & _guard14171;
wire _guard14173 = fsm_out == 1'd0;
wire _guard14174 = _guard14172 & _guard14173;
wire _guard14175 = _guard14169 | _guard14174;
wire _guard14176 = early_reset_static_par0_go_out;
wire _guard14177 = _guard14175 & _guard14176;
wire _guard14178 = fsm_out == 1'd0;
wire _guard14179 = cond_wire973_out;
wire _guard14180 = _guard14178 & _guard14179;
wire _guard14181 = fsm_out == 1'd0;
wire _guard14182 = _guard14180 & _guard14181;
wire _guard14183 = fsm_out == 1'd0;
wire _guard14184 = cond_wire975_out;
wire _guard14185 = _guard14183 & _guard14184;
wire _guard14186 = fsm_out == 1'd0;
wire _guard14187 = _guard14185 & _guard14186;
wire _guard14188 = _guard14182 | _guard14187;
wire _guard14189 = early_reset_static_par0_go_out;
wire _guard14190 = _guard14188 & _guard14189;
wire _guard14191 = fsm_out == 1'd0;
wire _guard14192 = cond_wire973_out;
wire _guard14193 = _guard14191 & _guard14192;
wire _guard14194 = fsm_out == 1'd0;
wire _guard14195 = _guard14193 & _guard14194;
wire _guard14196 = fsm_out == 1'd0;
wire _guard14197 = cond_wire975_out;
wire _guard14198 = _guard14196 & _guard14197;
wire _guard14199 = fsm_out == 1'd0;
wire _guard14200 = _guard14198 & _guard14199;
wire _guard14201 = _guard14195 | _guard14200;
wire _guard14202 = early_reset_static_par0_go_out;
wire _guard14203 = _guard14201 & _guard14202;
wire _guard14204 = cond_wire987_out;
wire _guard14205 = early_reset_static_par0_go_out;
wire _guard14206 = _guard14204 & _guard14205;
wire _guard14207 = cond_wire985_out;
wire _guard14208 = early_reset_static_par0_go_out;
wire _guard14209 = _guard14207 & _guard14208;
wire _guard14210 = fsm_out == 1'd0;
wire _guard14211 = cond_wire985_out;
wire _guard14212 = _guard14210 & _guard14211;
wire _guard14213 = fsm_out == 1'd0;
wire _guard14214 = _guard14212 & _guard14213;
wire _guard14215 = fsm_out == 1'd0;
wire _guard14216 = cond_wire987_out;
wire _guard14217 = _guard14215 & _guard14216;
wire _guard14218 = fsm_out == 1'd0;
wire _guard14219 = _guard14217 & _guard14218;
wire _guard14220 = _guard14214 | _guard14219;
wire _guard14221 = early_reset_static_par0_go_out;
wire _guard14222 = _guard14220 & _guard14221;
wire _guard14223 = fsm_out == 1'd0;
wire _guard14224 = cond_wire985_out;
wire _guard14225 = _guard14223 & _guard14224;
wire _guard14226 = fsm_out == 1'd0;
wire _guard14227 = _guard14225 & _guard14226;
wire _guard14228 = fsm_out == 1'd0;
wire _guard14229 = cond_wire987_out;
wire _guard14230 = _guard14228 & _guard14229;
wire _guard14231 = fsm_out == 1'd0;
wire _guard14232 = _guard14230 & _guard14231;
wire _guard14233 = _guard14227 | _guard14232;
wire _guard14234 = early_reset_static_par0_go_out;
wire _guard14235 = _guard14233 & _guard14234;
wire _guard14236 = fsm_out == 1'd0;
wire _guard14237 = cond_wire985_out;
wire _guard14238 = _guard14236 & _guard14237;
wire _guard14239 = fsm_out == 1'd0;
wire _guard14240 = _guard14238 & _guard14239;
wire _guard14241 = fsm_out == 1'd0;
wire _guard14242 = cond_wire987_out;
wire _guard14243 = _guard14241 & _guard14242;
wire _guard14244 = fsm_out == 1'd0;
wire _guard14245 = _guard14243 & _guard14244;
wire _guard14246 = _guard14240 | _guard14245;
wire _guard14247 = early_reset_static_par0_go_out;
wire _guard14248 = _guard14246 & _guard14247;
wire _guard14249 = cond_wire992_out;
wire _guard14250 = early_reset_static_par0_go_out;
wire _guard14251 = _guard14249 & _guard14250;
wire _guard14252 = cond_wire990_out;
wire _guard14253 = early_reset_static_par0_go_out;
wire _guard14254 = _guard14252 & _guard14253;
wire _guard14255 = fsm_out == 1'd0;
wire _guard14256 = cond_wire990_out;
wire _guard14257 = _guard14255 & _guard14256;
wire _guard14258 = fsm_out == 1'd0;
wire _guard14259 = _guard14257 & _guard14258;
wire _guard14260 = fsm_out == 1'd0;
wire _guard14261 = cond_wire992_out;
wire _guard14262 = _guard14260 & _guard14261;
wire _guard14263 = fsm_out == 1'd0;
wire _guard14264 = _guard14262 & _guard14263;
wire _guard14265 = _guard14259 | _guard14264;
wire _guard14266 = early_reset_static_par0_go_out;
wire _guard14267 = _guard14265 & _guard14266;
wire _guard14268 = fsm_out == 1'd0;
wire _guard14269 = cond_wire990_out;
wire _guard14270 = _guard14268 & _guard14269;
wire _guard14271 = fsm_out == 1'd0;
wire _guard14272 = _guard14270 & _guard14271;
wire _guard14273 = fsm_out == 1'd0;
wire _guard14274 = cond_wire992_out;
wire _guard14275 = _guard14273 & _guard14274;
wire _guard14276 = fsm_out == 1'd0;
wire _guard14277 = _guard14275 & _guard14276;
wire _guard14278 = _guard14272 | _guard14277;
wire _guard14279 = early_reset_static_par0_go_out;
wire _guard14280 = _guard14278 & _guard14279;
wire _guard14281 = fsm_out == 1'd0;
wire _guard14282 = cond_wire990_out;
wire _guard14283 = _guard14281 & _guard14282;
wire _guard14284 = fsm_out == 1'd0;
wire _guard14285 = _guard14283 & _guard14284;
wire _guard14286 = fsm_out == 1'd0;
wire _guard14287 = cond_wire992_out;
wire _guard14288 = _guard14286 & _guard14287;
wire _guard14289 = fsm_out == 1'd0;
wire _guard14290 = _guard14288 & _guard14289;
wire _guard14291 = _guard14285 | _guard14290;
wire _guard14292 = early_reset_static_par0_go_out;
wire _guard14293 = _guard14291 & _guard14292;
wire _guard14294 = cond_wire995_out;
wire _guard14295 = early_reset_static_par0_go_out;
wire _guard14296 = _guard14294 & _guard14295;
wire _guard14297 = cond_wire995_out;
wire _guard14298 = early_reset_static_par0_go_out;
wire _guard14299 = _guard14297 & _guard14298;
wire _guard14300 = cond_wire938_out;
wire _guard14301 = early_reset_static_par0_go_out;
wire _guard14302 = _guard14300 & _guard14301;
wire _guard14303 = cond_wire938_out;
wire _guard14304 = early_reset_static_par0_go_out;
wire _guard14305 = _guard14303 & _guard14304;
wire _guard14306 = cond_wire19_out;
wire _guard14307 = early_reset_static_par0_go_out;
wire _guard14308 = _guard14306 & _guard14307;
wire _guard14309 = cond_wire19_out;
wire _guard14310 = early_reset_static_par0_go_out;
wire _guard14311 = _guard14309 & _guard14310;
wire _guard14312 = fsm0_out == 6'd0;
wire _guard14313 = early_reset_static_seq_go_out;
wire _guard14314 = _guard14312 & _guard14313;
wire _guard14315 = cond_wire24_out;
wire _guard14316 = early_reset_static_par0_go_out;
wire _guard14317 = _guard14315 & _guard14316;
wire _guard14318 = _guard14314 | _guard14317;
wire _guard14319 = fsm0_out == 6'd0;
wire _guard14320 = early_reset_static_seq_go_out;
wire _guard14321 = _guard14319 & _guard14320;
wire _guard14322 = cond_wire24_out;
wire _guard14323 = early_reset_static_par0_go_out;
wire _guard14324 = _guard14322 & _guard14323;
wire _guard14325 = cond_wire29_out;
wire _guard14326 = early_reset_static_par0_go_out;
wire _guard14327 = _guard14325 & _guard14326;
wire _guard14328 = cond_wire29_out;
wire _guard14329 = early_reset_static_par0_go_out;
wire _guard14330 = _guard14328 & _guard14329;
wire _guard14331 = cond_wire49_out;
wire _guard14332 = early_reset_static_par0_go_out;
wire _guard14333 = _guard14331 & _guard14332;
wire _guard14334 = cond_wire49_out;
wire _guard14335 = early_reset_static_par0_go_out;
wire _guard14336 = _guard14334 & _guard14335;
wire _guard14337 = cond_wire74_out;
wire _guard14338 = early_reset_static_par0_go_out;
wire _guard14339 = _guard14337 & _guard14338;
wire _guard14340 = cond_wire74_out;
wire _guard14341 = early_reset_static_par0_go_out;
wire _guard14342 = _guard14340 & _guard14341;
wire _guard14343 = fsm0_out == 6'd0;
wire _guard14344 = early_reset_static_seq_go_out;
wire _guard14345 = _guard14343 & _guard14344;
wire _guard14346 = cond_wire924_out;
wire _guard14347 = early_reset_static_par0_go_out;
wire _guard14348 = _guard14346 & _guard14347;
wire _guard14349 = _guard14345 | _guard14348;
wire _guard14350 = fsm0_out == 6'd0;
wire _guard14351 = early_reset_static_seq_go_out;
wire _guard14352 = _guard14350 & _guard14351;
wire _guard14353 = cond_wire924_out;
wire _guard14354 = early_reset_static_par0_go_out;
wire _guard14355 = _guard14353 & _guard14354;
wire _guard14356 = fsm0_out == 6'd0;
wire _guard14357 = early_reset_static_seq_go_out;
wire _guard14358 = _guard14356 & _guard14357;
wire _guard14359 = early_reset_static_par0_go_out;
wire _guard14360 = _guard14358 | _guard14359;
wire _guard14361 = early_reset_static_par0_go_out;
wire _guard14362 = fsm0_out == 6'd0;
wire _guard14363 = early_reset_static_seq_go_out;
wire _guard14364 = _guard14362 & _guard14363;
wire _guard14365 = early_reset_static_par0_go_out;
wire _guard14366 = early_reset_static_par0_go_out;
wire _guard14367 = early_reset_static_par0_go_out;
wire _guard14368 = early_reset_static_par0_go_out;
wire _guard14369 = fsm0_out == 6'd0;
wire _guard14370 = early_reset_static_seq_go_out;
wire _guard14371 = _guard14369 & _guard14370;
wire _guard14372 = early_reset_static_par0_go_out;
wire _guard14373 = _guard14371 | _guard14372;
wire _guard14374 = fsm0_out == 6'd0;
wire _guard14375 = early_reset_static_seq_go_out;
wire _guard14376 = _guard14374 & _guard14375;
wire _guard14377 = early_reset_static_par0_go_out;
wire _guard14378 = early_reset_static_par0_go_out;
wire _guard14379 = early_reset_static_par0_go_out;
wire _guard14380 = early_reset_static_par0_go_out;
wire _guard14381 = early_reset_static_par0_go_out;
wire _guard14382 = fsm0_out == 6'd0;
wire _guard14383 = early_reset_static_seq_go_out;
wire _guard14384 = _guard14382 & _guard14383;
wire _guard14385 = early_reset_static_par0_go_out;
wire _guard14386 = _guard14384 | _guard14385;
wire _guard14387 = early_reset_static_par0_go_out;
wire _guard14388 = fsm0_out == 6'd0;
wire _guard14389 = early_reset_static_seq_go_out;
wire _guard14390 = _guard14388 & _guard14389;
wire _guard14391 = fsm0_out == 6'd0;
wire _guard14392 = early_reset_static_seq_go_out;
wire _guard14393 = _guard14391 & _guard14392;
wire _guard14394 = early_reset_static_par0_go_out;
wire _guard14395 = _guard14393 | _guard14394;
wire _guard14396 = early_reset_static_par0_go_out;
wire _guard14397 = fsm0_out == 6'd0;
wire _guard14398 = early_reset_static_seq_go_out;
wire _guard14399 = _guard14397 & _guard14398;
wire _guard14400 = fsm0_out == 6'd0;
wire _guard14401 = early_reset_static_seq_go_out;
wire _guard14402 = _guard14400 & _guard14401;
wire _guard14403 = early_reset_static_par0_go_out;
wire _guard14404 = _guard14402 | _guard14403;
wire _guard14405 = early_reset_static_par0_go_out;
wire _guard14406 = fsm0_out == 6'd0;
wire _guard14407 = early_reset_static_seq_go_out;
wire _guard14408 = _guard14406 & _guard14407;
wire _guard14409 = fsm0_out == 6'd0;
wire _guard14410 = early_reset_static_seq_go_out;
wire _guard14411 = _guard14409 & _guard14410;
wire _guard14412 = early_reset_static_par0_go_out;
wire _guard14413 = _guard14411 | _guard14412;
wire _guard14414 = fsm0_out == 6'd0;
wire _guard14415 = early_reset_static_seq_go_out;
wire _guard14416 = _guard14414 & _guard14415;
wire _guard14417 = early_reset_static_par0_go_out;
wire _guard14418 = fsm0_out == 6'd0;
wire _guard14419 = early_reset_static_seq_go_out;
wire _guard14420 = _guard14418 & _guard14419;
wire _guard14421 = early_reset_static_par0_go_out;
wire _guard14422 = _guard14420 | _guard14421;
wire _guard14423 = early_reset_static_par0_go_out;
wire _guard14424 = fsm0_out == 6'd0;
wire _guard14425 = early_reset_static_seq_go_out;
wire _guard14426 = _guard14424 & _guard14425;
wire _guard14427 = early_reset_static_par0_go_out;
wire _guard14428 = early_reset_static_par0_go_out;
wire _guard14429 = early_reset_static_par0_go_out;
wire _guard14430 = early_reset_static_par0_go_out;
wire _guard14431 = early_reset_static_par0_go_out;
wire _guard14432 = early_reset_static_par0_go_out;
wire _guard14433 = fsm0_out == 6'd0;
wire _guard14434 = early_reset_static_seq_go_out;
wire _guard14435 = _guard14433 & _guard14434;
wire _guard14436 = early_reset_static_par0_go_out;
wire _guard14437 = _guard14435 | _guard14436;
wire _guard14438 = early_reset_static_par0_go_out;
wire _guard14439 = fsm0_out == 6'd0;
wire _guard14440 = early_reset_static_seq_go_out;
wire _guard14441 = _guard14439 & _guard14440;
wire _guard14442 = early_reset_static_par0_go_out;
wire _guard14443 = early_reset_static_par0_go_out;
wire _guard14444 = early_reset_static_par0_go_out;
wire _guard14445 = early_reset_static_par0_go_out;
wire _guard14446 = early_reset_static_par0_go_out;
wire _guard14447 = ~_guard0;
wire _guard14448 = early_reset_static_par0_go_out;
wire _guard14449 = _guard14447 & _guard14448;
wire _guard14450 = early_reset_static_par0_go_out;
wire _guard14451 = early_reset_static_par0_go_out;
wire _guard14452 = early_reset_static_par0_go_out;
wire _guard14453 = early_reset_static_par0_go_out;
wire _guard14454 = early_reset_static_par0_go_out;
wire _guard14455 = ~_guard0;
wire _guard14456 = early_reset_static_par0_go_out;
wire _guard14457 = _guard14455 & _guard14456;
wire _guard14458 = early_reset_static_par0_go_out;
wire _guard14459 = early_reset_static_par0_go_out;
wire _guard14460 = early_reset_static_par0_go_out;
wire _guard14461 = early_reset_static_par0_go_out;
wire _guard14462 = early_reset_static_par0_go_out;
wire _guard14463 = early_reset_static_par0_go_out;
wire _guard14464 = early_reset_static_par0_go_out;
wire _guard14465 = early_reset_static_par0_go_out;
wire _guard14466 = early_reset_static_par0_go_out;
wire _guard14467 = early_reset_static_par0_go_out;
wire _guard14468 = early_reset_static_par0_go_out;
wire _guard14469 = early_reset_static_par0_go_out;
wire _guard14470 = ~_guard0;
wire _guard14471 = early_reset_static_par0_go_out;
wire _guard14472 = _guard14470 & _guard14471;
wire _guard14473 = early_reset_static_par0_go_out;
wire _guard14474 = ~_guard0;
wire _guard14475 = early_reset_static_par0_go_out;
wire _guard14476 = _guard14474 & _guard14475;
wire _guard14477 = early_reset_static_par0_go_out;
wire _guard14478 = early_reset_static_par0_go_out;
wire _guard14479 = ~_guard0;
wire _guard14480 = early_reset_static_par0_go_out;
wire _guard14481 = _guard14479 & _guard14480;
wire _guard14482 = early_reset_static_par0_go_out;
wire _guard14483 = early_reset_static_par0_go_out;
wire _guard14484 = early_reset_static_par0_go_out;
wire _guard14485 = early_reset_static_par0_go_out;
wire _guard14486 = early_reset_static_par0_go_out;
wire _guard14487 = early_reset_static_par0_go_out;
wire _guard14488 = ~_guard0;
wire _guard14489 = early_reset_static_par0_go_out;
wire _guard14490 = _guard14488 & _guard14489;
wire _guard14491 = early_reset_static_par0_go_out;
wire _guard14492 = early_reset_static_par0_go_out;
wire _guard14493 = early_reset_static_par0_go_out;
wire _guard14494 = early_reset_static_par0_go_out;
wire _guard14495 = early_reset_static_par0_go_out;
wire _guard14496 = early_reset_static_par0_go_out;
wire _guard14497 = ~_guard0;
wire _guard14498 = early_reset_static_par0_go_out;
wire _guard14499 = _guard14497 & _guard14498;
wire _guard14500 = early_reset_static_par0_go_out;
wire _guard14501 = early_reset_static_par0_go_out;
wire _guard14502 = early_reset_static_par0_go_out;
wire _guard14503 = ~_guard0;
wire _guard14504 = early_reset_static_par0_go_out;
wire _guard14505 = _guard14503 & _guard14504;
wire _guard14506 = early_reset_static_par0_go_out;
wire _guard14507 = early_reset_static_par0_go_out;
wire _guard14508 = early_reset_static_par0_go_out;
wire _guard14509 = early_reset_static_par0_go_out;
wire _guard14510 = ~_guard0;
wire _guard14511 = early_reset_static_par0_go_out;
wire _guard14512 = _guard14510 & _guard14511;
wire _guard14513 = early_reset_static_par0_go_out;
wire _guard14514 = early_reset_static_par0_go_out;
wire _guard14515 = early_reset_static_par0_go_out;
wire _guard14516 = early_reset_static_par0_go_out;
wire _guard14517 = early_reset_static_par0_go_out;
wire _guard14518 = early_reset_static_par0_go_out;
wire _guard14519 = ~_guard0;
wire _guard14520 = early_reset_static_par0_go_out;
wire _guard14521 = _guard14519 & _guard14520;
wire _guard14522 = early_reset_static_par0_go_out;
wire _guard14523 = early_reset_static_par0_go_out;
wire _guard14524 = early_reset_static_par0_go_out;
wire _guard14525 = ~_guard0;
wire _guard14526 = early_reset_static_par0_go_out;
wire _guard14527 = _guard14525 & _guard14526;
wire _guard14528 = early_reset_static_par0_go_out;
wire _guard14529 = ~_guard0;
wire _guard14530 = early_reset_static_par0_go_out;
wire _guard14531 = _guard14529 & _guard14530;
wire _guard14532 = early_reset_static_par0_go_out;
wire _guard14533 = early_reset_static_par0_go_out;
wire _guard14534 = early_reset_static_par0_go_out;
wire _guard14535 = ~_guard0;
wire _guard14536 = early_reset_static_par0_go_out;
wire _guard14537 = _guard14535 & _guard14536;
wire _guard14538 = early_reset_static_par0_go_out;
wire _guard14539 = early_reset_static_par0_go_out;
wire _guard14540 = early_reset_static_par0_go_out;
wire _guard14541 = early_reset_static_par0_go_out;
wire _guard14542 = early_reset_static_par0_go_out;
wire _guard14543 = ~_guard0;
wire _guard14544 = early_reset_static_par0_go_out;
wire _guard14545 = _guard14543 & _guard14544;
wire _guard14546 = ~_guard0;
wire _guard14547 = early_reset_static_par0_go_out;
wire _guard14548 = _guard14546 & _guard14547;
wire _guard14549 = early_reset_static_par0_go_out;
wire _guard14550 = early_reset_static_par0_go_out;
wire _guard14551 = early_reset_static_par0_go_out;
wire _guard14552 = ~_guard0;
wire _guard14553 = early_reset_static_par0_go_out;
wire _guard14554 = _guard14552 & _guard14553;
wire _guard14555 = early_reset_static_par0_go_out;
wire _guard14556 = early_reset_static_par0_go_out;
wire _guard14557 = ~_guard0;
wire _guard14558 = early_reset_static_par0_go_out;
wire _guard14559 = _guard14557 & _guard14558;
wire _guard14560 = early_reset_static_par0_go_out;
wire _guard14561 = ~_guard0;
wire _guard14562 = early_reset_static_par0_go_out;
wire _guard14563 = _guard14561 & _guard14562;
wire _guard14564 = early_reset_static_par0_go_out;
wire _guard14565 = early_reset_static_par0_go_out;
wire _guard14566 = early_reset_static_par0_go_out;
wire _guard14567 = early_reset_static_par0_go_out;
wire _guard14568 = early_reset_static_par0_go_out;
wire _guard14569 = early_reset_static_par0_go_out;
wire _guard14570 = early_reset_static_par0_go_out;
wire _guard14571 = early_reset_static_par0_go_out;
wire _guard14572 = early_reset_static_par0_go_out;
wire _guard14573 = ~_guard0;
wire _guard14574 = early_reset_static_par0_go_out;
wire _guard14575 = _guard14573 & _guard14574;
wire _guard14576 = ~_guard0;
wire _guard14577 = early_reset_static_par0_go_out;
wire _guard14578 = _guard14576 & _guard14577;
wire _guard14579 = early_reset_static_par0_go_out;
wire _guard14580 = ~_guard0;
wire _guard14581 = early_reset_static_par0_go_out;
wire _guard14582 = _guard14580 & _guard14581;
wire _guard14583 = early_reset_static_par0_go_out;
wire _guard14584 = early_reset_static_par0_go_out;
wire _guard14585 = ~_guard0;
wire _guard14586 = early_reset_static_par0_go_out;
wire _guard14587 = _guard14585 & _guard14586;
wire _guard14588 = ~_guard0;
wire _guard14589 = early_reset_static_par0_go_out;
wire _guard14590 = _guard14588 & _guard14589;
wire _guard14591 = early_reset_static_par0_go_out;
wire _guard14592 = ~_guard0;
wire _guard14593 = early_reset_static_par0_go_out;
wire _guard14594 = _guard14592 & _guard14593;
wire _guard14595 = early_reset_static_par0_go_out;
wire _guard14596 = ~_guard0;
wire _guard14597 = early_reset_static_par0_go_out;
wire _guard14598 = _guard14596 & _guard14597;
wire _guard14599 = early_reset_static_par0_go_out;
wire _guard14600 = early_reset_static_par0_go_out;
wire _guard14601 = ~_guard0;
wire _guard14602 = early_reset_static_par0_go_out;
wire _guard14603 = _guard14601 & _guard14602;
wire _guard14604 = early_reset_static_par0_go_out;
wire _guard14605 = ~_guard0;
wire _guard14606 = early_reset_static_par0_go_out;
wire _guard14607 = _guard14605 & _guard14606;
wire _guard14608 = early_reset_static_par0_go_out;
wire _guard14609 = early_reset_static_par0_go_out;
wire _guard14610 = ~_guard0;
wire _guard14611 = early_reset_static_par0_go_out;
wire _guard14612 = _guard14610 & _guard14611;
wire _guard14613 = early_reset_static_par0_go_out;
wire _guard14614 = early_reset_static_par0_go_out;
wire _guard14615 = early_reset_static_par0_go_out;
wire _guard14616 = early_reset_static_par0_go_out;
wire _guard14617 = early_reset_static_par0_go_out;
wire _guard14618 = early_reset_static_par0_go_out;
wire _guard14619 = ~_guard0;
wire _guard14620 = early_reset_static_par0_go_out;
wire _guard14621 = _guard14619 & _guard14620;
wire _guard14622 = early_reset_static_par0_go_out;
wire _guard14623 = early_reset_static_par0_go_out;
wire _guard14624 = early_reset_static_par0_go_out;
wire _guard14625 = ~_guard0;
wire _guard14626 = early_reset_static_par0_go_out;
wire _guard14627 = _guard14625 & _guard14626;
wire _guard14628 = early_reset_static_par0_go_out;
wire _guard14629 = early_reset_static_par0_go_out;
wire _guard14630 = early_reset_static_par0_go_out;
wire _guard14631 = ~_guard0;
wire _guard14632 = early_reset_static_par0_go_out;
wire _guard14633 = _guard14631 & _guard14632;
wire _guard14634 = early_reset_static_par0_go_out;
wire _guard14635 = early_reset_static_par0_go_out;
wire _guard14636 = early_reset_static_par0_go_out;
wire _guard14637 = early_reset_static_par0_go_out;
wire _guard14638 = early_reset_static_par0_go_out;
wire _guard14639 = early_reset_static_par0_go_out;
wire _guard14640 = early_reset_static_par0_go_out;
wire _guard14641 = early_reset_static_par0_go_out;
wire _guard14642 = early_reset_static_par0_go_out;
wire _guard14643 = early_reset_static_par0_go_out;
wire _guard14644 = ~_guard0;
wire _guard14645 = early_reset_static_par0_go_out;
wire _guard14646 = _guard14644 & _guard14645;
wire _guard14647 = early_reset_static_par0_go_out;
wire _guard14648 = early_reset_static_par0_go_out;
wire _guard14649 = ~_guard0;
wire _guard14650 = early_reset_static_par0_go_out;
wire _guard14651 = _guard14649 & _guard14650;
wire _guard14652 = early_reset_static_par0_go_out;
wire _guard14653 = early_reset_static_par0_go_out;
wire _guard14654 = early_reset_static_par0_go_out;
wire _guard14655 = early_reset_static_par0_go_out;
wire _guard14656 = early_reset_static_par0_go_out;
wire _guard14657 = early_reset_static_par0_go_out;
wire _guard14658 = early_reset_static_par0_go_out;
wire _guard14659 = early_reset_static_par0_go_out;
wire _guard14660 = early_reset_static_par0_go_out;
wire _guard14661 = early_reset_static_par0_go_out;
wire _guard14662 = early_reset_static_par0_go_out;
wire _guard14663 = early_reset_static_par0_go_out;
wire _guard14664 = early_reset_static_par0_go_out;
wire _guard14665 = ~_guard0;
wire _guard14666 = early_reset_static_par0_go_out;
wire _guard14667 = _guard14665 & _guard14666;
wire _guard14668 = early_reset_static_par0_go_out;
wire _guard14669 = ~_guard0;
wire _guard14670 = early_reset_static_par0_go_out;
wire _guard14671 = _guard14669 & _guard14670;
wire _guard14672 = early_reset_static_par0_go_out;
wire _guard14673 = early_reset_static_par0_go_out;
wire _guard14674 = early_reset_static_par0_go_out;
wire _guard14675 = ~_guard0;
wire _guard14676 = early_reset_static_par0_go_out;
wire _guard14677 = _guard14675 & _guard14676;
wire _guard14678 = early_reset_static_par0_go_out;
wire _guard14679 = early_reset_static_par0_go_out;
wire _guard14680 = ~_guard0;
wire _guard14681 = early_reset_static_par0_go_out;
wire _guard14682 = _guard14680 & _guard14681;
wire _guard14683 = early_reset_static_par0_go_out;
wire _guard14684 = early_reset_static_par0_go_out;
wire _guard14685 = early_reset_static_par0_go_out;
wire _guard14686 = early_reset_static_par0_go_out;
wire _guard14687 = early_reset_static_par0_go_out;
wire _guard14688 = early_reset_static_par0_go_out;
wire _guard14689 = ~_guard0;
wire _guard14690 = early_reset_static_par0_go_out;
wire _guard14691 = _guard14689 & _guard14690;
wire _guard14692 = early_reset_static_par0_go_out;
wire _guard14693 = early_reset_static_par0_go_out;
wire _guard14694 = early_reset_static_par0_go_out;
wire _guard14695 = early_reset_static_par0_go_out;
wire _guard14696 = early_reset_static_par0_go_out;
wire _guard14697 = ~_guard0;
wire _guard14698 = early_reset_static_par0_go_out;
wire _guard14699 = _guard14697 & _guard14698;
wire _guard14700 = early_reset_static_par0_go_out;
wire _guard14701 = early_reset_static_par0_go_out;
wire _guard14702 = ~_guard0;
wire _guard14703 = early_reset_static_par0_go_out;
wire _guard14704 = _guard14702 & _guard14703;
wire _guard14705 = early_reset_static_par0_go_out;
wire _guard14706 = early_reset_static_par0_go_out;
wire _guard14707 = ~_guard0;
wire _guard14708 = early_reset_static_par0_go_out;
wire _guard14709 = _guard14707 & _guard14708;
wire _guard14710 = ~_guard0;
wire _guard14711 = early_reset_static_par0_go_out;
wire _guard14712 = _guard14710 & _guard14711;
wire _guard14713 = early_reset_static_par0_go_out;
wire _guard14714 = ~_guard0;
wire _guard14715 = early_reset_static_par0_go_out;
wire _guard14716 = _guard14714 & _guard14715;
wire _guard14717 = early_reset_static_par0_go_out;
wire _guard14718 = early_reset_static_par0_go_out;
wire _guard14719 = early_reset_static_par0_go_out;
wire _guard14720 = ~_guard0;
wire _guard14721 = early_reset_static_par0_go_out;
wire _guard14722 = _guard14720 & _guard14721;
wire _guard14723 = early_reset_static_par0_go_out;
wire _guard14724 = early_reset_static_par0_go_out;
wire _guard14725 = early_reset_static_par0_go_out;
wire _guard14726 = ~_guard0;
wire _guard14727 = early_reset_static_par0_go_out;
wire _guard14728 = _guard14726 & _guard14727;
wire _guard14729 = early_reset_static_par0_go_out;
wire _guard14730 = early_reset_static_par0_go_out;
wire _guard14731 = early_reset_static_par0_go_out;
wire _guard14732 = early_reset_static_par0_go_out;
wire _guard14733 = early_reset_static_par0_go_out;
wire _guard14734 = ~_guard0;
wire _guard14735 = early_reset_static_par0_go_out;
wire _guard14736 = _guard14734 & _guard14735;
wire _guard14737 = early_reset_static_par0_go_out;
wire _guard14738 = ~_guard0;
wire _guard14739 = early_reset_static_par0_go_out;
wire _guard14740 = _guard14738 & _guard14739;
wire _guard14741 = early_reset_static_par0_go_out;
wire _guard14742 = early_reset_static_par0_go_out;
wire _guard14743 = early_reset_static_par0_go_out;
wire _guard14744 = ~_guard0;
wire _guard14745 = early_reset_static_par0_go_out;
wire _guard14746 = _guard14744 & _guard14745;
wire _guard14747 = early_reset_static_par0_go_out;
wire _guard14748 = early_reset_static_par0_go_out;
wire _guard14749 = early_reset_static_par0_go_out;
wire _guard14750 = early_reset_static_par0_go_out;
wire _guard14751 = early_reset_static_par0_go_out;
wire _guard14752 = ~_guard0;
wire _guard14753 = early_reset_static_par0_go_out;
wire _guard14754 = _guard14752 & _guard14753;
wire _guard14755 = early_reset_static_par0_go_out;
wire _guard14756 = early_reset_static_par0_go_out;
wire _guard14757 = early_reset_static_par0_go_out;
wire _guard14758 = early_reset_static_par0_go_out;
wire _guard14759 = ~_guard0;
wire _guard14760 = early_reset_static_par0_go_out;
wire _guard14761 = _guard14759 & _guard14760;
wire _guard14762 = early_reset_static_par0_go_out;
wire _guard14763 = early_reset_static_par0_go_out;
wire _guard14764 = early_reset_static_par0_go_out;
wire _guard14765 = early_reset_static_par0_go_out;
wire _guard14766 = early_reset_static_par0_go_out;
wire _guard14767 = early_reset_static_par0_go_out;
wire _guard14768 = ~_guard0;
wire _guard14769 = early_reset_static_par0_go_out;
wire _guard14770 = _guard14768 & _guard14769;
wire _guard14771 = early_reset_static_par0_go_out;
wire _guard14772 = early_reset_static_par0_go_out;
wire _guard14773 = early_reset_static_par0_go_out;
wire _guard14774 = early_reset_static_par0_go_out;
wire _guard14775 = early_reset_static_par0_go_out;
wire _guard14776 = early_reset_static_par0_go_out;
wire _guard14777 = early_reset_static_par0_go_out;
wire _guard14778 = early_reset_static_par0_go_out;
wire _guard14779 = ~_guard0;
wire _guard14780 = early_reset_static_par0_go_out;
wire _guard14781 = _guard14779 & _guard14780;
wire _guard14782 = ~_guard0;
wire _guard14783 = early_reset_static_par0_go_out;
wire _guard14784 = _guard14782 & _guard14783;
wire _guard14785 = early_reset_static_par0_go_out;
wire _guard14786 = ~_guard0;
wire _guard14787 = early_reset_static_par0_go_out;
wire _guard14788 = _guard14786 & _guard14787;
wire _guard14789 = early_reset_static_par0_go_out;
wire _guard14790 = ~_guard0;
wire _guard14791 = early_reset_static_par0_go_out;
wire _guard14792 = _guard14790 & _guard14791;
wire _guard14793 = early_reset_static_par0_go_out;
wire _guard14794 = early_reset_static_par0_go_out;
wire _guard14795 = early_reset_static_par0_go_out;
wire _guard14796 = early_reset_static_par0_go_out;
wire _guard14797 = early_reset_static_par0_go_out;
wire _guard14798 = early_reset_static_par0_go_out;
wire _guard14799 = early_reset_static_par0_go_out;
wire _guard14800 = early_reset_static_par0_go_out;
wire _guard14801 = ~_guard0;
wire _guard14802 = early_reset_static_par0_go_out;
wire _guard14803 = _guard14801 & _guard14802;
wire _guard14804 = early_reset_static_par0_go_out;
wire _guard14805 = early_reset_static_par0_go_out;
wire _guard14806 = ~_guard0;
wire _guard14807 = early_reset_static_par0_go_out;
wire _guard14808 = _guard14806 & _guard14807;
wire _guard14809 = early_reset_static_par0_go_out;
wire _guard14810 = early_reset_static_par0_go_out;
wire _guard14811 = early_reset_static_par0_go_out;
wire _guard14812 = early_reset_static_par0_go_out;
wire _guard14813 = early_reset_static_par0_go_out;
wire _guard14814 = early_reset_static_par0_go_out;
wire _guard14815 = early_reset_static_par0_go_out;
wire _guard14816 = early_reset_static_par0_go_out;
wire _guard14817 = ~_guard0;
wire _guard14818 = early_reset_static_par0_go_out;
wire _guard14819 = _guard14817 & _guard14818;
wire _guard14820 = early_reset_static_par0_go_out;
wire _guard14821 = early_reset_static_par0_go_out;
wire _guard14822 = early_reset_static_par0_go_out;
wire _guard14823 = ~_guard0;
wire _guard14824 = early_reset_static_par0_go_out;
wire _guard14825 = _guard14823 & _guard14824;
wire _guard14826 = early_reset_static_par0_go_out;
wire _guard14827 = ~_guard0;
wire _guard14828 = early_reset_static_par0_go_out;
wire _guard14829 = _guard14827 & _guard14828;
wire _guard14830 = early_reset_static_par0_go_out;
wire _guard14831 = early_reset_static_par0_go_out;
wire _guard14832 = early_reset_static_par0_go_out;
wire _guard14833 = ~_guard0;
wire _guard14834 = early_reset_static_par0_go_out;
wire _guard14835 = _guard14833 & _guard14834;
wire _guard14836 = early_reset_static_par0_go_out;
wire _guard14837 = early_reset_static_par0_go_out;
wire _guard14838 = early_reset_static_par0_go_out;
wire _guard14839 = early_reset_static_par0_go_out;
wire _guard14840 = ~_guard0;
wire _guard14841 = early_reset_static_par0_go_out;
wire _guard14842 = _guard14840 & _guard14841;
wire _guard14843 = early_reset_static_par0_go_out;
wire _guard14844 = ~_guard0;
wire _guard14845 = early_reset_static_par0_go_out;
wire _guard14846 = _guard14844 & _guard14845;
wire _guard14847 = early_reset_static_par0_go_out;
wire _guard14848 = early_reset_static_par0_go_out;
wire _guard14849 = early_reset_static_par0_go_out;
wire _guard14850 = early_reset_static_seq_go_out;
wire _guard14851 = fsm0_out != 6'd52;
wire _guard14852 = early_reset_static_seq_go_out;
wire _guard14853 = _guard14851 & _guard14852;
wire _guard14854 = fsm0_out == 6'd52;
wire _guard14855 = early_reset_static_seq_go_out;
wire _guard14856 = _guard14854 & _guard14855;
wire _guard14857 = cond_wire41_out;
wire _guard14858 = early_reset_static_par0_go_out;
wire _guard14859 = _guard14857 & _guard14858;
wire _guard14860 = cond_wire41_out;
wire _guard14861 = early_reset_static_par0_go_out;
wire _guard14862 = _guard14860 & _guard14861;
wire _guard14863 = cond_wire102_out;
wire _guard14864 = early_reset_static_par0_go_out;
wire _guard14865 = _guard14863 & _guard14864;
wire _guard14866 = cond_wire100_out;
wire _guard14867 = early_reset_static_par0_go_out;
wire _guard14868 = _guard14866 & _guard14867;
wire _guard14869 = fsm_out == 1'd0;
wire _guard14870 = cond_wire100_out;
wire _guard14871 = _guard14869 & _guard14870;
wire _guard14872 = fsm_out == 1'd0;
wire _guard14873 = _guard14871 & _guard14872;
wire _guard14874 = fsm_out == 1'd0;
wire _guard14875 = cond_wire102_out;
wire _guard14876 = _guard14874 & _guard14875;
wire _guard14877 = fsm_out == 1'd0;
wire _guard14878 = _guard14876 & _guard14877;
wire _guard14879 = _guard14873 | _guard14878;
wire _guard14880 = early_reset_static_par0_go_out;
wire _guard14881 = _guard14879 & _guard14880;
wire _guard14882 = fsm_out == 1'd0;
wire _guard14883 = cond_wire100_out;
wire _guard14884 = _guard14882 & _guard14883;
wire _guard14885 = fsm_out == 1'd0;
wire _guard14886 = _guard14884 & _guard14885;
wire _guard14887 = fsm_out == 1'd0;
wire _guard14888 = cond_wire102_out;
wire _guard14889 = _guard14887 & _guard14888;
wire _guard14890 = fsm_out == 1'd0;
wire _guard14891 = _guard14889 & _guard14890;
wire _guard14892 = _guard14886 | _guard14891;
wire _guard14893 = early_reset_static_par0_go_out;
wire _guard14894 = _guard14892 & _guard14893;
wire _guard14895 = fsm_out == 1'd0;
wire _guard14896 = cond_wire100_out;
wire _guard14897 = _guard14895 & _guard14896;
wire _guard14898 = fsm_out == 1'd0;
wire _guard14899 = _guard14897 & _guard14898;
wire _guard14900 = fsm_out == 1'd0;
wire _guard14901 = cond_wire102_out;
wire _guard14902 = _guard14900 & _guard14901;
wire _guard14903 = fsm_out == 1'd0;
wire _guard14904 = _guard14902 & _guard14903;
wire _guard14905 = _guard14899 | _guard14904;
wire _guard14906 = early_reset_static_par0_go_out;
wire _guard14907 = _guard14905 & _guard14906;
wire _guard14908 = cond_wire31_out;
wire _guard14909 = early_reset_static_par0_go_out;
wire _guard14910 = _guard14908 & _guard14909;
wire _guard14911 = cond_wire31_out;
wire _guard14912 = early_reset_static_par0_go_out;
wire _guard14913 = _guard14911 & _guard14912;
wire _guard14914 = cond_wire117_out;
wire _guard14915 = early_reset_static_par0_go_out;
wire _guard14916 = _guard14914 & _guard14915;
wire _guard14917 = cond_wire117_out;
wire _guard14918 = early_reset_static_par0_go_out;
wire _guard14919 = _guard14917 & _guard14918;
wire _guard14920 = cond_wire56_out;
wire _guard14921 = early_reset_static_par0_go_out;
wire _guard14922 = _guard14920 & _guard14921;
wire _guard14923 = cond_wire56_out;
wire _guard14924 = early_reset_static_par0_go_out;
wire _guard14925 = _guard14923 & _guard14924;
wire _guard14926 = cond_wire81_out;
wire _guard14927 = early_reset_static_par0_go_out;
wire _guard14928 = _guard14926 & _guard14927;
wire _guard14929 = cond_wire81_out;
wire _guard14930 = early_reset_static_par0_go_out;
wire _guard14931 = _guard14929 & _guard14930;
wire _guard14932 = cond_wire190_out;
wire _guard14933 = early_reset_static_par0_go_out;
wire _guard14934 = _guard14932 & _guard14933;
wire _guard14935 = cond_wire190_out;
wire _guard14936 = early_reset_static_par0_go_out;
wire _guard14937 = _guard14935 & _guard14936;
wire _guard14938 = cond_wire146_out;
wire _guard14939 = early_reset_static_par0_go_out;
wire _guard14940 = _guard14938 & _guard14939;
wire _guard14941 = cond_wire146_out;
wire _guard14942 = early_reset_static_par0_go_out;
wire _guard14943 = _guard14941 & _guard14942;
wire _guard14944 = cond_wire150_out;
wire _guard14945 = early_reset_static_par0_go_out;
wire _guard14946 = _guard14944 & _guard14945;
wire _guard14947 = cond_wire150_out;
wire _guard14948 = early_reset_static_par0_go_out;
wire _guard14949 = _guard14947 & _guard14948;
wire _guard14950 = cond_wire182_out;
wire _guard14951 = early_reset_static_par0_go_out;
wire _guard14952 = _guard14950 & _guard14951;
wire _guard14953 = cond_wire182_out;
wire _guard14954 = early_reset_static_par0_go_out;
wire _guard14955 = _guard14953 & _guard14954;
wire _guard14956 = cond_wire186_out;
wire _guard14957 = early_reset_static_par0_go_out;
wire _guard14958 = _guard14956 & _guard14957;
wire _guard14959 = cond_wire186_out;
wire _guard14960 = early_reset_static_par0_go_out;
wire _guard14961 = _guard14959 & _guard14960;
wire _guard14962 = cond_wire206_out;
wire _guard14963 = early_reset_static_par0_go_out;
wire _guard14964 = _guard14962 & _guard14963;
wire _guard14965 = cond_wire206_out;
wire _guard14966 = early_reset_static_par0_go_out;
wire _guard14967 = _guard14965 & _guard14966;
wire _guard14968 = cond_wire301_out;
wire _guard14969 = early_reset_static_par0_go_out;
wire _guard14970 = _guard14968 & _guard14969;
wire _guard14971 = cond_wire299_out;
wire _guard14972 = early_reset_static_par0_go_out;
wire _guard14973 = _guard14971 & _guard14972;
wire _guard14974 = fsm_out == 1'd0;
wire _guard14975 = cond_wire299_out;
wire _guard14976 = _guard14974 & _guard14975;
wire _guard14977 = fsm_out == 1'd0;
wire _guard14978 = _guard14976 & _guard14977;
wire _guard14979 = fsm_out == 1'd0;
wire _guard14980 = cond_wire301_out;
wire _guard14981 = _guard14979 & _guard14980;
wire _guard14982 = fsm_out == 1'd0;
wire _guard14983 = _guard14981 & _guard14982;
wire _guard14984 = _guard14978 | _guard14983;
wire _guard14985 = early_reset_static_par0_go_out;
wire _guard14986 = _guard14984 & _guard14985;
wire _guard14987 = fsm_out == 1'd0;
wire _guard14988 = cond_wire299_out;
wire _guard14989 = _guard14987 & _guard14988;
wire _guard14990 = fsm_out == 1'd0;
wire _guard14991 = _guard14989 & _guard14990;
wire _guard14992 = fsm_out == 1'd0;
wire _guard14993 = cond_wire301_out;
wire _guard14994 = _guard14992 & _guard14993;
wire _guard14995 = fsm_out == 1'd0;
wire _guard14996 = _guard14994 & _guard14995;
wire _guard14997 = _guard14991 | _guard14996;
wire _guard14998 = early_reset_static_par0_go_out;
wire _guard14999 = _guard14997 & _guard14998;
wire _guard15000 = fsm_out == 1'd0;
wire _guard15001 = cond_wire299_out;
wire _guard15002 = _guard15000 & _guard15001;
wire _guard15003 = fsm_out == 1'd0;
wire _guard15004 = _guard15002 & _guard15003;
wire _guard15005 = fsm_out == 1'd0;
wire _guard15006 = cond_wire301_out;
wire _guard15007 = _guard15005 & _guard15006;
wire _guard15008 = fsm_out == 1'd0;
wire _guard15009 = _guard15007 & _guard15008;
wire _guard15010 = _guard15004 | _guard15009;
wire _guard15011 = early_reset_static_par0_go_out;
wire _guard15012 = _guard15010 & _guard15011;
wire _guard15013 = cond_wire312_out;
wire _guard15014 = early_reset_static_par0_go_out;
wire _guard15015 = _guard15013 & _guard15014;
wire _guard15016 = cond_wire312_out;
wire _guard15017 = early_reset_static_par0_go_out;
wire _guard15018 = _guard15016 & _guard15017;
wire _guard15019 = cond_wire321_out;
wire _guard15020 = early_reset_static_par0_go_out;
wire _guard15021 = _guard15019 & _guard15020;
wire _guard15022 = cond_wire319_out;
wire _guard15023 = early_reset_static_par0_go_out;
wire _guard15024 = _guard15022 & _guard15023;
wire _guard15025 = fsm_out == 1'd0;
wire _guard15026 = cond_wire319_out;
wire _guard15027 = _guard15025 & _guard15026;
wire _guard15028 = fsm_out == 1'd0;
wire _guard15029 = _guard15027 & _guard15028;
wire _guard15030 = fsm_out == 1'd0;
wire _guard15031 = cond_wire321_out;
wire _guard15032 = _guard15030 & _guard15031;
wire _guard15033 = fsm_out == 1'd0;
wire _guard15034 = _guard15032 & _guard15033;
wire _guard15035 = _guard15029 | _guard15034;
wire _guard15036 = early_reset_static_par0_go_out;
wire _guard15037 = _guard15035 & _guard15036;
wire _guard15038 = fsm_out == 1'd0;
wire _guard15039 = cond_wire319_out;
wire _guard15040 = _guard15038 & _guard15039;
wire _guard15041 = fsm_out == 1'd0;
wire _guard15042 = _guard15040 & _guard15041;
wire _guard15043 = fsm_out == 1'd0;
wire _guard15044 = cond_wire321_out;
wire _guard15045 = _guard15043 & _guard15044;
wire _guard15046 = fsm_out == 1'd0;
wire _guard15047 = _guard15045 & _guard15046;
wire _guard15048 = _guard15042 | _guard15047;
wire _guard15049 = early_reset_static_par0_go_out;
wire _guard15050 = _guard15048 & _guard15049;
wire _guard15051 = fsm_out == 1'd0;
wire _guard15052 = cond_wire319_out;
wire _guard15053 = _guard15051 & _guard15052;
wire _guard15054 = fsm_out == 1'd0;
wire _guard15055 = _guard15053 & _guard15054;
wire _guard15056 = fsm_out == 1'd0;
wire _guard15057 = cond_wire321_out;
wire _guard15058 = _guard15056 & _guard15057;
wire _guard15059 = fsm_out == 1'd0;
wire _guard15060 = _guard15058 & _guard15059;
wire _guard15061 = _guard15055 | _guard15060;
wire _guard15062 = early_reset_static_par0_go_out;
wire _guard15063 = _guard15061 & _guard15062;
wire _guard15064 = cond_wire284_out;
wire _guard15065 = early_reset_static_par0_go_out;
wire _guard15066 = _guard15064 & _guard15065;
wire _guard15067 = cond_wire284_out;
wire _guard15068 = early_reset_static_par0_go_out;
wire _guard15069 = _guard15067 & _guard15068;
wire _guard15070 = cond_wire292_out;
wire _guard15071 = early_reset_static_par0_go_out;
wire _guard15072 = _guard15070 & _guard15071;
wire _guard15073 = cond_wire292_out;
wire _guard15074 = early_reset_static_par0_go_out;
wire _guard15075 = _guard15073 & _guard15074;
wire _guard15076 = cond_wire377_out;
wire _guard15077 = early_reset_static_par0_go_out;
wire _guard15078 = _guard15076 & _guard15077;
wire _guard15079 = cond_wire377_out;
wire _guard15080 = early_reset_static_par0_go_out;
wire _guard15081 = _guard15079 & _guard15080;
wire _guard15082 = cond_wire328_out;
wire _guard15083 = early_reset_static_par0_go_out;
wire _guard15084 = _guard15082 & _guard15083;
wire _guard15085 = cond_wire328_out;
wire _guard15086 = early_reset_static_par0_go_out;
wire _guard15087 = _guard15085 & _guard15086;
wire _guard15088 = cond_wire397_out;
wire _guard15089 = early_reset_static_par0_go_out;
wire _guard15090 = _guard15088 & _guard15089;
wire _guard15091 = cond_wire397_out;
wire _guard15092 = early_reset_static_par0_go_out;
wire _guard15093 = _guard15091 & _guard15092;
wire _guard15094 = cond_wire458_out;
wire _guard15095 = early_reset_static_par0_go_out;
wire _guard15096 = _guard15094 & _guard15095;
wire _guard15097 = cond_wire458_out;
wire _guard15098 = early_reset_static_par0_go_out;
wire _guard15099 = _guard15097 & _guard15098;
wire _guard15100 = cond_wire462_out;
wire _guard15101 = early_reset_static_par0_go_out;
wire _guard15102 = _guard15100 & _guard15101;
wire _guard15103 = cond_wire462_out;
wire _guard15104 = early_reset_static_par0_go_out;
wire _guard15105 = _guard15103 & _guard15104;
wire _guard15106 = cond_wire495_out;
wire _guard15107 = early_reset_static_par0_go_out;
wire _guard15108 = _guard15106 & _guard15107;
wire _guard15109 = cond_wire495_out;
wire _guard15110 = early_reset_static_par0_go_out;
wire _guard15111 = _guard15109 & _guard15110;
wire _guard15112 = cond_wire568_out;
wire _guard15113 = early_reset_static_par0_go_out;
wire _guard15114 = _guard15112 & _guard15113;
wire _guard15115 = cond_wire568_out;
wire _guard15116 = early_reset_static_par0_go_out;
wire _guard15117 = _guard15115 & _guard15116;
wire _guard15118 = cond_wire580_out;
wire _guard15119 = early_reset_static_par0_go_out;
wire _guard15120 = _guard15118 & _guard15119;
wire _guard15121 = cond_wire580_out;
wire _guard15122 = early_reset_static_par0_go_out;
wire _guard15123 = _guard15121 & _guard15122;
wire _guard15124 = cond_wire523_out;
wire _guard15125 = early_reset_static_par0_go_out;
wire _guard15126 = _guard15124 & _guard15125;
wire _guard15127 = cond_wire523_out;
wire _guard15128 = early_reset_static_par0_go_out;
wire _guard15129 = _guard15127 & _guard15128;
wire _guard15130 = cond_wire642_out;
wire _guard15131 = early_reset_static_par0_go_out;
wire _guard15132 = _guard15130 & _guard15131;
wire _guard15133 = cond_wire640_out;
wire _guard15134 = early_reset_static_par0_go_out;
wire _guard15135 = _guard15133 & _guard15134;
wire _guard15136 = fsm_out == 1'd0;
wire _guard15137 = cond_wire640_out;
wire _guard15138 = _guard15136 & _guard15137;
wire _guard15139 = fsm_out == 1'd0;
wire _guard15140 = _guard15138 & _guard15139;
wire _guard15141 = fsm_out == 1'd0;
wire _guard15142 = cond_wire642_out;
wire _guard15143 = _guard15141 & _guard15142;
wire _guard15144 = fsm_out == 1'd0;
wire _guard15145 = _guard15143 & _guard15144;
wire _guard15146 = _guard15140 | _guard15145;
wire _guard15147 = early_reset_static_par0_go_out;
wire _guard15148 = _guard15146 & _guard15147;
wire _guard15149 = fsm_out == 1'd0;
wire _guard15150 = cond_wire640_out;
wire _guard15151 = _guard15149 & _guard15150;
wire _guard15152 = fsm_out == 1'd0;
wire _guard15153 = _guard15151 & _guard15152;
wire _guard15154 = fsm_out == 1'd0;
wire _guard15155 = cond_wire642_out;
wire _guard15156 = _guard15154 & _guard15155;
wire _guard15157 = fsm_out == 1'd0;
wire _guard15158 = _guard15156 & _guard15157;
wire _guard15159 = _guard15153 | _guard15158;
wire _guard15160 = early_reset_static_par0_go_out;
wire _guard15161 = _guard15159 & _guard15160;
wire _guard15162 = fsm_out == 1'd0;
wire _guard15163 = cond_wire640_out;
wire _guard15164 = _guard15162 & _guard15163;
wire _guard15165 = fsm_out == 1'd0;
wire _guard15166 = _guard15164 & _guard15165;
wire _guard15167 = fsm_out == 1'd0;
wire _guard15168 = cond_wire642_out;
wire _guard15169 = _guard15167 & _guard15168;
wire _guard15170 = fsm_out == 1'd0;
wire _guard15171 = _guard15169 & _guard15170;
wire _guard15172 = _guard15166 | _guard15171;
wire _guard15173 = early_reset_static_par0_go_out;
wire _guard15174 = _guard15172 & _guard15173;
wire _guard15175 = cond_wire650_out;
wire _guard15176 = early_reset_static_par0_go_out;
wire _guard15177 = _guard15175 & _guard15176;
wire _guard15178 = cond_wire648_out;
wire _guard15179 = early_reset_static_par0_go_out;
wire _guard15180 = _guard15178 & _guard15179;
wire _guard15181 = fsm_out == 1'd0;
wire _guard15182 = cond_wire648_out;
wire _guard15183 = _guard15181 & _guard15182;
wire _guard15184 = fsm_out == 1'd0;
wire _guard15185 = _guard15183 & _guard15184;
wire _guard15186 = fsm_out == 1'd0;
wire _guard15187 = cond_wire650_out;
wire _guard15188 = _guard15186 & _guard15187;
wire _guard15189 = fsm_out == 1'd0;
wire _guard15190 = _guard15188 & _guard15189;
wire _guard15191 = _guard15185 | _guard15190;
wire _guard15192 = early_reset_static_par0_go_out;
wire _guard15193 = _guard15191 & _guard15192;
wire _guard15194 = fsm_out == 1'd0;
wire _guard15195 = cond_wire648_out;
wire _guard15196 = _guard15194 & _guard15195;
wire _guard15197 = fsm_out == 1'd0;
wire _guard15198 = _guard15196 & _guard15197;
wire _guard15199 = fsm_out == 1'd0;
wire _guard15200 = cond_wire650_out;
wire _guard15201 = _guard15199 & _guard15200;
wire _guard15202 = fsm_out == 1'd0;
wire _guard15203 = _guard15201 & _guard15202;
wire _guard15204 = _guard15198 | _guard15203;
wire _guard15205 = early_reset_static_par0_go_out;
wire _guard15206 = _guard15204 & _guard15205;
wire _guard15207 = fsm_out == 1'd0;
wire _guard15208 = cond_wire648_out;
wire _guard15209 = _guard15207 & _guard15208;
wire _guard15210 = fsm_out == 1'd0;
wire _guard15211 = _guard15209 & _guard15210;
wire _guard15212 = fsm_out == 1'd0;
wire _guard15213 = cond_wire650_out;
wire _guard15214 = _guard15212 & _guard15213;
wire _guard15215 = fsm_out == 1'd0;
wire _guard15216 = _guard15214 & _guard15215;
wire _guard15217 = _guard15211 | _guard15216;
wire _guard15218 = early_reset_static_par0_go_out;
wire _guard15219 = _guard15217 & _guard15218;
wire _guard15220 = cond_wire605_out;
wire _guard15221 = early_reset_static_par0_go_out;
wire _guard15222 = _guard15220 & _guard15221;
wire _guard15223 = cond_wire605_out;
wire _guard15224 = early_reset_static_par0_go_out;
wire _guard15225 = _guard15223 & _guard15224;
wire _guard15226 = cond_wire723_out;
wire _guard15227 = early_reset_static_par0_go_out;
wire _guard15228 = _guard15226 & _guard15227;
wire _guard15229 = cond_wire721_out;
wire _guard15230 = early_reset_static_par0_go_out;
wire _guard15231 = _guard15229 & _guard15230;
wire _guard15232 = fsm_out == 1'd0;
wire _guard15233 = cond_wire721_out;
wire _guard15234 = _guard15232 & _guard15233;
wire _guard15235 = fsm_out == 1'd0;
wire _guard15236 = _guard15234 & _guard15235;
wire _guard15237 = fsm_out == 1'd0;
wire _guard15238 = cond_wire723_out;
wire _guard15239 = _guard15237 & _guard15238;
wire _guard15240 = fsm_out == 1'd0;
wire _guard15241 = _guard15239 & _guard15240;
wire _guard15242 = _guard15236 | _guard15241;
wire _guard15243 = early_reset_static_par0_go_out;
wire _guard15244 = _guard15242 & _guard15243;
wire _guard15245 = fsm_out == 1'd0;
wire _guard15246 = cond_wire721_out;
wire _guard15247 = _guard15245 & _guard15246;
wire _guard15248 = fsm_out == 1'd0;
wire _guard15249 = _guard15247 & _guard15248;
wire _guard15250 = fsm_out == 1'd0;
wire _guard15251 = cond_wire723_out;
wire _guard15252 = _guard15250 & _guard15251;
wire _guard15253 = fsm_out == 1'd0;
wire _guard15254 = _guard15252 & _guard15253;
wire _guard15255 = _guard15249 | _guard15254;
wire _guard15256 = early_reset_static_par0_go_out;
wire _guard15257 = _guard15255 & _guard15256;
wire _guard15258 = fsm_out == 1'd0;
wire _guard15259 = cond_wire721_out;
wire _guard15260 = _guard15258 & _guard15259;
wire _guard15261 = fsm_out == 1'd0;
wire _guard15262 = _guard15260 & _guard15261;
wire _guard15263 = fsm_out == 1'd0;
wire _guard15264 = cond_wire723_out;
wire _guard15265 = _guard15263 & _guard15264;
wire _guard15266 = fsm_out == 1'd0;
wire _guard15267 = _guard15265 & _guard15266;
wire _guard15268 = _guard15262 | _guard15267;
wire _guard15269 = early_reset_static_par0_go_out;
wire _guard15270 = _guard15268 & _guard15269;
wire _guard15271 = cond_wire722_out;
wire _guard15272 = early_reset_static_par0_go_out;
wire _guard15273 = _guard15271 & _guard15272;
wire _guard15274 = cond_wire722_out;
wire _guard15275 = early_reset_static_par0_go_out;
wire _guard15276 = _guard15274 & _guard15275;
wire _guard15277 = cond_wire740_out;
wire _guard15278 = early_reset_static_par0_go_out;
wire _guard15279 = _guard15277 & _guard15278;
wire _guard15280 = cond_wire738_out;
wire _guard15281 = early_reset_static_par0_go_out;
wire _guard15282 = _guard15280 & _guard15281;
wire _guard15283 = fsm_out == 1'd0;
wire _guard15284 = cond_wire738_out;
wire _guard15285 = _guard15283 & _guard15284;
wire _guard15286 = fsm_out == 1'd0;
wire _guard15287 = _guard15285 & _guard15286;
wire _guard15288 = fsm_out == 1'd0;
wire _guard15289 = cond_wire740_out;
wire _guard15290 = _guard15288 & _guard15289;
wire _guard15291 = fsm_out == 1'd0;
wire _guard15292 = _guard15290 & _guard15291;
wire _guard15293 = _guard15287 | _guard15292;
wire _guard15294 = early_reset_static_par0_go_out;
wire _guard15295 = _guard15293 & _guard15294;
wire _guard15296 = fsm_out == 1'd0;
wire _guard15297 = cond_wire738_out;
wire _guard15298 = _guard15296 & _guard15297;
wire _guard15299 = fsm_out == 1'd0;
wire _guard15300 = _guard15298 & _guard15299;
wire _guard15301 = fsm_out == 1'd0;
wire _guard15302 = cond_wire740_out;
wire _guard15303 = _guard15301 & _guard15302;
wire _guard15304 = fsm_out == 1'd0;
wire _guard15305 = _guard15303 & _guard15304;
wire _guard15306 = _guard15300 | _guard15305;
wire _guard15307 = early_reset_static_par0_go_out;
wire _guard15308 = _guard15306 & _guard15307;
wire _guard15309 = fsm_out == 1'd0;
wire _guard15310 = cond_wire738_out;
wire _guard15311 = _guard15309 & _guard15310;
wire _guard15312 = fsm_out == 1'd0;
wire _guard15313 = _guard15311 & _guard15312;
wire _guard15314 = fsm_out == 1'd0;
wire _guard15315 = cond_wire740_out;
wire _guard15316 = _guard15314 & _guard15315;
wire _guard15317 = fsm_out == 1'd0;
wire _guard15318 = _guard15316 & _guard15317;
wire _guard15319 = _guard15313 | _guard15318;
wire _guard15320 = early_reset_static_par0_go_out;
wire _guard15321 = _guard15319 & _guard15320;
wire _guard15322 = cond_wire674_out;
wire _guard15323 = early_reset_static_par0_go_out;
wire _guard15324 = _guard15322 & _guard15323;
wire _guard15325 = cond_wire674_out;
wire _guard15326 = early_reset_static_par0_go_out;
wire _guard15327 = _guard15325 & _guard15326;
wire _guard15328 = cond_wire744_out;
wire _guard15329 = early_reset_static_par0_go_out;
wire _guard15330 = _guard15328 & _guard15329;
wire _guard15331 = cond_wire742_out;
wire _guard15332 = early_reset_static_par0_go_out;
wire _guard15333 = _guard15331 & _guard15332;
wire _guard15334 = fsm_out == 1'd0;
wire _guard15335 = cond_wire742_out;
wire _guard15336 = _guard15334 & _guard15335;
wire _guard15337 = fsm_out == 1'd0;
wire _guard15338 = _guard15336 & _guard15337;
wire _guard15339 = fsm_out == 1'd0;
wire _guard15340 = cond_wire744_out;
wire _guard15341 = _guard15339 & _guard15340;
wire _guard15342 = fsm_out == 1'd0;
wire _guard15343 = _guard15341 & _guard15342;
wire _guard15344 = _guard15338 | _guard15343;
wire _guard15345 = early_reset_static_par0_go_out;
wire _guard15346 = _guard15344 & _guard15345;
wire _guard15347 = fsm_out == 1'd0;
wire _guard15348 = cond_wire742_out;
wire _guard15349 = _guard15347 & _guard15348;
wire _guard15350 = fsm_out == 1'd0;
wire _guard15351 = _guard15349 & _guard15350;
wire _guard15352 = fsm_out == 1'd0;
wire _guard15353 = cond_wire744_out;
wire _guard15354 = _guard15352 & _guard15353;
wire _guard15355 = fsm_out == 1'd0;
wire _guard15356 = _guard15354 & _guard15355;
wire _guard15357 = _guard15351 | _guard15356;
wire _guard15358 = early_reset_static_par0_go_out;
wire _guard15359 = _guard15357 & _guard15358;
wire _guard15360 = fsm_out == 1'd0;
wire _guard15361 = cond_wire742_out;
wire _guard15362 = _guard15360 & _guard15361;
wire _guard15363 = fsm_out == 1'd0;
wire _guard15364 = _guard15362 & _guard15363;
wire _guard15365 = fsm_out == 1'd0;
wire _guard15366 = cond_wire744_out;
wire _guard15367 = _guard15365 & _guard15366;
wire _guard15368 = fsm_out == 1'd0;
wire _guard15369 = _guard15367 & _guard15368;
wire _guard15370 = _guard15364 | _guard15369;
wire _guard15371 = early_reset_static_par0_go_out;
wire _guard15372 = _guard15370 & _guard15371;
wire _guard15373 = cond_wire690_out;
wire _guard15374 = early_reset_static_par0_go_out;
wire _guard15375 = _guard15373 & _guard15374;
wire _guard15376 = cond_wire690_out;
wire _guard15377 = early_reset_static_par0_go_out;
wire _guard15378 = _guard15376 & _guard15377;
wire _guard15379 = cond_wire722_out;
wire _guard15380 = early_reset_static_par0_go_out;
wire _guard15381 = _guard15379 & _guard15380;
wire _guard15382 = cond_wire722_out;
wire _guard15383 = early_reset_static_par0_go_out;
wire _guard15384 = _guard15382 & _guard15383;
wire _guard15385 = cond_wire804_out;
wire _guard15386 = early_reset_static_par0_go_out;
wire _guard15387 = _guard15385 & _guard15386;
wire _guard15388 = cond_wire804_out;
wire _guard15389 = early_reset_static_par0_go_out;
wire _guard15390 = _guard15388 & _guard15389;
wire _guard15391 = cond_wire783_out;
wire _guard15392 = early_reset_static_par0_go_out;
wire _guard15393 = _guard15391 & _guard15392;
wire _guard15394 = cond_wire783_out;
wire _guard15395 = early_reset_static_par0_go_out;
wire _guard15396 = _guard15394 & _guard15395;
wire _guard15397 = cond_wire866_out;
wire _guard15398 = early_reset_static_par0_go_out;
wire _guard15399 = _guard15397 & _guard15398;
wire _guard15400 = cond_wire864_out;
wire _guard15401 = early_reset_static_par0_go_out;
wire _guard15402 = _guard15400 & _guard15401;
wire _guard15403 = fsm_out == 1'd0;
wire _guard15404 = cond_wire864_out;
wire _guard15405 = _guard15403 & _guard15404;
wire _guard15406 = fsm_out == 1'd0;
wire _guard15407 = _guard15405 & _guard15406;
wire _guard15408 = fsm_out == 1'd0;
wire _guard15409 = cond_wire866_out;
wire _guard15410 = _guard15408 & _guard15409;
wire _guard15411 = fsm_out == 1'd0;
wire _guard15412 = _guard15410 & _guard15411;
wire _guard15413 = _guard15407 | _guard15412;
wire _guard15414 = early_reset_static_par0_go_out;
wire _guard15415 = _guard15413 & _guard15414;
wire _guard15416 = fsm_out == 1'd0;
wire _guard15417 = cond_wire864_out;
wire _guard15418 = _guard15416 & _guard15417;
wire _guard15419 = fsm_out == 1'd0;
wire _guard15420 = _guard15418 & _guard15419;
wire _guard15421 = fsm_out == 1'd0;
wire _guard15422 = cond_wire866_out;
wire _guard15423 = _guard15421 & _guard15422;
wire _guard15424 = fsm_out == 1'd0;
wire _guard15425 = _guard15423 & _guard15424;
wire _guard15426 = _guard15420 | _guard15425;
wire _guard15427 = early_reset_static_par0_go_out;
wire _guard15428 = _guard15426 & _guard15427;
wire _guard15429 = fsm_out == 1'd0;
wire _guard15430 = cond_wire864_out;
wire _guard15431 = _guard15429 & _guard15430;
wire _guard15432 = fsm_out == 1'd0;
wire _guard15433 = _guard15431 & _guard15432;
wire _guard15434 = fsm_out == 1'd0;
wire _guard15435 = cond_wire866_out;
wire _guard15436 = _guard15434 & _guard15435;
wire _guard15437 = fsm_out == 1'd0;
wire _guard15438 = _guard15436 & _guard15437;
wire _guard15439 = _guard15433 | _guard15438;
wire _guard15440 = early_reset_static_par0_go_out;
wire _guard15441 = _guard15439 & _guard15440;
wire _guard15442 = cond_wire800_out;
wire _guard15443 = early_reset_static_par0_go_out;
wire _guard15444 = _guard15442 & _guard15443;
wire _guard15445 = cond_wire800_out;
wire _guard15446 = early_reset_static_par0_go_out;
wire _guard15447 = _guard15445 & _guard15446;
wire _guard15448 = cond_wire927_out;
wire _guard15449 = early_reset_static_par0_go_out;
wire _guard15450 = _guard15448 & _guard15449;
wire _guard15451 = cond_wire925_out;
wire _guard15452 = early_reset_static_par0_go_out;
wire _guard15453 = _guard15451 & _guard15452;
wire _guard15454 = fsm_out == 1'd0;
wire _guard15455 = cond_wire925_out;
wire _guard15456 = _guard15454 & _guard15455;
wire _guard15457 = fsm_out == 1'd0;
wire _guard15458 = _guard15456 & _guard15457;
wire _guard15459 = fsm_out == 1'd0;
wire _guard15460 = cond_wire927_out;
wire _guard15461 = _guard15459 & _guard15460;
wire _guard15462 = fsm_out == 1'd0;
wire _guard15463 = _guard15461 & _guard15462;
wire _guard15464 = _guard15458 | _guard15463;
wire _guard15465 = early_reset_static_par0_go_out;
wire _guard15466 = _guard15464 & _guard15465;
wire _guard15467 = fsm_out == 1'd0;
wire _guard15468 = cond_wire925_out;
wire _guard15469 = _guard15467 & _guard15468;
wire _guard15470 = fsm_out == 1'd0;
wire _guard15471 = _guard15469 & _guard15470;
wire _guard15472 = fsm_out == 1'd0;
wire _guard15473 = cond_wire927_out;
wire _guard15474 = _guard15472 & _guard15473;
wire _guard15475 = fsm_out == 1'd0;
wire _guard15476 = _guard15474 & _guard15475;
wire _guard15477 = _guard15471 | _guard15476;
wire _guard15478 = early_reset_static_par0_go_out;
wire _guard15479 = _guard15477 & _guard15478;
wire _guard15480 = fsm_out == 1'd0;
wire _guard15481 = cond_wire925_out;
wire _guard15482 = _guard15480 & _guard15481;
wire _guard15483 = fsm_out == 1'd0;
wire _guard15484 = _guard15482 & _guard15483;
wire _guard15485 = fsm_out == 1'd0;
wire _guard15486 = cond_wire927_out;
wire _guard15487 = _guard15485 & _guard15486;
wire _guard15488 = fsm_out == 1'd0;
wire _guard15489 = _guard15487 & _guard15488;
wire _guard15490 = _guard15484 | _guard15489;
wire _guard15491 = early_reset_static_par0_go_out;
wire _guard15492 = _guard15490 & _guard15491;
wire _guard15493 = cond_wire947_out;
wire _guard15494 = early_reset_static_par0_go_out;
wire _guard15495 = _guard15493 & _guard15494;
wire _guard15496 = cond_wire945_out;
wire _guard15497 = early_reset_static_par0_go_out;
wire _guard15498 = _guard15496 & _guard15497;
wire _guard15499 = fsm_out == 1'd0;
wire _guard15500 = cond_wire945_out;
wire _guard15501 = _guard15499 & _guard15500;
wire _guard15502 = fsm_out == 1'd0;
wire _guard15503 = _guard15501 & _guard15502;
wire _guard15504 = fsm_out == 1'd0;
wire _guard15505 = cond_wire947_out;
wire _guard15506 = _guard15504 & _guard15505;
wire _guard15507 = fsm_out == 1'd0;
wire _guard15508 = _guard15506 & _guard15507;
wire _guard15509 = _guard15503 | _guard15508;
wire _guard15510 = early_reset_static_par0_go_out;
wire _guard15511 = _guard15509 & _guard15510;
wire _guard15512 = fsm_out == 1'd0;
wire _guard15513 = cond_wire945_out;
wire _guard15514 = _guard15512 & _guard15513;
wire _guard15515 = fsm_out == 1'd0;
wire _guard15516 = _guard15514 & _guard15515;
wire _guard15517 = fsm_out == 1'd0;
wire _guard15518 = cond_wire947_out;
wire _guard15519 = _guard15517 & _guard15518;
wire _guard15520 = fsm_out == 1'd0;
wire _guard15521 = _guard15519 & _guard15520;
wire _guard15522 = _guard15516 | _guard15521;
wire _guard15523 = early_reset_static_par0_go_out;
wire _guard15524 = _guard15522 & _guard15523;
wire _guard15525 = fsm_out == 1'd0;
wire _guard15526 = cond_wire945_out;
wire _guard15527 = _guard15525 & _guard15526;
wire _guard15528 = fsm_out == 1'd0;
wire _guard15529 = _guard15527 & _guard15528;
wire _guard15530 = fsm_out == 1'd0;
wire _guard15531 = cond_wire947_out;
wire _guard15532 = _guard15530 & _guard15531;
wire _guard15533 = fsm_out == 1'd0;
wire _guard15534 = _guard15532 & _guard15533;
wire _guard15535 = _guard15529 | _guard15534;
wire _guard15536 = early_reset_static_par0_go_out;
wire _guard15537 = _guard15535 & _guard15536;
wire _guard15538 = cond_wire881_out;
wire _guard15539 = early_reset_static_par0_go_out;
wire _guard15540 = _guard15538 & _guard15539;
wire _guard15541 = cond_wire881_out;
wire _guard15542 = early_reset_static_par0_go_out;
wire _guard15543 = _guard15541 & _guard15542;
wire _guard15544 = cond_wire1007_out;
wire _guard15545 = early_reset_static_par0_go_out;
wire _guard15546 = _guard15544 & _guard15545;
wire _guard15547 = cond_wire1007_out;
wire _guard15548 = early_reset_static_par0_go_out;
wire _guard15549 = _guard15547 & _guard15548;
wire _guard15550 = cond_wire1040_out;
wire _guard15551 = early_reset_static_par0_go_out;
wire _guard15552 = _guard15550 & _guard15551;
wire _guard15553 = cond_wire1038_out;
wire _guard15554 = early_reset_static_par0_go_out;
wire _guard15555 = _guard15553 & _guard15554;
wire _guard15556 = fsm_out == 1'd0;
wire _guard15557 = cond_wire1038_out;
wire _guard15558 = _guard15556 & _guard15557;
wire _guard15559 = fsm_out == 1'd0;
wire _guard15560 = _guard15558 & _guard15559;
wire _guard15561 = fsm_out == 1'd0;
wire _guard15562 = cond_wire1040_out;
wire _guard15563 = _guard15561 & _guard15562;
wire _guard15564 = fsm_out == 1'd0;
wire _guard15565 = _guard15563 & _guard15564;
wire _guard15566 = _guard15560 | _guard15565;
wire _guard15567 = early_reset_static_par0_go_out;
wire _guard15568 = _guard15566 & _guard15567;
wire _guard15569 = fsm_out == 1'd0;
wire _guard15570 = cond_wire1038_out;
wire _guard15571 = _guard15569 & _guard15570;
wire _guard15572 = fsm_out == 1'd0;
wire _guard15573 = _guard15571 & _guard15572;
wire _guard15574 = fsm_out == 1'd0;
wire _guard15575 = cond_wire1040_out;
wire _guard15576 = _guard15574 & _guard15575;
wire _guard15577 = fsm_out == 1'd0;
wire _guard15578 = _guard15576 & _guard15577;
wire _guard15579 = _guard15573 | _guard15578;
wire _guard15580 = early_reset_static_par0_go_out;
wire _guard15581 = _guard15579 & _guard15580;
wire _guard15582 = fsm_out == 1'd0;
wire _guard15583 = cond_wire1038_out;
wire _guard15584 = _guard15582 & _guard15583;
wire _guard15585 = fsm_out == 1'd0;
wire _guard15586 = _guard15584 & _guard15585;
wire _guard15587 = fsm_out == 1'd0;
wire _guard15588 = cond_wire1040_out;
wire _guard15589 = _guard15587 & _guard15588;
wire _guard15590 = fsm_out == 1'd0;
wire _guard15591 = _guard15589 & _guard15590;
wire _guard15592 = _guard15586 | _guard15591;
wire _guard15593 = early_reset_static_par0_go_out;
wire _guard15594 = _guard15592 & _guard15593;
wire _guard15595 = cond_wire34_out;
wire _guard15596 = early_reset_static_par0_go_out;
wire _guard15597 = _guard15595 & _guard15596;
wire _guard15598 = cond_wire34_out;
wire _guard15599 = early_reset_static_par0_go_out;
wire _guard15600 = _guard15598 & _guard15599;
wire _guard15601 = cond_wire64_out;
wire _guard15602 = early_reset_static_par0_go_out;
wire _guard15603 = _guard15601 & _guard15602;
wire _guard15604 = cond_wire64_out;
wire _guard15605 = early_reset_static_par0_go_out;
wire _guard15606 = _guard15604 & _guard15605;
wire _guard15607 = fsm0_out == 6'd0;
wire _guard15608 = early_reset_static_seq_go_out;
wire _guard15609 = _guard15607 & _guard15608;
wire _guard15610 = cond_wire274_out;
wire _guard15611 = early_reset_static_par0_go_out;
wire _guard15612 = _guard15610 & _guard15611;
wire _guard15613 = _guard15609 | _guard15612;
wire _guard15614 = fsm0_out == 6'd0;
wire _guard15615 = early_reset_static_seq_go_out;
wire _guard15616 = _guard15614 & _guard15615;
wire _guard15617 = cond_wire274_out;
wire _guard15618 = early_reset_static_par0_go_out;
wire _guard15619 = _guard15617 & _guard15618;
wire _guard15620 = cond_wire664_out;
wire _guard15621 = early_reset_static_par0_go_out;
wire _guard15622 = _guard15620 & _guard15621;
wire _guard15623 = cond_wire664_out;
wire _guard15624 = early_reset_static_par0_go_out;
wire _guard15625 = _guard15623 & _guard15624;
wire _guard15626 = fsm0_out == 6'd0;
wire _guard15627 = early_reset_static_seq_go_out;
wire _guard15628 = _guard15626 & _guard15627;
wire _guard15629 = cond_wire989_out;
wire _guard15630 = early_reset_static_par0_go_out;
wire _guard15631 = _guard15629 & _guard15630;
wire _guard15632 = _guard15628 | _guard15631;
wire _guard15633 = cond_wire989_out;
wire _guard15634 = early_reset_static_par0_go_out;
wire _guard15635 = _guard15633 & _guard15634;
wire _guard15636 = fsm0_out == 6'd0;
wire _guard15637 = early_reset_static_seq_go_out;
wire _guard15638 = _guard15636 & _guard15637;
wire _guard15639 = fsm0_out == 6'd0;
wire _guard15640 = early_reset_static_seq_go_out;
wire _guard15641 = _guard15639 & _guard15640;
wire _guard15642 = early_reset_static_par0_go_out;
wire _guard15643 = _guard15641 | _guard15642;
wire _guard15644 = early_reset_static_par0_go_out;
wire _guard15645 = fsm0_out == 6'd0;
wire _guard15646 = early_reset_static_seq_go_out;
wire _guard15647 = _guard15645 & _guard15646;
wire _guard15648 = fsm0_out == 6'd0;
wire _guard15649 = early_reset_static_seq_go_out;
wire _guard15650 = _guard15648 & _guard15649;
wire _guard15651 = early_reset_static_par0_go_out;
wire _guard15652 = _guard15650 | _guard15651;
wire _guard15653 = early_reset_static_par0_go_out;
wire _guard15654 = fsm0_out == 6'd0;
wire _guard15655 = early_reset_static_seq_go_out;
wire _guard15656 = _guard15654 & _guard15655;
wire _guard15657 = fsm0_out == 6'd0;
wire _guard15658 = early_reset_static_seq_go_out;
wire _guard15659 = _guard15657 & _guard15658;
wire _guard15660 = early_reset_static_par0_go_out;
wire _guard15661 = _guard15659 | _guard15660;
wire _guard15662 = early_reset_static_par0_go_out;
wire _guard15663 = fsm0_out == 6'd0;
wire _guard15664 = early_reset_static_seq_go_out;
wire _guard15665 = _guard15663 & _guard15664;
wire _guard15666 = early_reset_static_par0_go_out;
wire _guard15667 = early_reset_static_par0_go_out;
wire _guard15668 = early_reset_static_par0_go_out;
wire _guard15669 = early_reset_static_par0_go_out;
wire _guard15670 = fsm0_out == 6'd0;
wire _guard15671 = early_reset_static_seq_go_out;
wire _guard15672 = _guard15670 & _guard15671;
wire _guard15673 = early_reset_static_par0_go_out;
wire _guard15674 = _guard15672 | _guard15673;
wire _guard15675 = fsm0_out == 6'd0;
wire _guard15676 = early_reset_static_seq_go_out;
wire _guard15677 = _guard15675 & _guard15676;
wire _guard15678 = early_reset_static_par0_go_out;
wire _guard15679 = early_reset_static_par0_go_out;
wire _guard15680 = early_reset_static_par0_go_out;
wire _guard15681 = early_reset_static_par0_go_out;
wire _guard15682 = early_reset_static_par0_go_out;
wire _guard15683 = early_reset_static_par0_go_out;
wire _guard15684 = early_reset_static_par0_go_out;
wire _guard15685 = early_reset_static_par0_go_out;
wire _guard15686 = early_reset_static_par0_go_out;
wire _guard15687 = early_reset_static_par0_go_out;
wire _guard15688 = early_reset_static_par0_go_out;
wire _guard15689 = early_reset_static_par0_go_out;
wire _guard15690 = early_reset_static_par0_go_out;
wire _guard15691 = early_reset_static_par0_go_out;
wire _guard15692 = early_reset_static_par0_go_out;
wire _guard15693 = fsm0_out == 6'd0;
wire _guard15694 = early_reset_static_seq_go_out;
wire _guard15695 = _guard15693 & _guard15694;
wire _guard15696 = early_reset_static_par0_go_out;
wire _guard15697 = _guard15695 | _guard15696;
wire _guard15698 = early_reset_static_par0_go_out;
wire _guard15699 = fsm0_out == 6'd0;
wire _guard15700 = early_reset_static_seq_go_out;
wire _guard15701 = _guard15699 & _guard15700;
wire _guard15702 = early_reset_static_par0_go_out;
wire _guard15703 = early_reset_static_par0_go_out;
wire _guard15704 = early_reset_static_par0_go_out;
wire _guard15705 = early_reset_static_par0_go_out;
wire _guard15706 = early_reset_static_par0_go_out;
wire _guard15707 = early_reset_static_par0_go_out;
wire _guard15708 = early_reset_static_par0_go_out;
wire _guard15709 = early_reset_static_par0_go_out;
wire _guard15710 = early_reset_static_par0_go_out;
wire _guard15711 = early_reset_static_par0_go_out;
wire _guard15712 = early_reset_static_par0_go_out;
wire _guard15713 = early_reset_static_par0_go_out;
wire _guard15714 = early_reset_static_par0_go_out;
wire _guard15715 = ~_guard0;
wire _guard15716 = early_reset_static_par0_go_out;
wire _guard15717 = _guard15715 & _guard15716;
wire _guard15718 = early_reset_static_par0_go_out;
wire _guard15719 = early_reset_static_par0_go_out;
wire _guard15720 = early_reset_static_par0_go_out;
wire _guard15721 = early_reset_static_par0_go_out;
wire _guard15722 = early_reset_static_par0_go_out;
wire _guard15723 = ~_guard0;
wire _guard15724 = early_reset_static_par0_go_out;
wire _guard15725 = _guard15723 & _guard15724;
wire _guard15726 = early_reset_static_par0_go_out;
wire _guard15727 = early_reset_static_par0_go_out;
wire _guard15728 = early_reset_static_par0_go_out;
wire _guard15729 = early_reset_static_par0_go_out;
wire _guard15730 = early_reset_static_par0_go_out;
wire _guard15731 = ~_guard0;
wire _guard15732 = early_reset_static_par0_go_out;
wire _guard15733 = _guard15731 & _guard15732;
wire _guard15734 = early_reset_static_par0_go_out;
wire _guard15735 = early_reset_static_par0_go_out;
wire _guard15736 = ~_guard0;
wire _guard15737 = early_reset_static_par0_go_out;
wire _guard15738 = _guard15736 & _guard15737;
wire _guard15739 = early_reset_static_par0_go_out;
wire _guard15740 = early_reset_static_par0_go_out;
wire _guard15741 = ~_guard0;
wire _guard15742 = early_reset_static_par0_go_out;
wire _guard15743 = _guard15741 & _guard15742;
wire _guard15744 = ~_guard0;
wire _guard15745 = early_reset_static_par0_go_out;
wire _guard15746 = _guard15744 & _guard15745;
wire _guard15747 = early_reset_static_par0_go_out;
wire _guard15748 = early_reset_static_par0_go_out;
wire _guard15749 = ~_guard0;
wire _guard15750 = early_reset_static_par0_go_out;
wire _guard15751 = _guard15749 & _guard15750;
wire _guard15752 = early_reset_static_par0_go_out;
wire _guard15753 = early_reset_static_par0_go_out;
wire _guard15754 = early_reset_static_par0_go_out;
wire _guard15755 = ~_guard0;
wire _guard15756 = early_reset_static_par0_go_out;
wire _guard15757 = _guard15755 & _guard15756;
wire _guard15758 = early_reset_static_par0_go_out;
wire _guard15759 = ~_guard0;
wire _guard15760 = early_reset_static_par0_go_out;
wire _guard15761 = _guard15759 & _guard15760;
wire _guard15762 = early_reset_static_par0_go_out;
wire _guard15763 = early_reset_static_par0_go_out;
wire _guard15764 = ~_guard0;
wire _guard15765 = early_reset_static_par0_go_out;
wire _guard15766 = _guard15764 & _guard15765;
wire _guard15767 = early_reset_static_par0_go_out;
wire _guard15768 = early_reset_static_par0_go_out;
wire _guard15769 = early_reset_static_par0_go_out;
wire _guard15770 = early_reset_static_par0_go_out;
wire _guard15771 = ~_guard0;
wire _guard15772 = early_reset_static_par0_go_out;
wire _guard15773 = _guard15771 & _guard15772;
wire _guard15774 = early_reset_static_par0_go_out;
wire _guard15775 = ~_guard0;
wire _guard15776 = early_reset_static_par0_go_out;
wire _guard15777 = _guard15775 & _guard15776;
wire _guard15778 = early_reset_static_par0_go_out;
wire _guard15779 = ~_guard0;
wire _guard15780 = early_reset_static_par0_go_out;
wire _guard15781 = _guard15779 & _guard15780;
wire _guard15782 = early_reset_static_par0_go_out;
wire _guard15783 = ~_guard0;
wire _guard15784 = early_reset_static_par0_go_out;
wire _guard15785 = _guard15783 & _guard15784;
wire _guard15786 = early_reset_static_par0_go_out;
wire _guard15787 = early_reset_static_par0_go_out;
wire _guard15788 = early_reset_static_par0_go_out;
wire _guard15789 = early_reset_static_par0_go_out;
wire _guard15790 = early_reset_static_par0_go_out;
wire _guard15791 = early_reset_static_par0_go_out;
wire _guard15792 = early_reset_static_par0_go_out;
wire _guard15793 = ~_guard0;
wire _guard15794 = early_reset_static_par0_go_out;
wire _guard15795 = _guard15793 & _guard15794;
wire _guard15796 = early_reset_static_par0_go_out;
wire _guard15797 = ~_guard0;
wire _guard15798 = early_reset_static_par0_go_out;
wire _guard15799 = _guard15797 & _guard15798;
wire _guard15800 = early_reset_static_par0_go_out;
wire _guard15801 = early_reset_static_par0_go_out;
wire _guard15802 = early_reset_static_par0_go_out;
wire _guard15803 = early_reset_static_par0_go_out;
wire _guard15804 = early_reset_static_par0_go_out;
wire _guard15805 = early_reset_static_par0_go_out;
wire _guard15806 = ~_guard0;
wire _guard15807 = early_reset_static_par0_go_out;
wire _guard15808 = _guard15806 & _guard15807;
wire _guard15809 = early_reset_static_par0_go_out;
wire _guard15810 = early_reset_static_par0_go_out;
wire _guard15811 = ~_guard0;
wire _guard15812 = early_reset_static_par0_go_out;
wire _guard15813 = _guard15811 & _guard15812;
wire _guard15814 = early_reset_static_par0_go_out;
wire _guard15815 = early_reset_static_par0_go_out;
wire _guard15816 = early_reset_static_par0_go_out;
wire _guard15817 = early_reset_static_par0_go_out;
wire _guard15818 = early_reset_static_par0_go_out;
wire _guard15819 = early_reset_static_par0_go_out;
wire _guard15820 = early_reset_static_par0_go_out;
wire _guard15821 = early_reset_static_par0_go_out;
wire _guard15822 = early_reset_static_par0_go_out;
wire _guard15823 = early_reset_static_par0_go_out;
wire _guard15824 = early_reset_static_par0_go_out;
wire _guard15825 = early_reset_static_par0_go_out;
wire _guard15826 = ~_guard0;
wire _guard15827 = early_reset_static_par0_go_out;
wire _guard15828 = _guard15826 & _guard15827;
wire _guard15829 = early_reset_static_par0_go_out;
wire _guard15830 = early_reset_static_par0_go_out;
wire _guard15831 = ~_guard0;
wire _guard15832 = early_reset_static_par0_go_out;
wire _guard15833 = _guard15831 & _guard15832;
wire _guard15834 = early_reset_static_par0_go_out;
wire _guard15835 = ~_guard0;
wire _guard15836 = early_reset_static_par0_go_out;
wire _guard15837 = _guard15835 & _guard15836;
wire _guard15838 = early_reset_static_par0_go_out;
wire _guard15839 = early_reset_static_par0_go_out;
wire _guard15840 = early_reset_static_par0_go_out;
wire _guard15841 = early_reset_static_par0_go_out;
wire _guard15842 = early_reset_static_par0_go_out;
wire _guard15843 = early_reset_static_par0_go_out;
wire _guard15844 = early_reset_static_par0_go_out;
wire _guard15845 = ~_guard0;
wire _guard15846 = early_reset_static_par0_go_out;
wire _guard15847 = _guard15845 & _guard15846;
wire _guard15848 = early_reset_static_par0_go_out;
wire _guard15849 = early_reset_static_par0_go_out;
wire _guard15850 = early_reset_static_par0_go_out;
wire _guard15851 = early_reset_static_par0_go_out;
wire _guard15852 = early_reset_static_par0_go_out;
wire _guard15853 = ~_guard0;
wire _guard15854 = early_reset_static_par0_go_out;
wire _guard15855 = _guard15853 & _guard15854;
wire _guard15856 = ~_guard0;
wire _guard15857 = early_reset_static_par0_go_out;
wire _guard15858 = _guard15856 & _guard15857;
wire _guard15859 = early_reset_static_par0_go_out;
wire _guard15860 = early_reset_static_par0_go_out;
wire _guard15861 = early_reset_static_par0_go_out;
wire _guard15862 = early_reset_static_par0_go_out;
wire _guard15863 = ~_guard0;
wire _guard15864 = early_reset_static_par0_go_out;
wire _guard15865 = _guard15863 & _guard15864;
wire _guard15866 = early_reset_static_par0_go_out;
wire _guard15867 = ~_guard0;
wire _guard15868 = early_reset_static_par0_go_out;
wire _guard15869 = _guard15867 & _guard15868;
wire _guard15870 = early_reset_static_par0_go_out;
wire _guard15871 = early_reset_static_par0_go_out;
wire _guard15872 = early_reset_static_par0_go_out;
wire _guard15873 = early_reset_static_par0_go_out;
wire _guard15874 = ~_guard0;
wire _guard15875 = early_reset_static_par0_go_out;
wire _guard15876 = _guard15874 & _guard15875;
wire _guard15877 = early_reset_static_par0_go_out;
wire _guard15878 = early_reset_static_par0_go_out;
wire _guard15879 = ~_guard0;
wire _guard15880 = early_reset_static_par0_go_out;
wire _guard15881 = _guard15879 & _guard15880;
wire _guard15882 = early_reset_static_par0_go_out;
wire _guard15883 = early_reset_static_par0_go_out;
wire _guard15884 = early_reset_static_par0_go_out;
wire _guard15885 = ~_guard0;
wire _guard15886 = early_reset_static_par0_go_out;
wire _guard15887 = _guard15885 & _guard15886;
wire _guard15888 = ~_guard0;
wire _guard15889 = early_reset_static_par0_go_out;
wire _guard15890 = _guard15888 & _guard15889;
wire _guard15891 = early_reset_static_par0_go_out;
wire _guard15892 = early_reset_static_par0_go_out;
wire _guard15893 = early_reset_static_par0_go_out;
wire _guard15894 = early_reset_static_par0_go_out;
wire _guard15895 = early_reset_static_par0_go_out;
wire _guard15896 = early_reset_static_par0_go_out;
wire _guard15897 = early_reset_static_par0_go_out;
wire _guard15898 = early_reset_static_par0_go_out;
wire _guard15899 = ~_guard0;
wire _guard15900 = early_reset_static_par0_go_out;
wire _guard15901 = _guard15899 & _guard15900;
wire _guard15902 = ~_guard0;
wire _guard15903 = early_reset_static_par0_go_out;
wire _guard15904 = _guard15902 & _guard15903;
wire _guard15905 = early_reset_static_par0_go_out;
wire _guard15906 = early_reset_static_par0_go_out;
wire _guard15907 = early_reset_static_par0_go_out;
wire _guard15908 = ~_guard0;
wire _guard15909 = early_reset_static_par0_go_out;
wire _guard15910 = _guard15908 & _guard15909;
wire _guard15911 = early_reset_static_par0_go_out;
wire _guard15912 = early_reset_static_par0_go_out;
wire _guard15913 = early_reset_static_par0_go_out;
wire _guard15914 = early_reset_static_par0_go_out;
wire _guard15915 = early_reset_static_par0_go_out;
wire _guard15916 = early_reset_static_par0_go_out;
wire _guard15917 = early_reset_static_par0_go_out;
wire _guard15918 = early_reset_static_par0_go_out;
wire _guard15919 = early_reset_static_par0_go_out;
wire _guard15920 = early_reset_static_par0_go_out;
wire _guard15921 = ~_guard0;
wire _guard15922 = early_reset_static_par0_go_out;
wire _guard15923 = _guard15921 & _guard15922;
wire _guard15924 = early_reset_static_par0_go_out;
wire _guard15925 = early_reset_static_par0_go_out;
wire _guard15926 = early_reset_static_par0_go_out;
wire _guard15927 = early_reset_static_par0_go_out;
wire _guard15928 = early_reset_static_par0_go_out;
wire _guard15929 = ~_guard0;
wire _guard15930 = early_reset_static_par0_go_out;
wire _guard15931 = _guard15929 & _guard15930;
wire _guard15932 = early_reset_static_par0_go_out;
wire _guard15933 = ~_guard0;
wire _guard15934 = early_reset_static_par0_go_out;
wire _guard15935 = _guard15933 & _guard15934;
wire _guard15936 = early_reset_static_par0_go_out;
wire _guard15937 = early_reset_static_par0_go_out;
wire _guard15938 = ~_guard0;
wire _guard15939 = early_reset_static_par0_go_out;
wire _guard15940 = _guard15938 & _guard15939;
wire _guard15941 = early_reset_static_par0_go_out;
wire _guard15942 = early_reset_static_par0_go_out;
wire _guard15943 = early_reset_static_par0_go_out;
wire _guard15944 = early_reset_static_par0_go_out;
wire _guard15945 = early_reset_static_par0_go_out;
wire _guard15946 = early_reset_static_par0_go_out;
wire _guard15947 = early_reset_static_par0_go_out;
wire _guard15948 = early_reset_static_par0_go_out;
wire _guard15949 = ~_guard0;
wire _guard15950 = early_reset_static_par0_go_out;
wire _guard15951 = _guard15949 & _guard15950;
wire _guard15952 = ~_guard0;
wire _guard15953 = early_reset_static_par0_go_out;
wire _guard15954 = _guard15952 & _guard15953;
wire _guard15955 = early_reset_static_par0_go_out;
wire _guard15956 = early_reset_static_par0_go_out;
wire _guard15957 = early_reset_static_par0_go_out;
wire _guard15958 = ~_guard0;
wire _guard15959 = early_reset_static_par0_go_out;
wire _guard15960 = _guard15958 & _guard15959;
wire _guard15961 = early_reset_static_par0_go_out;
wire _guard15962 = ~_guard0;
wire _guard15963 = early_reset_static_par0_go_out;
wire _guard15964 = _guard15962 & _guard15963;
wire _guard15965 = early_reset_static_par0_go_out;
wire _guard15966 = ~_guard0;
wire _guard15967 = early_reset_static_par0_go_out;
wire _guard15968 = _guard15966 & _guard15967;
wire _guard15969 = early_reset_static_par0_go_out;
wire _guard15970 = early_reset_static_par0_go_out;
wire _guard15971 = ~_guard0;
wire _guard15972 = early_reset_static_par0_go_out;
wire _guard15973 = _guard15971 & _guard15972;
wire _guard15974 = ~_guard0;
wire _guard15975 = early_reset_static_par0_go_out;
wire _guard15976 = _guard15974 & _guard15975;
wire _guard15977 = early_reset_static_par0_go_out;
wire _guard15978 = ~_guard0;
wire _guard15979 = early_reset_static_par0_go_out;
wire _guard15980 = _guard15978 & _guard15979;
wire _guard15981 = early_reset_static_par0_go_out;
wire _guard15982 = early_reset_static_par0_go_out;
wire _guard15983 = early_reset_static_par0_go_out;
wire _guard15984 = early_reset_static_par0_go_out;
wire _guard15985 = early_reset_static_par0_go_out;
wire _guard15986 = early_reset_static_par0_go_out;
wire _guard15987 = early_reset_static_par0_go_out;
wire _guard15988 = ~_guard0;
wire _guard15989 = early_reset_static_par0_go_out;
wire _guard15990 = _guard15988 & _guard15989;
wire _guard15991 = early_reset_static_par0_go_out;
wire _guard15992 = early_reset_static_par0_go_out;
wire _guard15993 = early_reset_static_par0_go_out;
wire _guard15994 = early_reset_static_par0_go_out;
wire _guard15995 = early_reset_static_par0_go_out;
wire _guard15996 = early_reset_static_par0_go_out;
wire _guard15997 = early_reset_static_par0_go_out;
wire _guard15998 = ~_guard0;
wire _guard15999 = early_reset_static_par0_go_out;
wire _guard16000 = _guard15998 & _guard15999;
wire _guard16001 = early_reset_static_par0_go_out;
wire _guard16002 = early_reset_static_par0_go_out;
wire _guard16003 = ~_guard0;
wire _guard16004 = early_reset_static_par0_go_out;
wire _guard16005 = _guard16003 & _guard16004;
wire _guard16006 = early_reset_static_par0_go_out;
wire _guard16007 = early_reset_static_par0_go_out;
wire _guard16008 = ~_guard0;
wire _guard16009 = early_reset_static_par0_go_out;
wire _guard16010 = _guard16008 & _guard16009;
wire _guard16011 = early_reset_static_par0_go_out;
wire _guard16012 = early_reset_static_par0_go_out;
wire _guard16013 = early_reset_static_par0_go_out;
wire _guard16014 = ~_guard0;
wire _guard16015 = early_reset_static_par0_go_out;
wire _guard16016 = _guard16014 & _guard16015;
wire _guard16017 = early_reset_static_par0_go_out;
wire _guard16018 = early_reset_static_par0_go_out;
wire _guard16019 = ~_guard0;
wire _guard16020 = early_reset_static_par0_go_out;
wire _guard16021 = _guard16019 & _guard16020;
wire _guard16022 = ~_guard0;
wire _guard16023 = early_reset_static_par0_go_out;
wire _guard16024 = _guard16022 & _guard16023;
wire _guard16025 = early_reset_static_par0_go_out;
wire _guard16026 = ~_guard0;
wire _guard16027 = early_reset_static_par0_go_out;
wire _guard16028 = _guard16026 & _guard16027;
wire _guard16029 = early_reset_static_par0_go_out;
wire _guard16030 = fsm0_out == 6'd0;
wire _guard16031 = signal_reg_out;
wire _guard16032 = _guard16030 & _guard16031;
wire _guard16033 = cond_wire4_out;
wire _guard16034 = early_reset_static_par0_go_out;
wire _guard16035 = _guard16033 & _guard16034;
wire _guard16036 = cond_wire4_out;
wire _guard16037 = early_reset_static_par0_go_out;
wire _guard16038 = _guard16036 & _guard16037;
wire _guard16039 = cond_wire6_out;
wire _guard16040 = early_reset_static_par0_go_out;
wire _guard16041 = _guard16039 & _guard16040;
wire _guard16042 = cond_wire6_out;
wire _guard16043 = early_reset_static_par0_go_out;
wire _guard16044 = _guard16042 & _guard16043;
wire _guard16045 = cond_wire22_out;
wire _guard16046 = early_reset_static_par0_go_out;
wire _guard16047 = _guard16045 & _guard16046;
wire _guard16048 = cond_wire20_out;
wire _guard16049 = early_reset_static_par0_go_out;
wire _guard16050 = _guard16048 & _guard16049;
wire _guard16051 = fsm_out == 1'd0;
wire _guard16052 = cond_wire20_out;
wire _guard16053 = _guard16051 & _guard16052;
wire _guard16054 = fsm_out == 1'd0;
wire _guard16055 = _guard16053 & _guard16054;
wire _guard16056 = fsm_out == 1'd0;
wire _guard16057 = cond_wire22_out;
wire _guard16058 = _guard16056 & _guard16057;
wire _guard16059 = fsm_out == 1'd0;
wire _guard16060 = _guard16058 & _guard16059;
wire _guard16061 = _guard16055 | _guard16060;
wire _guard16062 = early_reset_static_par0_go_out;
wire _guard16063 = _guard16061 & _guard16062;
wire _guard16064 = fsm_out == 1'd0;
wire _guard16065 = cond_wire20_out;
wire _guard16066 = _guard16064 & _guard16065;
wire _guard16067 = fsm_out == 1'd0;
wire _guard16068 = _guard16066 & _guard16067;
wire _guard16069 = fsm_out == 1'd0;
wire _guard16070 = cond_wire22_out;
wire _guard16071 = _guard16069 & _guard16070;
wire _guard16072 = fsm_out == 1'd0;
wire _guard16073 = _guard16071 & _guard16072;
wire _guard16074 = _guard16068 | _guard16073;
wire _guard16075 = early_reset_static_par0_go_out;
wire _guard16076 = _guard16074 & _guard16075;
wire _guard16077 = fsm_out == 1'd0;
wire _guard16078 = cond_wire20_out;
wire _guard16079 = _guard16077 & _guard16078;
wire _guard16080 = fsm_out == 1'd0;
wire _guard16081 = _guard16079 & _guard16080;
wire _guard16082 = fsm_out == 1'd0;
wire _guard16083 = cond_wire22_out;
wire _guard16084 = _guard16082 & _guard16083;
wire _guard16085 = fsm_out == 1'd0;
wire _guard16086 = _guard16084 & _guard16085;
wire _guard16087 = _guard16081 | _guard16086;
wire _guard16088 = early_reset_static_par0_go_out;
wire _guard16089 = _guard16087 & _guard16088;
wire _guard16090 = cond_wire44_out;
wire _guard16091 = early_reset_static_par0_go_out;
wire _guard16092 = _guard16090 & _guard16091;
wire _guard16093 = cond_wire44_out;
wire _guard16094 = early_reset_static_par0_go_out;
wire _guard16095 = _guard16093 & _guard16094;
wire _guard16096 = cond_wire46_out;
wire _guard16097 = early_reset_static_par0_go_out;
wire _guard16098 = _guard16096 & _guard16097;
wire _guard16099 = cond_wire46_out;
wire _guard16100 = early_reset_static_par0_go_out;
wire _guard16101 = _guard16099 & _guard16100;
wire _guard16102 = cond_wire72_out;
wire _guard16103 = early_reset_static_par0_go_out;
wire _guard16104 = _guard16102 & _guard16103;
wire _guard16105 = cond_wire70_out;
wire _guard16106 = early_reset_static_par0_go_out;
wire _guard16107 = _guard16105 & _guard16106;
wire _guard16108 = fsm_out == 1'd0;
wire _guard16109 = cond_wire70_out;
wire _guard16110 = _guard16108 & _guard16109;
wire _guard16111 = fsm_out == 1'd0;
wire _guard16112 = _guard16110 & _guard16111;
wire _guard16113 = fsm_out == 1'd0;
wire _guard16114 = cond_wire72_out;
wire _guard16115 = _guard16113 & _guard16114;
wire _guard16116 = fsm_out == 1'd0;
wire _guard16117 = _guard16115 & _guard16116;
wire _guard16118 = _guard16112 | _guard16117;
wire _guard16119 = early_reset_static_par0_go_out;
wire _guard16120 = _guard16118 & _guard16119;
wire _guard16121 = fsm_out == 1'd0;
wire _guard16122 = cond_wire70_out;
wire _guard16123 = _guard16121 & _guard16122;
wire _guard16124 = fsm_out == 1'd0;
wire _guard16125 = _guard16123 & _guard16124;
wire _guard16126 = fsm_out == 1'd0;
wire _guard16127 = cond_wire72_out;
wire _guard16128 = _guard16126 & _guard16127;
wire _guard16129 = fsm_out == 1'd0;
wire _guard16130 = _guard16128 & _guard16129;
wire _guard16131 = _guard16125 | _guard16130;
wire _guard16132 = early_reset_static_par0_go_out;
wire _guard16133 = _guard16131 & _guard16132;
wire _guard16134 = fsm_out == 1'd0;
wire _guard16135 = cond_wire70_out;
wire _guard16136 = _guard16134 & _guard16135;
wire _guard16137 = fsm_out == 1'd0;
wire _guard16138 = _guard16136 & _guard16137;
wire _guard16139 = fsm_out == 1'd0;
wire _guard16140 = cond_wire72_out;
wire _guard16141 = _guard16139 & _guard16140;
wire _guard16142 = fsm_out == 1'd0;
wire _guard16143 = _guard16141 & _guard16142;
wire _guard16144 = _guard16138 | _guard16143;
wire _guard16145 = early_reset_static_par0_go_out;
wire _guard16146 = _guard16144 & _guard16145;
wire _guard16147 = cond_wire118_out;
wire _guard16148 = early_reset_static_par0_go_out;
wire _guard16149 = _guard16147 & _guard16148;
wire _guard16150 = cond_wire116_out;
wire _guard16151 = early_reset_static_par0_go_out;
wire _guard16152 = _guard16150 & _guard16151;
wire _guard16153 = fsm_out == 1'd0;
wire _guard16154 = cond_wire116_out;
wire _guard16155 = _guard16153 & _guard16154;
wire _guard16156 = fsm_out == 1'd0;
wire _guard16157 = _guard16155 & _guard16156;
wire _guard16158 = fsm_out == 1'd0;
wire _guard16159 = cond_wire118_out;
wire _guard16160 = _guard16158 & _guard16159;
wire _guard16161 = fsm_out == 1'd0;
wire _guard16162 = _guard16160 & _guard16161;
wire _guard16163 = _guard16157 | _guard16162;
wire _guard16164 = early_reset_static_par0_go_out;
wire _guard16165 = _guard16163 & _guard16164;
wire _guard16166 = fsm_out == 1'd0;
wire _guard16167 = cond_wire116_out;
wire _guard16168 = _guard16166 & _guard16167;
wire _guard16169 = fsm_out == 1'd0;
wire _guard16170 = _guard16168 & _guard16169;
wire _guard16171 = fsm_out == 1'd0;
wire _guard16172 = cond_wire118_out;
wire _guard16173 = _guard16171 & _guard16172;
wire _guard16174 = fsm_out == 1'd0;
wire _guard16175 = _guard16173 & _guard16174;
wire _guard16176 = _guard16170 | _guard16175;
wire _guard16177 = early_reset_static_par0_go_out;
wire _guard16178 = _guard16176 & _guard16177;
wire _guard16179 = fsm_out == 1'd0;
wire _guard16180 = cond_wire116_out;
wire _guard16181 = _guard16179 & _guard16180;
wire _guard16182 = fsm_out == 1'd0;
wire _guard16183 = _guard16181 & _guard16182;
wire _guard16184 = fsm_out == 1'd0;
wire _guard16185 = cond_wire118_out;
wire _guard16186 = _guard16184 & _guard16185;
wire _guard16187 = fsm_out == 1'd0;
wire _guard16188 = _guard16186 & _guard16187;
wire _guard16189 = _guard16183 | _guard16188;
wire _guard16190 = early_reset_static_par0_go_out;
wire _guard16191 = _guard16189 & _guard16190;
wire _guard16192 = cond_wire93_out;
wire _guard16193 = early_reset_static_par0_go_out;
wire _guard16194 = _guard16192 & _guard16193;
wire _guard16195 = cond_wire93_out;
wire _guard16196 = early_reset_static_par0_go_out;
wire _guard16197 = _guard16195 & _guard16196;
wire _guard16198 = cond_wire171_out;
wire _guard16199 = early_reset_static_par0_go_out;
wire _guard16200 = _guard16198 & _guard16199;
wire _guard16201 = cond_wire169_out;
wire _guard16202 = early_reset_static_par0_go_out;
wire _guard16203 = _guard16201 & _guard16202;
wire _guard16204 = fsm_out == 1'd0;
wire _guard16205 = cond_wire169_out;
wire _guard16206 = _guard16204 & _guard16205;
wire _guard16207 = fsm_out == 1'd0;
wire _guard16208 = _guard16206 & _guard16207;
wire _guard16209 = fsm_out == 1'd0;
wire _guard16210 = cond_wire171_out;
wire _guard16211 = _guard16209 & _guard16210;
wire _guard16212 = fsm_out == 1'd0;
wire _guard16213 = _guard16211 & _guard16212;
wire _guard16214 = _guard16208 | _guard16213;
wire _guard16215 = early_reset_static_par0_go_out;
wire _guard16216 = _guard16214 & _guard16215;
wire _guard16217 = fsm_out == 1'd0;
wire _guard16218 = cond_wire169_out;
wire _guard16219 = _guard16217 & _guard16218;
wire _guard16220 = fsm_out == 1'd0;
wire _guard16221 = _guard16219 & _guard16220;
wire _guard16222 = fsm_out == 1'd0;
wire _guard16223 = cond_wire171_out;
wire _guard16224 = _guard16222 & _guard16223;
wire _guard16225 = fsm_out == 1'd0;
wire _guard16226 = _guard16224 & _guard16225;
wire _guard16227 = _guard16221 | _guard16226;
wire _guard16228 = early_reset_static_par0_go_out;
wire _guard16229 = _guard16227 & _guard16228;
wire _guard16230 = fsm_out == 1'd0;
wire _guard16231 = cond_wire169_out;
wire _guard16232 = _guard16230 & _guard16231;
wire _guard16233 = fsm_out == 1'd0;
wire _guard16234 = _guard16232 & _guard16233;
wire _guard16235 = fsm_out == 1'd0;
wire _guard16236 = cond_wire171_out;
wire _guard16237 = _guard16235 & _guard16236;
wire _guard16238 = fsm_out == 1'd0;
wire _guard16239 = _guard16237 & _guard16238;
wire _guard16240 = _guard16234 | _guard16239;
wire _guard16241 = early_reset_static_par0_go_out;
wire _guard16242 = _guard16240 & _guard16241;
wire _guard16243 = cond_wire179_out;
wire _guard16244 = early_reset_static_par0_go_out;
wire _guard16245 = _guard16243 & _guard16244;
wire _guard16246 = cond_wire177_out;
wire _guard16247 = early_reset_static_par0_go_out;
wire _guard16248 = _guard16246 & _guard16247;
wire _guard16249 = fsm_out == 1'd0;
wire _guard16250 = cond_wire177_out;
wire _guard16251 = _guard16249 & _guard16250;
wire _guard16252 = fsm_out == 1'd0;
wire _guard16253 = _guard16251 & _guard16252;
wire _guard16254 = fsm_out == 1'd0;
wire _guard16255 = cond_wire179_out;
wire _guard16256 = _guard16254 & _guard16255;
wire _guard16257 = fsm_out == 1'd0;
wire _guard16258 = _guard16256 & _guard16257;
wire _guard16259 = _guard16253 | _guard16258;
wire _guard16260 = early_reset_static_par0_go_out;
wire _guard16261 = _guard16259 & _guard16260;
wire _guard16262 = fsm_out == 1'd0;
wire _guard16263 = cond_wire177_out;
wire _guard16264 = _guard16262 & _guard16263;
wire _guard16265 = fsm_out == 1'd0;
wire _guard16266 = _guard16264 & _guard16265;
wire _guard16267 = fsm_out == 1'd0;
wire _guard16268 = cond_wire179_out;
wire _guard16269 = _guard16267 & _guard16268;
wire _guard16270 = fsm_out == 1'd0;
wire _guard16271 = _guard16269 & _guard16270;
wire _guard16272 = _guard16266 | _guard16271;
wire _guard16273 = early_reset_static_par0_go_out;
wire _guard16274 = _guard16272 & _guard16273;
wire _guard16275 = fsm_out == 1'd0;
wire _guard16276 = cond_wire177_out;
wire _guard16277 = _guard16275 & _guard16276;
wire _guard16278 = fsm_out == 1'd0;
wire _guard16279 = _guard16277 & _guard16278;
wire _guard16280 = fsm_out == 1'd0;
wire _guard16281 = cond_wire179_out;
wire _guard16282 = _guard16280 & _guard16281;
wire _guard16283 = fsm_out == 1'd0;
wire _guard16284 = _guard16282 & _guard16283;
wire _guard16285 = _guard16279 | _guard16284;
wire _guard16286 = early_reset_static_par0_go_out;
wire _guard16287 = _guard16285 & _guard16286;
wire _guard16288 = cond_wire133_out;
wire _guard16289 = early_reset_static_par0_go_out;
wire _guard16290 = _guard16288 & _guard16289;
wire _guard16291 = cond_wire133_out;
wire _guard16292 = early_reset_static_par0_go_out;
wire _guard16293 = _guard16291 & _guard16292;
wire _guard16294 = cond_wire209_out;
wire _guard16295 = early_reset_static_par0_go_out;
wire _guard16296 = _guard16294 & _guard16295;
wire _guard16297 = cond_wire209_out;
wire _guard16298 = early_reset_static_par0_go_out;
wire _guard16299 = _guard16297 & _guard16298;
wire _guard16300 = cond_wire248_out;
wire _guard16301 = early_reset_static_par0_go_out;
wire _guard16302 = _guard16300 & _guard16301;
wire _guard16303 = cond_wire246_out;
wire _guard16304 = early_reset_static_par0_go_out;
wire _guard16305 = _guard16303 & _guard16304;
wire _guard16306 = fsm_out == 1'd0;
wire _guard16307 = cond_wire246_out;
wire _guard16308 = _guard16306 & _guard16307;
wire _guard16309 = fsm_out == 1'd0;
wire _guard16310 = _guard16308 & _guard16309;
wire _guard16311 = fsm_out == 1'd0;
wire _guard16312 = cond_wire248_out;
wire _guard16313 = _guard16311 & _guard16312;
wire _guard16314 = fsm_out == 1'd0;
wire _guard16315 = _guard16313 & _guard16314;
wire _guard16316 = _guard16310 | _guard16315;
wire _guard16317 = early_reset_static_par0_go_out;
wire _guard16318 = _guard16316 & _guard16317;
wire _guard16319 = fsm_out == 1'd0;
wire _guard16320 = cond_wire246_out;
wire _guard16321 = _guard16319 & _guard16320;
wire _guard16322 = fsm_out == 1'd0;
wire _guard16323 = _guard16321 & _guard16322;
wire _guard16324 = fsm_out == 1'd0;
wire _guard16325 = cond_wire248_out;
wire _guard16326 = _guard16324 & _guard16325;
wire _guard16327 = fsm_out == 1'd0;
wire _guard16328 = _guard16326 & _guard16327;
wire _guard16329 = _guard16323 | _guard16328;
wire _guard16330 = early_reset_static_par0_go_out;
wire _guard16331 = _guard16329 & _guard16330;
wire _guard16332 = fsm_out == 1'd0;
wire _guard16333 = cond_wire246_out;
wire _guard16334 = _guard16332 & _guard16333;
wire _guard16335 = fsm_out == 1'd0;
wire _guard16336 = _guard16334 & _guard16335;
wire _guard16337 = fsm_out == 1'd0;
wire _guard16338 = cond_wire248_out;
wire _guard16339 = _guard16337 & _guard16338;
wire _guard16340 = fsm_out == 1'd0;
wire _guard16341 = _guard16339 & _guard16340;
wire _guard16342 = _guard16336 | _guard16341;
wire _guard16343 = early_reset_static_par0_go_out;
wire _guard16344 = _guard16342 & _guard16343;
wire _guard16345 = cond_wire256_out;
wire _guard16346 = early_reset_static_par0_go_out;
wire _guard16347 = _guard16345 & _guard16346;
wire _guard16348 = cond_wire254_out;
wire _guard16349 = early_reset_static_par0_go_out;
wire _guard16350 = _guard16348 & _guard16349;
wire _guard16351 = fsm_out == 1'd0;
wire _guard16352 = cond_wire254_out;
wire _guard16353 = _guard16351 & _guard16352;
wire _guard16354 = fsm_out == 1'd0;
wire _guard16355 = _guard16353 & _guard16354;
wire _guard16356 = fsm_out == 1'd0;
wire _guard16357 = cond_wire256_out;
wire _guard16358 = _guard16356 & _guard16357;
wire _guard16359 = fsm_out == 1'd0;
wire _guard16360 = _guard16358 & _guard16359;
wire _guard16361 = _guard16355 | _guard16360;
wire _guard16362 = early_reset_static_par0_go_out;
wire _guard16363 = _guard16361 & _guard16362;
wire _guard16364 = fsm_out == 1'd0;
wire _guard16365 = cond_wire254_out;
wire _guard16366 = _guard16364 & _guard16365;
wire _guard16367 = fsm_out == 1'd0;
wire _guard16368 = _guard16366 & _guard16367;
wire _guard16369 = fsm_out == 1'd0;
wire _guard16370 = cond_wire256_out;
wire _guard16371 = _guard16369 & _guard16370;
wire _guard16372 = fsm_out == 1'd0;
wire _guard16373 = _guard16371 & _guard16372;
wire _guard16374 = _guard16368 | _guard16373;
wire _guard16375 = early_reset_static_par0_go_out;
wire _guard16376 = _guard16374 & _guard16375;
wire _guard16377 = fsm_out == 1'd0;
wire _guard16378 = cond_wire254_out;
wire _guard16379 = _guard16377 & _guard16378;
wire _guard16380 = fsm_out == 1'd0;
wire _guard16381 = _guard16379 & _guard16380;
wire _guard16382 = fsm_out == 1'd0;
wire _guard16383 = cond_wire256_out;
wire _guard16384 = _guard16382 & _guard16383;
wire _guard16385 = fsm_out == 1'd0;
wire _guard16386 = _guard16384 & _guard16385;
wire _guard16387 = _guard16381 | _guard16386;
wire _guard16388 = early_reset_static_par0_go_out;
wire _guard16389 = _guard16387 & _guard16388;
wire _guard16390 = cond_wire285_out;
wire _guard16391 = early_reset_static_par0_go_out;
wire _guard16392 = _guard16390 & _guard16391;
wire _guard16393 = cond_wire283_out;
wire _guard16394 = early_reset_static_par0_go_out;
wire _guard16395 = _guard16393 & _guard16394;
wire _guard16396 = fsm_out == 1'd0;
wire _guard16397 = cond_wire283_out;
wire _guard16398 = _guard16396 & _guard16397;
wire _guard16399 = fsm_out == 1'd0;
wire _guard16400 = _guard16398 & _guard16399;
wire _guard16401 = fsm_out == 1'd0;
wire _guard16402 = cond_wire285_out;
wire _guard16403 = _guard16401 & _guard16402;
wire _guard16404 = fsm_out == 1'd0;
wire _guard16405 = _guard16403 & _guard16404;
wire _guard16406 = _guard16400 | _guard16405;
wire _guard16407 = early_reset_static_par0_go_out;
wire _guard16408 = _guard16406 & _guard16407;
wire _guard16409 = fsm_out == 1'd0;
wire _guard16410 = cond_wire283_out;
wire _guard16411 = _guard16409 & _guard16410;
wire _guard16412 = fsm_out == 1'd0;
wire _guard16413 = _guard16411 & _guard16412;
wire _guard16414 = fsm_out == 1'd0;
wire _guard16415 = cond_wire285_out;
wire _guard16416 = _guard16414 & _guard16415;
wire _guard16417 = fsm_out == 1'd0;
wire _guard16418 = _guard16416 & _guard16417;
wire _guard16419 = _guard16413 | _guard16418;
wire _guard16420 = early_reset_static_par0_go_out;
wire _guard16421 = _guard16419 & _guard16420;
wire _guard16422 = fsm_out == 1'd0;
wire _guard16423 = cond_wire283_out;
wire _guard16424 = _guard16422 & _guard16423;
wire _guard16425 = fsm_out == 1'd0;
wire _guard16426 = _guard16424 & _guard16425;
wire _guard16427 = fsm_out == 1'd0;
wire _guard16428 = cond_wire285_out;
wire _guard16429 = _guard16427 & _guard16428;
wire _guard16430 = fsm_out == 1'd0;
wire _guard16431 = _guard16429 & _guard16430;
wire _guard16432 = _guard16426 | _guard16431;
wire _guard16433 = early_reset_static_par0_go_out;
wire _guard16434 = _guard16432 & _guard16433;
wire _guard16435 = cond_wire309_out;
wire _guard16436 = early_reset_static_par0_go_out;
wire _guard16437 = _guard16435 & _guard16436;
wire _guard16438 = cond_wire307_out;
wire _guard16439 = early_reset_static_par0_go_out;
wire _guard16440 = _guard16438 & _guard16439;
wire _guard16441 = fsm_out == 1'd0;
wire _guard16442 = cond_wire307_out;
wire _guard16443 = _guard16441 & _guard16442;
wire _guard16444 = fsm_out == 1'd0;
wire _guard16445 = _guard16443 & _guard16444;
wire _guard16446 = fsm_out == 1'd0;
wire _guard16447 = cond_wire309_out;
wire _guard16448 = _guard16446 & _guard16447;
wire _guard16449 = fsm_out == 1'd0;
wire _guard16450 = _guard16448 & _guard16449;
wire _guard16451 = _guard16445 | _guard16450;
wire _guard16452 = early_reset_static_par0_go_out;
wire _guard16453 = _guard16451 & _guard16452;
wire _guard16454 = fsm_out == 1'd0;
wire _guard16455 = cond_wire307_out;
wire _guard16456 = _guard16454 & _guard16455;
wire _guard16457 = fsm_out == 1'd0;
wire _guard16458 = _guard16456 & _guard16457;
wire _guard16459 = fsm_out == 1'd0;
wire _guard16460 = cond_wire309_out;
wire _guard16461 = _guard16459 & _guard16460;
wire _guard16462 = fsm_out == 1'd0;
wire _guard16463 = _guard16461 & _guard16462;
wire _guard16464 = _guard16458 | _guard16463;
wire _guard16465 = early_reset_static_par0_go_out;
wire _guard16466 = _guard16464 & _guard16465;
wire _guard16467 = fsm_out == 1'd0;
wire _guard16468 = cond_wire307_out;
wire _guard16469 = _guard16467 & _guard16468;
wire _guard16470 = fsm_out == 1'd0;
wire _guard16471 = _guard16469 & _guard16470;
wire _guard16472 = fsm_out == 1'd0;
wire _guard16473 = cond_wire309_out;
wire _guard16474 = _guard16472 & _guard16473;
wire _guard16475 = fsm_out == 1'd0;
wire _guard16476 = _guard16474 & _guard16475;
wire _guard16477 = _guard16471 | _guard16476;
wire _guard16478 = early_reset_static_par0_go_out;
wire _guard16479 = _guard16477 & _guard16478;
wire _guard16480 = cond_wire280_out;
wire _guard16481 = early_reset_static_par0_go_out;
wire _guard16482 = _guard16480 & _guard16481;
wire _guard16483 = cond_wire280_out;
wire _guard16484 = early_reset_static_par0_go_out;
wire _guard16485 = _guard16483 & _guard16484;
wire _guard16486 = cond_wire353_out;
wire _guard16487 = early_reset_static_par0_go_out;
wire _guard16488 = _guard16486 & _guard16487;
wire _guard16489 = cond_wire353_out;
wire _guard16490 = early_reset_static_par0_go_out;
wire _guard16491 = _guard16489 & _guard16490;
wire _guard16492 = cond_wire393_out;
wire _guard16493 = early_reset_static_par0_go_out;
wire _guard16494 = _guard16492 & _guard16493;
wire _guard16495 = cond_wire393_out;
wire _guard16496 = early_reset_static_par0_go_out;
wire _guard16497 = _guard16495 & _guard16496;
wire _guard16498 = cond_wire435_out;
wire _guard16499 = early_reset_static_par0_go_out;
wire _guard16500 = _guard16498 & _guard16499;
wire _guard16501 = cond_wire433_out;
wire _guard16502 = early_reset_static_par0_go_out;
wire _guard16503 = _guard16501 & _guard16502;
wire _guard16504 = fsm_out == 1'd0;
wire _guard16505 = cond_wire433_out;
wire _guard16506 = _guard16504 & _guard16505;
wire _guard16507 = fsm_out == 1'd0;
wire _guard16508 = _guard16506 & _guard16507;
wire _guard16509 = fsm_out == 1'd0;
wire _guard16510 = cond_wire435_out;
wire _guard16511 = _guard16509 & _guard16510;
wire _guard16512 = fsm_out == 1'd0;
wire _guard16513 = _guard16511 & _guard16512;
wire _guard16514 = _guard16508 | _guard16513;
wire _guard16515 = early_reset_static_par0_go_out;
wire _guard16516 = _guard16514 & _guard16515;
wire _guard16517 = fsm_out == 1'd0;
wire _guard16518 = cond_wire433_out;
wire _guard16519 = _guard16517 & _guard16518;
wire _guard16520 = fsm_out == 1'd0;
wire _guard16521 = _guard16519 & _guard16520;
wire _guard16522 = fsm_out == 1'd0;
wire _guard16523 = cond_wire435_out;
wire _guard16524 = _guard16522 & _guard16523;
wire _guard16525 = fsm_out == 1'd0;
wire _guard16526 = _guard16524 & _guard16525;
wire _guard16527 = _guard16521 | _guard16526;
wire _guard16528 = early_reset_static_par0_go_out;
wire _guard16529 = _guard16527 & _guard16528;
wire _guard16530 = fsm_out == 1'd0;
wire _guard16531 = cond_wire433_out;
wire _guard16532 = _guard16530 & _guard16531;
wire _guard16533 = fsm_out == 1'd0;
wire _guard16534 = _guard16532 & _guard16533;
wire _guard16535 = fsm_out == 1'd0;
wire _guard16536 = cond_wire435_out;
wire _guard16537 = _guard16535 & _guard16536;
wire _guard16538 = fsm_out == 1'd0;
wire _guard16539 = _guard16537 & _guard16538;
wire _guard16540 = _guard16534 | _guard16539;
wire _guard16541 = early_reset_static_par0_go_out;
wire _guard16542 = _guard16540 & _guard16541;
wire _guard16543 = cond_wire385_out;
wire _guard16544 = early_reset_static_par0_go_out;
wire _guard16545 = _guard16543 & _guard16544;
wire _guard16546 = cond_wire385_out;
wire _guard16547 = early_reset_static_par0_go_out;
wire _guard16548 = _guard16546 & _guard16547;
wire _guard16549 = cond_wire459_out;
wire _guard16550 = early_reset_static_par0_go_out;
wire _guard16551 = _guard16549 & _guard16550;
wire _guard16552 = cond_wire457_out;
wire _guard16553 = early_reset_static_par0_go_out;
wire _guard16554 = _guard16552 & _guard16553;
wire _guard16555 = fsm_out == 1'd0;
wire _guard16556 = cond_wire457_out;
wire _guard16557 = _guard16555 & _guard16556;
wire _guard16558 = fsm_out == 1'd0;
wire _guard16559 = _guard16557 & _guard16558;
wire _guard16560 = fsm_out == 1'd0;
wire _guard16561 = cond_wire459_out;
wire _guard16562 = _guard16560 & _guard16561;
wire _guard16563 = fsm_out == 1'd0;
wire _guard16564 = _guard16562 & _guard16563;
wire _guard16565 = _guard16559 | _guard16564;
wire _guard16566 = early_reset_static_par0_go_out;
wire _guard16567 = _guard16565 & _guard16566;
wire _guard16568 = fsm_out == 1'd0;
wire _guard16569 = cond_wire457_out;
wire _guard16570 = _guard16568 & _guard16569;
wire _guard16571 = fsm_out == 1'd0;
wire _guard16572 = _guard16570 & _guard16571;
wire _guard16573 = fsm_out == 1'd0;
wire _guard16574 = cond_wire459_out;
wire _guard16575 = _guard16573 & _guard16574;
wire _guard16576 = fsm_out == 1'd0;
wire _guard16577 = _guard16575 & _guard16576;
wire _guard16578 = _guard16572 | _guard16577;
wire _guard16579 = early_reset_static_par0_go_out;
wire _guard16580 = _guard16578 & _guard16579;
wire _guard16581 = fsm_out == 1'd0;
wire _guard16582 = cond_wire457_out;
wire _guard16583 = _guard16581 & _guard16582;
wire _guard16584 = fsm_out == 1'd0;
wire _guard16585 = _guard16583 & _guard16584;
wire _guard16586 = fsm_out == 1'd0;
wire _guard16587 = cond_wire459_out;
wire _guard16588 = _guard16586 & _guard16587;
wire _guard16589 = fsm_out == 1'd0;
wire _guard16590 = _guard16588 & _guard16589;
wire _guard16591 = _guard16585 | _guard16590;
wire _guard16592 = early_reset_static_par0_go_out;
wire _guard16593 = _guard16591 & _guard16592;
wire _guard16594 = cond_wire463_out;
wire _guard16595 = early_reset_static_par0_go_out;
wire _guard16596 = _guard16594 & _guard16595;
wire _guard16597 = cond_wire461_out;
wire _guard16598 = early_reset_static_par0_go_out;
wire _guard16599 = _guard16597 & _guard16598;
wire _guard16600 = fsm_out == 1'd0;
wire _guard16601 = cond_wire461_out;
wire _guard16602 = _guard16600 & _guard16601;
wire _guard16603 = fsm_out == 1'd0;
wire _guard16604 = _guard16602 & _guard16603;
wire _guard16605 = fsm_out == 1'd0;
wire _guard16606 = cond_wire463_out;
wire _guard16607 = _guard16605 & _guard16606;
wire _guard16608 = fsm_out == 1'd0;
wire _guard16609 = _guard16607 & _guard16608;
wire _guard16610 = _guard16604 | _guard16609;
wire _guard16611 = early_reset_static_par0_go_out;
wire _guard16612 = _guard16610 & _guard16611;
wire _guard16613 = fsm_out == 1'd0;
wire _guard16614 = cond_wire461_out;
wire _guard16615 = _guard16613 & _guard16614;
wire _guard16616 = fsm_out == 1'd0;
wire _guard16617 = _guard16615 & _guard16616;
wire _guard16618 = fsm_out == 1'd0;
wire _guard16619 = cond_wire463_out;
wire _guard16620 = _guard16618 & _guard16619;
wire _guard16621 = fsm_out == 1'd0;
wire _guard16622 = _guard16620 & _guard16621;
wire _guard16623 = _guard16617 | _guard16622;
wire _guard16624 = early_reset_static_par0_go_out;
wire _guard16625 = _guard16623 & _guard16624;
wire _guard16626 = fsm_out == 1'd0;
wire _guard16627 = cond_wire461_out;
wire _guard16628 = _guard16626 & _guard16627;
wire _guard16629 = fsm_out == 1'd0;
wire _guard16630 = _guard16628 & _guard16629;
wire _guard16631 = fsm_out == 1'd0;
wire _guard16632 = cond_wire463_out;
wire _guard16633 = _guard16631 & _guard16632;
wire _guard16634 = fsm_out == 1'd0;
wire _guard16635 = _guard16633 & _guard16634;
wire _guard16636 = _guard16630 | _guard16635;
wire _guard16637 = early_reset_static_par0_go_out;
wire _guard16638 = _guard16636 & _guard16637;
wire _guard16639 = cond_wire467_out;
wire _guard16640 = early_reset_static_par0_go_out;
wire _guard16641 = _guard16639 & _guard16640;
wire _guard16642 = cond_wire465_out;
wire _guard16643 = early_reset_static_par0_go_out;
wire _guard16644 = _guard16642 & _guard16643;
wire _guard16645 = fsm_out == 1'd0;
wire _guard16646 = cond_wire465_out;
wire _guard16647 = _guard16645 & _guard16646;
wire _guard16648 = fsm_out == 1'd0;
wire _guard16649 = _guard16647 & _guard16648;
wire _guard16650 = fsm_out == 1'd0;
wire _guard16651 = cond_wire467_out;
wire _guard16652 = _guard16650 & _guard16651;
wire _guard16653 = fsm_out == 1'd0;
wire _guard16654 = _guard16652 & _guard16653;
wire _guard16655 = _guard16649 | _guard16654;
wire _guard16656 = early_reset_static_par0_go_out;
wire _guard16657 = _guard16655 & _guard16656;
wire _guard16658 = fsm_out == 1'd0;
wire _guard16659 = cond_wire465_out;
wire _guard16660 = _guard16658 & _guard16659;
wire _guard16661 = fsm_out == 1'd0;
wire _guard16662 = _guard16660 & _guard16661;
wire _guard16663 = fsm_out == 1'd0;
wire _guard16664 = cond_wire467_out;
wire _guard16665 = _guard16663 & _guard16664;
wire _guard16666 = fsm_out == 1'd0;
wire _guard16667 = _guard16665 & _guard16666;
wire _guard16668 = _guard16662 | _guard16667;
wire _guard16669 = early_reset_static_par0_go_out;
wire _guard16670 = _guard16668 & _guard16669;
wire _guard16671 = fsm_out == 1'd0;
wire _guard16672 = cond_wire465_out;
wire _guard16673 = _guard16671 & _guard16672;
wire _guard16674 = fsm_out == 1'd0;
wire _guard16675 = _guard16673 & _guard16674;
wire _guard16676 = fsm_out == 1'd0;
wire _guard16677 = cond_wire467_out;
wire _guard16678 = _guard16676 & _guard16677;
wire _guard16679 = fsm_out == 1'd0;
wire _guard16680 = _guard16678 & _guard16679;
wire _guard16681 = _guard16675 | _guard16680;
wire _guard16682 = early_reset_static_par0_go_out;
wire _guard16683 = _guard16681 & _guard16682;
wire _guard16684 = cond_wire544_out;
wire _guard16685 = early_reset_static_par0_go_out;
wire _guard16686 = _guard16684 & _guard16685;
wire _guard16687 = cond_wire544_out;
wire _guard16688 = early_reset_static_par0_go_out;
wire _guard16689 = _guard16687 & _guard16688;
wire _guard16690 = cond_wire602_out;
wire _guard16691 = early_reset_static_par0_go_out;
wire _guard16692 = _guard16690 & _guard16691;
wire _guard16693 = cond_wire600_out;
wire _guard16694 = early_reset_static_par0_go_out;
wire _guard16695 = _guard16693 & _guard16694;
wire _guard16696 = fsm_out == 1'd0;
wire _guard16697 = cond_wire600_out;
wire _guard16698 = _guard16696 & _guard16697;
wire _guard16699 = fsm_out == 1'd0;
wire _guard16700 = _guard16698 & _guard16699;
wire _guard16701 = fsm_out == 1'd0;
wire _guard16702 = cond_wire602_out;
wire _guard16703 = _guard16701 & _guard16702;
wire _guard16704 = fsm_out == 1'd0;
wire _guard16705 = _guard16703 & _guard16704;
wire _guard16706 = _guard16700 | _guard16705;
wire _guard16707 = early_reset_static_par0_go_out;
wire _guard16708 = _guard16706 & _guard16707;
wire _guard16709 = fsm_out == 1'd0;
wire _guard16710 = cond_wire600_out;
wire _guard16711 = _guard16709 & _guard16710;
wire _guard16712 = fsm_out == 1'd0;
wire _guard16713 = _guard16711 & _guard16712;
wire _guard16714 = fsm_out == 1'd0;
wire _guard16715 = cond_wire602_out;
wire _guard16716 = _guard16714 & _guard16715;
wire _guard16717 = fsm_out == 1'd0;
wire _guard16718 = _guard16716 & _guard16717;
wire _guard16719 = _guard16713 | _guard16718;
wire _guard16720 = early_reset_static_par0_go_out;
wire _guard16721 = _guard16719 & _guard16720;
wire _guard16722 = fsm_out == 1'd0;
wire _guard16723 = cond_wire600_out;
wire _guard16724 = _guard16722 & _guard16723;
wire _guard16725 = fsm_out == 1'd0;
wire _guard16726 = _guard16724 & _guard16725;
wire _guard16727 = fsm_out == 1'd0;
wire _guard16728 = cond_wire602_out;
wire _guard16729 = _guard16727 & _guard16728;
wire _guard16730 = fsm_out == 1'd0;
wire _guard16731 = _guard16729 & _guard16730;
wire _guard16732 = _guard16726 | _guard16731;
wire _guard16733 = early_reset_static_par0_go_out;
wire _guard16734 = _guard16732 & _guard16733;
wire _guard16735 = cond_wire601_out;
wire _guard16736 = early_reset_static_par0_go_out;
wire _guard16737 = _guard16735 & _guard16736;
wire _guard16738 = cond_wire601_out;
wire _guard16739 = early_reset_static_par0_go_out;
wire _guard16740 = _guard16738 & _guard16739;
wire _guard16741 = cond_wire605_out;
wire _guard16742 = early_reset_static_par0_go_out;
wire _guard16743 = _guard16741 & _guard16742;
wire _guard16744 = cond_wire605_out;
wire _guard16745 = early_reset_static_par0_go_out;
wire _guard16746 = _guard16744 & _guard16745;
wire _guard16747 = cond_wire618_out;
wire _guard16748 = early_reset_static_par0_go_out;
wire _guard16749 = _guard16747 & _guard16748;
wire _guard16750 = cond_wire616_out;
wire _guard16751 = early_reset_static_par0_go_out;
wire _guard16752 = _guard16750 & _guard16751;
wire _guard16753 = fsm_out == 1'd0;
wire _guard16754 = cond_wire616_out;
wire _guard16755 = _guard16753 & _guard16754;
wire _guard16756 = fsm_out == 1'd0;
wire _guard16757 = _guard16755 & _guard16756;
wire _guard16758 = fsm_out == 1'd0;
wire _guard16759 = cond_wire618_out;
wire _guard16760 = _guard16758 & _guard16759;
wire _guard16761 = fsm_out == 1'd0;
wire _guard16762 = _guard16760 & _guard16761;
wire _guard16763 = _guard16757 | _guard16762;
wire _guard16764 = early_reset_static_par0_go_out;
wire _guard16765 = _guard16763 & _guard16764;
wire _guard16766 = fsm_out == 1'd0;
wire _guard16767 = cond_wire616_out;
wire _guard16768 = _guard16766 & _guard16767;
wire _guard16769 = fsm_out == 1'd0;
wire _guard16770 = _guard16768 & _guard16769;
wire _guard16771 = fsm_out == 1'd0;
wire _guard16772 = cond_wire618_out;
wire _guard16773 = _guard16771 & _guard16772;
wire _guard16774 = fsm_out == 1'd0;
wire _guard16775 = _guard16773 & _guard16774;
wire _guard16776 = _guard16770 | _guard16775;
wire _guard16777 = early_reset_static_par0_go_out;
wire _guard16778 = _guard16776 & _guard16777;
wire _guard16779 = fsm_out == 1'd0;
wire _guard16780 = cond_wire616_out;
wire _guard16781 = _guard16779 & _guard16780;
wire _guard16782 = fsm_out == 1'd0;
wire _guard16783 = _guard16781 & _guard16782;
wire _guard16784 = fsm_out == 1'd0;
wire _guard16785 = cond_wire618_out;
wire _guard16786 = _guard16784 & _guard16785;
wire _guard16787 = fsm_out == 1'd0;
wire _guard16788 = _guard16786 & _guard16787;
wire _guard16789 = _guard16783 | _guard16788;
wire _guard16790 = early_reset_static_par0_go_out;
wire _guard16791 = _guard16789 & _guard16790;
wire _guard16792 = cond_wire653_out;
wire _guard16793 = early_reset_static_par0_go_out;
wire _guard16794 = _guard16792 & _guard16793;
wire _guard16795 = cond_wire653_out;
wire _guard16796 = early_reset_static_par0_go_out;
wire _guard16797 = _guard16795 & _guard16796;
wire _guard16798 = cond_wire657_out;
wire _guard16799 = early_reset_static_par0_go_out;
wire _guard16800 = _guard16798 & _guard16799;
wire _guard16801 = cond_wire657_out;
wire _guard16802 = early_reset_static_par0_go_out;
wire _guard16803 = _guard16801 & _guard16802;
wire _guard16804 = cond_wire707_out;
wire _guard16805 = early_reset_static_par0_go_out;
wire _guard16806 = _guard16804 & _guard16805;
wire _guard16807 = cond_wire705_out;
wire _guard16808 = early_reset_static_par0_go_out;
wire _guard16809 = _guard16807 & _guard16808;
wire _guard16810 = fsm_out == 1'd0;
wire _guard16811 = cond_wire705_out;
wire _guard16812 = _guard16810 & _guard16811;
wire _guard16813 = fsm_out == 1'd0;
wire _guard16814 = _guard16812 & _guard16813;
wire _guard16815 = fsm_out == 1'd0;
wire _guard16816 = cond_wire707_out;
wire _guard16817 = _guard16815 & _guard16816;
wire _guard16818 = fsm_out == 1'd0;
wire _guard16819 = _guard16817 & _guard16818;
wire _guard16820 = _guard16814 | _guard16819;
wire _guard16821 = early_reset_static_par0_go_out;
wire _guard16822 = _guard16820 & _guard16821;
wire _guard16823 = fsm_out == 1'd0;
wire _guard16824 = cond_wire705_out;
wire _guard16825 = _guard16823 & _guard16824;
wire _guard16826 = fsm_out == 1'd0;
wire _guard16827 = _guard16825 & _guard16826;
wire _guard16828 = fsm_out == 1'd0;
wire _guard16829 = cond_wire707_out;
wire _guard16830 = _guard16828 & _guard16829;
wire _guard16831 = fsm_out == 1'd0;
wire _guard16832 = _guard16830 & _guard16831;
wire _guard16833 = _guard16827 | _guard16832;
wire _guard16834 = early_reset_static_par0_go_out;
wire _guard16835 = _guard16833 & _guard16834;
wire _guard16836 = fsm_out == 1'd0;
wire _guard16837 = cond_wire705_out;
wire _guard16838 = _guard16836 & _guard16837;
wire _guard16839 = fsm_out == 1'd0;
wire _guard16840 = _guard16838 & _guard16839;
wire _guard16841 = fsm_out == 1'd0;
wire _guard16842 = cond_wire707_out;
wire _guard16843 = _guard16841 & _guard16842;
wire _guard16844 = fsm_out == 1'd0;
wire _guard16845 = _guard16843 & _guard16844;
wire _guard16846 = _guard16840 | _guard16845;
wire _guard16847 = early_reset_static_par0_go_out;
wire _guard16848 = _guard16846 & _guard16847;
wire _guard16849 = cond_wire641_out;
wire _guard16850 = early_reset_static_par0_go_out;
wire _guard16851 = _guard16849 & _guard16850;
wire _guard16852 = cond_wire641_out;
wire _guard16853 = early_reset_static_par0_go_out;
wire _guard16854 = _guard16852 & _guard16853;
wire _guard16855 = cond_wire801_out;
wire _guard16856 = early_reset_static_par0_go_out;
wire _guard16857 = _guard16855 & _guard16856;
wire _guard16858 = cond_wire799_out;
wire _guard16859 = early_reset_static_par0_go_out;
wire _guard16860 = _guard16858 & _guard16859;
wire _guard16861 = fsm_out == 1'd0;
wire _guard16862 = cond_wire799_out;
wire _guard16863 = _guard16861 & _guard16862;
wire _guard16864 = fsm_out == 1'd0;
wire _guard16865 = _guard16863 & _guard16864;
wire _guard16866 = fsm_out == 1'd0;
wire _guard16867 = cond_wire801_out;
wire _guard16868 = _guard16866 & _guard16867;
wire _guard16869 = fsm_out == 1'd0;
wire _guard16870 = _guard16868 & _guard16869;
wire _guard16871 = _guard16865 | _guard16870;
wire _guard16872 = early_reset_static_par0_go_out;
wire _guard16873 = _guard16871 & _guard16872;
wire _guard16874 = fsm_out == 1'd0;
wire _guard16875 = cond_wire799_out;
wire _guard16876 = _guard16874 & _guard16875;
wire _guard16877 = fsm_out == 1'd0;
wire _guard16878 = _guard16876 & _guard16877;
wire _guard16879 = fsm_out == 1'd0;
wire _guard16880 = cond_wire801_out;
wire _guard16881 = _guard16879 & _guard16880;
wire _guard16882 = fsm_out == 1'd0;
wire _guard16883 = _guard16881 & _guard16882;
wire _guard16884 = _guard16878 | _guard16883;
wire _guard16885 = early_reset_static_par0_go_out;
wire _guard16886 = _guard16884 & _guard16885;
wire _guard16887 = fsm_out == 1'd0;
wire _guard16888 = cond_wire799_out;
wire _guard16889 = _guard16887 & _guard16888;
wire _guard16890 = fsm_out == 1'd0;
wire _guard16891 = _guard16889 & _guard16890;
wire _guard16892 = fsm_out == 1'd0;
wire _guard16893 = cond_wire801_out;
wire _guard16894 = _guard16892 & _guard16893;
wire _guard16895 = fsm_out == 1'd0;
wire _guard16896 = _guard16894 & _guard16895;
wire _guard16897 = _guard16891 | _guard16896;
wire _guard16898 = early_reset_static_par0_go_out;
wire _guard16899 = _guard16897 & _guard16898;
wire _guard16900 = cond_wire796_out;
wire _guard16901 = early_reset_static_par0_go_out;
wire _guard16902 = _guard16900 & _guard16901;
wire _guard16903 = cond_wire796_out;
wire _guard16904 = early_reset_static_par0_go_out;
wire _guard16905 = _guard16903 & _guard16904;
wire _guard16906 = cond_wire751_out;
wire _guard16907 = early_reset_static_par0_go_out;
wire _guard16908 = _guard16906 & _guard16907;
wire _guard16909 = cond_wire751_out;
wire _guard16910 = early_reset_static_par0_go_out;
wire _guard16911 = _guard16909 & _guard16910;
wire _guard16912 = cond_wire825_out;
wire _guard16913 = early_reset_static_par0_go_out;
wire _guard16914 = _guard16912 & _guard16913;
wire _guard16915 = cond_wire823_out;
wire _guard16916 = early_reset_static_par0_go_out;
wire _guard16917 = _guard16915 & _guard16916;
wire _guard16918 = fsm_out == 1'd0;
wire _guard16919 = cond_wire823_out;
wire _guard16920 = _guard16918 & _guard16919;
wire _guard16921 = fsm_out == 1'd0;
wire _guard16922 = _guard16920 & _guard16921;
wire _guard16923 = fsm_out == 1'd0;
wire _guard16924 = cond_wire825_out;
wire _guard16925 = _guard16923 & _guard16924;
wire _guard16926 = fsm_out == 1'd0;
wire _guard16927 = _guard16925 & _guard16926;
wire _guard16928 = _guard16922 | _guard16927;
wire _guard16929 = early_reset_static_par0_go_out;
wire _guard16930 = _guard16928 & _guard16929;
wire _guard16931 = fsm_out == 1'd0;
wire _guard16932 = cond_wire823_out;
wire _guard16933 = _guard16931 & _guard16932;
wire _guard16934 = fsm_out == 1'd0;
wire _guard16935 = _guard16933 & _guard16934;
wire _guard16936 = fsm_out == 1'd0;
wire _guard16937 = cond_wire825_out;
wire _guard16938 = _guard16936 & _guard16937;
wire _guard16939 = fsm_out == 1'd0;
wire _guard16940 = _guard16938 & _guard16939;
wire _guard16941 = _guard16935 | _guard16940;
wire _guard16942 = early_reset_static_par0_go_out;
wire _guard16943 = _guard16941 & _guard16942;
wire _guard16944 = fsm_out == 1'd0;
wire _guard16945 = cond_wire823_out;
wire _guard16946 = _guard16944 & _guard16945;
wire _guard16947 = fsm_out == 1'd0;
wire _guard16948 = _guard16946 & _guard16947;
wire _guard16949 = fsm_out == 1'd0;
wire _guard16950 = cond_wire825_out;
wire _guard16951 = _guard16949 & _guard16950;
wire _guard16952 = fsm_out == 1'd0;
wire _guard16953 = _guard16951 & _guard16952;
wire _guard16954 = _guard16948 | _guard16953;
wire _guard16955 = early_reset_static_par0_go_out;
wire _guard16956 = _guard16954 & _guard16955;
wire _guard16957 = cond_wire841_out;
wire _guard16958 = early_reset_static_par0_go_out;
wire _guard16959 = _guard16957 & _guard16958;
wire _guard16960 = cond_wire839_out;
wire _guard16961 = early_reset_static_par0_go_out;
wire _guard16962 = _guard16960 & _guard16961;
wire _guard16963 = fsm_out == 1'd0;
wire _guard16964 = cond_wire839_out;
wire _guard16965 = _guard16963 & _guard16964;
wire _guard16966 = fsm_out == 1'd0;
wire _guard16967 = _guard16965 & _guard16966;
wire _guard16968 = fsm_out == 1'd0;
wire _guard16969 = cond_wire841_out;
wire _guard16970 = _guard16968 & _guard16969;
wire _guard16971 = fsm_out == 1'd0;
wire _guard16972 = _guard16970 & _guard16971;
wire _guard16973 = _guard16967 | _guard16972;
wire _guard16974 = early_reset_static_par0_go_out;
wire _guard16975 = _guard16973 & _guard16974;
wire _guard16976 = fsm_out == 1'd0;
wire _guard16977 = cond_wire839_out;
wire _guard16978 = _guard16976 & _guard16977;
wire _guard16979 = fsm_out == 1'd0;
wire _guard16980 = _guard16978 & _guard16979;
wire _guard16981 = fsm_out == 1'd0;
wire _guard16982 = cond_wire841_out;
wire _guard16983 = _guard16981 & _guard16982;
wire _guard16984 = fsm_out == 1'd0;
wire _guard16985 = _guard16983 & _guard16984;
wire _guard16986 = _guard16980 | _guard16985;
wire _guard16987 = early_reset_static_par0_go_out;
wire _guard16988 = _guard16986 & _guard16987;
wire _guard16989 = fsm_out == 1'd0;
wire _guard16990 = cond_wire839_out;
wire _guard16991 = _guard16989 & _guard16990;
wire _guard16992 = fsm_out == 1'd0;
wire _guard16993 = _guard16991 & _guard16992;
wire _guard16994 = fsm_out == 1'd0;
wire _guard16995 = cond_wire841_out;
wire _guard16996 = _guard16994 & _guard16995;
wire _guard16997 = fsm_out == 1'd0;
wire _guard16998 = _guard16996 & _guard16997;
wire _guard16999 = _guard16993 | _guard16998;
wire _guard17000 = early_reset_static_par0_go_out;
wire _guard17001 = _guard16999 & _guard17000;
wire _guard17002 = cond_wire808_out;
wire _guard17003 = early_reset_static_par0_go_out;
wire _guard17004 = _guard17002 & _guard17003;
wire _guard17005 = cond_wire808_out;
wire _guard17006 = early_reset_static_par0_go_out;
wire _guard17007 = _guard17005 & _guard17006;
wire _guard17008 = cond_wire828_out;
wire _guard17009 = early_reset_static_par0_go_out;
wire _guard17010 = _guard17008 & _guard17009;
wire _guard17011 = cond_wire828_out;
wire _guard17012 = early_reset_static_par0_go_out;
wire _guard17013 = _guard17011 & _guard17012;
wire _guard17014 = cond_wire906_out;
wire _guard17015 = early_reset_static_par0_go_out;
wire _guard17016 = _guard17014 & _guard17015;
wire _guard17017 = cond_wire904_out;
wire _guard17018 = early_reset_static_par0_go_out;
wire _guard17019 = _guard17017 & _guard17018;
wire _guard17020 = fsm_out == 1'd0;
wire _guard17021 = cond_wire904_out;
wire _guard17022 = _guard17020 & _guard17021;
wire _guard17023 = fsm_out == 1'd0;
wire _guard17024 = _guard17022 & _guard17023;
wire _guard17025 = fsm_out == 1'd0;
wire _guard17026 = cond_wire906_out;
wire _guard17027 = _guard17025 & _guard17026;
wire _guard17028 = fsm_out == 1'd0;
wire _guard17029 = _guard17027 & _guard17028;
wire _guard17030 = _guard17024 | _guard17029;
wire _guard17031 = early_reset_static_par0_go_out;
wire _guard17032 = _guard17030 & _guard17031;
wire _guard17033 = fsm_out == 1'd0;
wire _guard17034 = cond_wire904_out;
wire _guard17035 = _guard17033 & _guard17034;
wire _guard17036 = fsm_out == 1'd0;
wire _guard17037 = _guard17035 & _guard17036;
wire _guard17038 = fsm_out == 1'd0;
wire _guard17039 = cond_wire906_out;
wire _guard17040 = _guard17038 & _guard17039;
wire _guard17041 = fsm_out == 1'd0;
wire _guard17042 = _guard17040 & _guard17041;
wire _guard17043 = _guard17037 | _guard17042;
wire _guard17044 = early_reset_static_par0_go_out;
wire _guard17045 = _guard17043 & _guard17044;
wire _guard17046 = fsm_out == 1'd0;
wire _guard17047 = cond_wire904_out;
wire _guard17048 = _guard17046 & _guard17047;
wire _guard17049 = fsm_out == 1'd0;
wire _guard17050 = _guard17048 & _guard17049;
wire _guard17051 = fsm_out == 1'd0;
wire _guard17052 = cond_wire906_out;
wire _guard17053 = _guard17051 & _guard17052;
wire _guard17054 = fsm_out == 1'd0;
wire _guard17055 = _guard17053 & _guard17054;
wire _guard17056 = _guard17050 | _guard17055;
wire _guard17057 = early_reset_static_par0_go_out;
wire _guard17058 = _guard17056 & _guard17057;
wire _guard17059 = cond_wire913_out;
wire _guard17060 = early_reset_static_par0_go_out;
wire _guard17061 = _guard17059 & _guard17060;
wire _guard17062 = cond_wire913_out;
wire _guard17063 = early_reset_static_par0_go_out;
wire _guard17064 = _guard17062 & _guard17063;
wire _guard17065 = cond_wire889_out;
wire _guard17066 = early_reset_static_par0_go_out;
wire _guard17067 = _guard17065 & _guard17066;
wire _guard17068 = cond_wire889_out;
wire _guard17069 = early_reset_static_par0_go_out;
wire _guard17070 = _guard17068 & _guard17069;
wire _guard17071 = cond_wire970_out;
wire _guard17072 = early_reset_static_par0_go_out;
wire _guard17073 = _guard17071 & _guard17072;
wire _guard17074 = cond_wire970_out;
wire _guard17075 = early_reset_static_par0_go_out;
wire _guard17076 = _guard17074 & _guard17075;
wire _guard17077 = cond_wire974_out;
wire _guard17078 = early_reset_static_par0_go_out;
wire _guard17079 = _guard17077 & _guard17078;
wire _guard17080 = cond_wire974_out;
wire _guard17081 = early_reset_static_par0_go_out;
wire _guard17082 = _guard17080 & _guard17081;
wire _guard17083 = cond_wire989_out;
wire _guard17084 = early_reset_static_par0_go_out;
wire _guard17085 = _guard17083 & _guard17084;
wire _guard17086 = cond_wire989_out;
wire _guard17087 = early_reset_static_par0_go_out;
wire _guard17088 = _guard17086 & _guard17087;
wire _guard17089 = cond_wire950_out;
wire _guard17090 = early_reset_static_par0_go_out;
wire _guard17091 = _guard17089 & _guard17090;
wire _guard17092 = cond_wire950_out;
wire _guard17093 = early_reset_static_par0_go_out;
wire _guard17094 = _guard17092 & _guard17093;
wire _guard17095 = cond_wire966_out;
wire _guard17096 = early_reset_static_par0_go_out;
wire _guard17097 = _guard17095 & _guard17096;
wire _guard17098 = cond_wire966_out;
wire _guard17099 = early_reset_static_par0_go_out;
wire _guard17100 = _guard17098 & _guard17099;
wire _guard17101 = cond_wire1036_out;
wire _guard17102 = early_reset_static_par0_go_out;
wire _guard17103 = _guard17101 & _guard17102;
wire _guard17104 = cond_wire1034_out;
wire _guard17105 = early_reset_static_par0_go_out;
wire _guard17106 = _guard17104 & _guard17105;
wire _guard17107 = fsm_out == 1'd0;
wire _guard17108 = cond_wire1034_out;
wire _guard17109 = _guard17107 & _guard17108;
wire _guard17110 = fsm_out == 1'd0;
wire _guard17111 = _guard17109 & _guard17110;
wire _guard17112 = fsm_out == 1'd0;
wire _guard17113 = cond_wire1036_out;
wire _guard17114 = _guard17112 & _guard17113;
wire _guard17115 = fsm_out == 1'd0;
wire _guard17116 = _guard17114 & _guard17115;
wire _guard17117 = _guard17111 | _guard17116;
wire _guard17118 = early_reset_static_par0_go_out;
wire _guard17119 = _guard17117 & _guard17118;
wire _guard17120 = fsm_out == 1'd0;
wire _guard17121 = cond_wire1034_out;
wire _guard17122 = _guard17120 & _guard17121;
wire _guard17123 = fsm_out == 1'd0;
wire _guard17124 = _guard17122 & _guard17123;
wire _guard17125 = fsm_out == 1'd0;
wire _guard17126 = cond_wire1036_out;
wire _guard17127 = _guard17125 & _guard17126;
wire _guard17128 = fsm_out == 1'd0;
wire _guard17129 = _guard17127 & _guard17128;
wire _guard17130 = _guard17124 | _guard17129;
wire _guard17131 = early_reset_static_par0_go_out;
wire _guard17132 = _guard17130 & _guard17131;
wire _guard17133 = fsm_out == 1'd0;
wire _guard17134 = cond_wire1034_out;
wire _guard17135 = _guard17133 & _guard17134;
wire _guard17136 = fsm_out == 1'd0;
wire _guard17137 = _guard17135 & _guard17136;
wire _guard17138 = fsm_out == 1'd0;
wire _guard17139 = cond_wire1036_out;
wire _guard17140 = _guard17138 & _guard17139;
wire _guard17141 = fsm_out == 1'd0;
wire _guard17142 = _guard17140 & _guard17141;
wire _guard17143 = _guard17137 | _guard17142;
wire _guard17144 = early_reset_static_par0_go_out;
wire _guard17145 = _guard17143 & _guard17144;
wire _guard17146 = cond_wire69_out;
wire _guard17147 = early_reset_static_par0_go_out;
wire _guard17148 = _guard17146 & _guard17147;
wire _guard17149 = cond_wire69_out;
wire _guard17150 = early_reset_static_par0_go_out;
wire _guard17151 = _guard17149 & _guard17150;
wire _guard17152 = cond_wire469_out;
wire _guard17153 = early_reset_static_par0_go_out;
wire _guard17154 = _guard17152 & _guard17153;
wire _guard17155 = cond_wire469_out;
wire _guard17156 = early_reset_static_par0_go_out;
wire _guard17157 = _guard17155 & _guard17156;
wire _guard17158 = cond_wire794_out;
wire _guard17159 = early_reset_static_par0_go_out;
wire _guard17160 = _guard17158 & _guard17159;
wire _guard17161 = cond_wire794_out;
wire _guard17162 = early_reset_static_par0_go_out;
wire _guard17163 = _guard17161 & _guard17162;
wire _guard17164 = early_reset_static_par0_go_out;
wire _guard17165 = early_reset_static_par0_go_out;
wire _guard17166 = early_reset_static_par0_go_out;
wire _guard17167 = early_reset_static_par0_go_out;
wire _guard17168 = early_reset_static_par0_go_out;
wire _guard17169 = early_reset_static_par0_go_out;
wire _guard17170 = fsm0_out == 6'd0;
wire _guard17171 = early_reset_static_seq_go_out;
wire _guard17172 = _guard17170 & _guard17171;
wire _guard17173 = early_reset_static_par0_go_out;
wire _guard17174 = _guard17172 | _guard17173;
wire _guard17175 = early_reset_static_par0_go_out;
wire _guard17176 = fsm0_out == 6'd0;
wire _guard17177 = early_reset_static_seq_go_out;
wire _guard17178 = _guard17176 & _guard17177;
wire _guard17179 = fsm0_out == 6'd0;
wire _guard17180 = early_reset_static_seq_go_out;
wire _guard17181 = _guard17179 & _guard17180;
wire _guard17182 = early_reset_static_par0_go_out;
wire _guard17183 = _guard17181 | _guard17182;
wire _guard17184 = early_reset_static_par0_go_out;
wire _guard17185 = fsm0_out == 6'd0;
wire _guard17186 = early_reset_static_seq_go_out;
wire _guard17187 = _guard17185 & _guard17186;
wire _guard17188 = early_reset_static_par0_go_out;
wire _guard17189 = early_reset_static_par0_go_out;
wire _guard17190 = early_reset_static_par0_go_out;
wire _guard17191 = early_reset_static_par0_go_out;
wire _guard17192 = early_reset_static_par0_go_out;
wire _guard17193 = early_reset_static_par0_go_out;
wire _guard17194 = early_reset_static_par0_go_out;
wire _guard17195 = early_reset_static_par0_go_out;
wire _guard17196 = fsm0_out == 6'd0;
wire _guard17197 = early_reset_static_seq_go_out;
wire _guard17198 = _guard17196 & _guard17197;
wire _guard17199 = early_reset_static_par0_go_out;
wire _guard17200 = _guard17198 | _guard17199;
wire _guard17201 = fsm0_out == 6'd0;
wire _guard17202 = early_reset_static_seq_go_out;
wire _guard17203 = _guard17201 & _guard17202;
wire _guard17204 = early_reset_static_par0_go_out;
wire _guard17205 = fsm0_out == 6'd0;
wire _guard17206 = early_reset_static_seq_go_out;
wire _guard17207 = _guard17205 & _guard17206;
wire _guard17208 = early_reset_static_par0_go_out;
wire _guard17209 = _guard17207 | _guard17208;
wire _guard17210 = early_reset_static_par0_go_out;
wire _guard17211 = fsm0_out == 6'd0;
wire _guard17212 = early_reset_static_seq_go_out;
wire _guard17213 = _guard17211 & _guard17212;
wire _guard17214 = early_reset_static_par0_go_out;
wire _guard17215 = early_reset_static_par0_go_out;
wire _guard17216 = early_reset_static_par0_go_out;
wire _guard17217 = early_reset_static_par0_go_out;
wire _guard17218 = early_reset_static_par0_go_out;
wire _guard17219 = early_reset_static_par0_go_out;
wire _guard17220 = fsm0_out == 6'd0;
wire _guard17221 = early_reset_static_seq_go_out;
wire _guard17222 = _guard17220 & _guard17221;
wire _guard17223 = early_reset_static_par0_go_out;
wire _guard17224 = _guard17222 | _guard17223;
wire _guard17225 = fsm0_out == 6'd0;
wire _guard17226 = early_reset_static_seq_go_out;
wire _guard17227 = _guard17225 & _guard17226;
wire _guard17228 = early_reset_static_par0_go_out;
wire _guard17229 = early_reset_static_par0_go_out;
wire _guard17230 = early_reset_static_par0_go_out;
wire _guard17231 = early_reset_static_par0_go_out;
wire _guard17232 = early_reset_static_par0_go_out;
wire _guard17233 = early_reset_static_par0_go_out;
wire _guard17234 = early_reset_static_par0_go_out;
wire _guard17235 = early_reset_static_par0_go_out;
wire _guard17236 = early_reset_static_par0_go_out;
wire _guard17237 = ~_guard0;
wire _guard17238 = early_reset_static_par0_go_out;
wire _guard17239 = _guard17237 & _guard17238;
wire _guard17240 = early_reset_static_par0_go_out;
wire _guard17241 = early_reset_static_par0_go_out;
wire _guard17242 = early_reset_static_par0_go_out;
wire _guard17243 = ~_guard0;
wire _guard17244 = early_reset_static_par0_go_out;
wire _guard17245 = _guard17243 & _guard17244;
wire _guard17246 = early_reset_static_par0_go_out;
wire _guard17247 = early_reset_static_par0_go_out;
wire _guard17248 = early_reset_static_par0_go_out;
wire _guard17249 = early_reset_static_par0_go_out;
wire _guard17250 = ~_guard0;
wire _guard17251 = early_reset_static_par0_go_out;
wire _guard17252 = _guard17250 & _guard17251;
wire _guard17253 = early_reset_static_par0_go_out;
wire _guard17254 = early_reset_static_par0_go_out;
wire _guard17255 = early_reset_static_par0_go_out;
wire _guard17256 = ~_guard0;
wire _guard17257 = early_reset_static_par0_go_out;
wire _guard17258 = _guard17256 & _guard17257;
wire _guard17259 = ~_guard0;
wire _guard17260 = early_reset_static_par0_go_out;
wire _guard17261 = _guard17259 & _guard17260;
wire _guard17262 = early_reset_static_par0_go_out;
wire _guard17263 = early_reset_static_par0_go_out;
wire _guard17264 = ~_guard0;
wire _guard17265 = early_reset_static_par0_go_out;
wire _guard17266 = _guard17264 & _guard17265;
wire _guard17267 = early_reset_static_par0_go_out;
wire _guard17268 = early_reset_static_par0_go_out;
wire _guard17269 = early_reset_static_par0_go_out;
wire _guard17270 = early_reset_static_par0_go_out;
wire _guard17271 = ~_guard0;
wire _guard17272 = early_reset_static_par0_go_out;
wire _guard17273 = _guard17271 & _guard17272;
wire _guard17274 = early_reset_static_par0_go_out;
wire _guard17275 = early_reset_static_par0_go_out;
wire _guard17276 = early_reset_static_par0_go_out;
wire _guard17277 = early_reset_static_par0_go_out;
wire _guard17278 = early_reset_static_par0_go_out;
wire _guard17279 = ~_guard0;
wire _guard17280 = early_reset_static_par0_go_out;
wire _guard17281 = _guard17279 & _guard17280;
wire _guard17282 = early_reset_static_par0_go_out;
wire _guard17283 = early_reset_static_par0_go_out;
wire _guard17284 = early_reset_static_par0_go_out;
wire _guard17285 = early_reset_static_par0_go_out;
wire _guard17286 = early_reset_static_par0_go_out;
wire _guard17287 = early_reset_static_par0_go_out;
wire _guard17288 = ~_guard0;
wire _guard17289 = early_reset_static_par0_go_out;
wire _guard17290 = _guard17288 & _guard17289;
wire _guard17291 = ~_guard0;
wire _guard17292 = early_reset_static_par0_go_out;
wire _guard17293 = _guard17291 & _guard17292;
wire _guard17294 = early_reset_static_par0_go_out;
wire _guard17295 = early_reset_static_par0_go_out;
wire _guard17296 = ~_guard0;
wire _guard17297 = early_reset_static_par0_go_out;
wire _guard17298 = _guard17296 & _guard17297;
wire _guard17299 = early_reset_static_par0_go_out;
wire _guard17300 = early_reset_static_par0_go_out;
wire _guard17301 = ~_guard0;
wire _guard17302 = early_reset_static_par0_go_out;
wire _guard17303 = _guard17301 & _guard17302;
wire _guard17304 = early_reset_static_par0_go_out;
wire _guard17305 = early_reset_static_par0_go_out;
wire _guard17306 = early_reset_static_par0_go_out;
wire _guard17307 = early_reset_static_par0_go_out;
wire _guard17308 = early_reset_static_par0_go_out;
wire _guard17309 = ~_guard0;
wire _guard17310 = early_reset_static_par0_go_out;
wire _guard17311 = _guard17309 & _guard17310;
wire _guard17312 = early_reset_static_par0_go_out;
wire _guard17313 = early_reset_static_par0_go_out;
wire _guard17314 = ~_guard0;
wire _guard17315 = early_reset_static_par0_go_out;
wire _guard17316 = _guard17314 & _guard17315;
wire _guard17317 = ~_guard0;
wire _guard17318 = early_reset_static_par0_go_out;
wire _guard17319 = _guard17317 & _guard17318;
wire _guard17320 = early_reset_static_par0_go_out;
wire _guard17321 = ~_guard0;
wire _guard17322 = early_reset_static_par0_go_out;
wire _guard17323 = _guard17321 & _guard17322;
wire _guard17324 = early_reset_static_par0_go_out;
wire _guard17325 = early_reset_static_par0_go_out;
wire _guard17326 = early_reset_static_par0_go_out;
wire _guard17327 = early_reset_static_par0_go_out;
wire _guard17328 = early_reset_static_par0_go_out;
wire _guard17329 = early_reset_static_par0_go_out;
wire _guard17330 = early_reset_static_par0_go_out;
wire _guard17331 = early_reset_static_par0_go_out;
wire _guard17332 = ~_guard0;
wire _guard17333 = early_reset_static_par0_go_out;
wire _guard17334 = _guard17332 & _guard17333;
wire _guard17335 = early_reset_static_par0_go_out;
wire _guard17336 = early_reset_static_par0_go_out;
wire _guard17337 = early_reset_static_par0_go_out;
wire _guard17338 = ~_guard0;
wire _guard17339 = early_reset_static_par0_go_out;
wire _guard17340 = _guard17338 & _guard17339;
wire _guard17341 = ~_guard0;
wire _guard17342 = early_reset_static_par0_go_out;
wire _guard17343 = _guard17341 & _guard17342;
wire _guard17344 = early_reset_static_par0_go_out;
wire _guard17345 = ~_guard0;
wire _guard17346 = early_reset_static_par0_go_out;
wire _guard17347 = _guard17345 & _guard17346;
wire _guard17348 = early_reset_static_par0_go_out;
wire _guard17349 = early_reset_static_par0_go_out;
wire _guard17350 = early_reset_static_par0_go_out;
wire _guard17351 = early_reset_static_par0_go_out;
wire _guard17352 = ~_guard0;
wire _guard17353 = early_reset_static_par0_go_out;
wire _guard17354 = _guard17352 & _guard17353;
wire _guard17355 = early_reset_static_par0_go_out;
wire _guard17356 = early_reset_static_par0_go_out;
wire _guard17357 = early_reset_static_par0_go_out;
wire _guard17358 = early_reset_static_par0_go_out;
wire _guard17359 = early_reset_static_par0_go_out;
wire _guard17360 = ~_guard0;
wire _guard17361 = early_reset_static_par0_go_out;
wire _guard17362 = _guard17360 & _guard17361;
wire _guard17363 = ~_guard0;
wire _guard17364 = early_reset_static_par0_go_out;
wire _guard17365 = _guard17363 & _guard17364;
wire _guard17366 = early_reset_static_par0_go_out;
wire _guard17367 = early_reset_static_par0_go_out;
wire _guard17368 = ~_guard0;
wire _guard17369 = early_reset_static_par0_go_out;
wire _guard17370 = _guard17368 & _guard17369;
wire _guard17371 = ~_guard0;
wire _guard17372 = early_reset_static_par0_go_out;
wire _guard17373 = _guard17371 & _guard17372;
wire _guard17374 = early_reset_static_par0_go_out;
wire _guard17375 = ~_guard0;
wire _guard17376 = early_reset_static_par0_go_out;
wire _guard17377 = _guard17375 & _guard17376;
wire _guard17378 = early_reset_static_par0_go_out;
wire _guard17379 = ~_guard0;
wire _guard17380 = early_reset_static_par0_go_out;
wire _guard17381 = _guard17379 & _guard17380;
wire _guard17382 = early_reset_static_par0_go_out;
wire _guard17383 = early_reset_static_par0_go_out;
wire _guard17384 = ~_guard0;
wire _guard17385 = early_reset_static_par0_go_out;
wire _guard17386 = _guard17384 & _guard17385;
wire _guard17387 = early_reset_static_par0_go_out;
wire _guard17388 = early_reset_static_par0_go_out;
wire _guard17389 = early_reset_static_par0_go_out;
wire _guard17390 = ~_guard0;
wire _guard17391 = early_reset_static_par0_go_out;
wire _guard17392 = _guard17390 & _guard17391;
wire _guard17393 = early_reset_static_par0_go_out;
wire _guard17394 = early_reset_static_par0_go_out;
wire _guard17395 = early_reset_static_par0_go_out;
wire _guard17396 = ~_guard0;
wire _guard17397 = early_reset_static_par0_go_out;
wire _guard17398 = _guard17396 & _guard17397;
wire _guard17399 = early_reset_static_par0_go_out;
wire _guard17400 = early_reset_static_par0_go_out;
wire _guard17401 = early_reset_static_par0_go_out;
wire _guard17402 = ~_guard0;
wire _guard17403 = early_reset_static_par0_go_out;
wire _guard17404 = _guard17402 & _guard17403;
wire _guard17405 = ~_guard0;
wire _guard17406 = early_reset_static_par0_go_out;
wire _guard17407 = _guard17405 & _guard17406;
wire _guard17408 = early_reset_static_par0_go_out;
wire _guard17409 = early_reset_static_par0_go_out;
wire _guard17410 = ~_guard0;
wire _guard17411 = early_reset_static_par0_go_out;
wire _guard17412 = _guard17410 & _guard17411;
wire _guard17413 = ~_guard0;
wire _guard17414 = early_reset_static_par0_go_out;
wire _guard17415 = _guard17413 & _guard17414;
wire _guard17416 = early_reset_static_par0_go_out;
wire _guard17417 = ~_guard0;
wire _guard17418 = early_reset_static_par0_go_out;
wire _guard17419 = _guard17417 & _guard17418;
wire _guard17420 = early_reset_static_par0_go_out;
wire _guard17421 = ~_guard0;
wire _guard17422 = early_reset_static_par0_go_out;
wire _guard17423 = _guard17421 & _guard17422;
wire _guard17424 = early_reset_static_par0_go_out;
wire _guard17425 = early_reset_static_par0_go_out;
wire _guard17426 = early_reset_static_par0_go_out;
wire _guard17427 = early_reset_static_par0_go_out;
wire _guard17428 = early_reset_static_par0_go_out;
wire _guard17429 = ~_guard0;
wire _guard17430 = early_reset_static_par0_go_out;
wire _guard17431 = _guard17429 & _guard17430;
wire _guard17432 = early_reset_static_par0_go_out;
wire _guard17433 = early_reset_static_par0_go_out;
wire _guard17434 = early_reset_static_par0_go_out;
wire _guard17435 = early_reset_static_par0_go_out;
wire _guard17436 = ~_guard0;
wire _guard17437 = early_reset_static_par0_go_out;
wire _guard17438 = _guard17436 & _guard17437;
wire _guard17439 = early_reset_static_par0_go_out;
wire _guard17440 = early_reset_static_par0_go_out;
wire _guard17441 = early_reset_static_par0_go_out;
wire _guard17442 = early_reset_static_par0_go_out;
wire _guard17443 = early_reset_static_par0_go_out;
wire _guard17444 = ~_guard0;
wire _guard17445 = early_reset_static_par0_go_out;
wire _guard17446 = _guard17444 & _guard17445;
wire _guard17447 = early_reset_static_par0_go_out;
wire _guard17448 = early_reset_static_par0_go_out;
wire _guard17449 = early_reset_static_par0_go_out;
wire _guard17450 = early_reset_static_par0_go_out;
wire _guard17451 = early_reset_static_par0_go_out;
wire _guard17452 = early_reset_static_par0_go_out;
wire _guard17453 = early_reset_static_par0_go_out;
wire _guard17454 = early_reset_static_par0_go_out;
wire _guard17455 = early_reset_static_par0_go_out;
wire _guard17456 = early_reset_static_par0_go_out;
wire _guard17457 = ~_guard0;
wire _guard17458 = early_reset_static_par0_go_out;
wire _guard17459 = _guard17457 & _guard17458;
wire _guard17460 = early_reset_static_par0_go_out;
wire _guard17461 = early_reset_static_par0_go_out;
wire _guard17462 = early_reset_static_par0_go_out;
wire _guard17463 = early_reset_static_par0_go_out;
wire _guard17464 = early_reset_static_par0_go_out;
wire _guard17465 = ~_guard0;
wire _guard17466 = early_reset_static_par0_go_out;
wire _guard17467 = _guard17465 & _guard17466;
wire _guard17468 = early_reset_static_par0_go_out;
wire _guard17469 = early_reset_static_par0_go_out;
wire _guard17470 = early_reset_static_par0_go_out;
wire _guard17471 = early_reset_static_par0_go_out;
wire _guard17472 = early_reset_static_par0_go_out;
wire _guard17473 = early_reset_static_par0_go_out;
wire _guard17474 = early_reset_static_par0_go_out;
wire _guard17475 = early_reset_static_par0_go_out;
wire _guard17476 = ~_guard0;
wire _guard17477 = early_reset_static_par0_go_out;
wire _guard17478 = _guard17476 & _guard17477;
wire _guard17479 = ~_guard0;
wire _guard17480 = early_reset_static_par0_go_out;
wire _guard17481 = _guard17479 & _guard17480;
wire _guard17482 = early_reset_static_par0_go_out;
wire _guard17483 = early_reset_static_par0_go_out;
wire _guard17484 = early_reset_static_par0_go_out;
wire _guard17485 = ~_guard0;
wire _guard17486 = early_reset_static_par0_go_out;
wire _guard17487 = _guard17485 & _guard17486;
wire _guard17488 = early_reset_static_par0_go_out;
wire _guard17489 = early_reset_static_par0_go_out;
wire _guard17490 = early_reset_static_par0_go_out;
wire _guard17491 = early_reset_static_par0_go_out;
wire _guard17492 = early_reset_static_par0_go_out;
wire _guard17493 = early_reset_static_par0_go_out;
wire _guard17494 = early_reset_static_par0_go_out;
wire _guard17495 = early_reset_static_par0_go_out;
wire _guard17496 = early_reset_static_par0_go_out;
wire _guard17497 = early_reset_static_par0_go_out;
wire _guard17498 = ~_guard0;
wire _guard17499 = early_reset_static_par0_go_out;
wire _guard17500 = _guard17498 & _guard17499;
wire _guard17501 = early_reset_static_par0_go_out;
wire _guard17502 = early_reset_static_par0_go_out;
wire _guard17503 = early_reset_static_par0_go_out;
wire _guard17504 = early_reset_static_par0_go_out;
wire _guard17505 = early_reset_static_par0_go_out;
wire _guard17506 = ~_guard0;
wire _guard17507 = early_reset_static_par0_go_out;
wire _guard17508 = _guard17506 & _guard17507;
wire _guard17509 = early_reset_static_par0_go_out;
wire _guard17510 = early_reset_static_par0_go_out;
wire _guard17511 = ~_guard0;
wire _guard17512 = early_reset_static_par0_go_out;
wire _guard17513 = _guard17511 & _guard17512;
wire _guard17514 = early_reset_static_par0_go_out;
wire _guard17515 = early_reset_static_par0_go_out;
wire _guard17516 = ~_guard0;
wire _guard17517 = early_reset_static_par0_go_out;
wire _guard17518 = _guard17516 & _guard17517;
wire _guard17519 = ~_guard0;
wire _guard17520 = early_reset_static_par0_go_out;
wire _guard17521 = _guard17519 & _guard17520;
wire _guard17522 = early_reset_static_par0_go_out;
wire _guard17523 = early_reset_static_par0_go_out;
wire _guard17524 = ~_guard0;
wire _guard17525 = early_reset_static_par0_go_out;
wire _guard17526 = _guard17524 & _guard17525;
wire _guard17527 = early_reset_static_par0_go_out;
wire _guard17528 = ~_guard0;
wire _guard17529 = early_reset_static_par0_go_out;
wire _guard17530 = _guard17528 & _guard17529;
wire _guard17531 = early_reset_static_par0_go_out;
wire _guard17532 = early_reset_static_par0_go_out;
wire _guard17533 = early_reset_static_par0_go_out;
wire _guard17534 = ~_guard0;
wire _guard17535 = early_reset_static_par0_go_out;
wire _guard17536 = _guard17534 & _guard17535;
wire _guard17537 = early_reset_static_par0_go_out;
wire _guard17538 = ~_guard0;
wire _guard17539 = early_reset_static_par0_go_out;
wire _guard17540 = _guard17538 & _guard17539;
wire _guard17541 = early_reset_static_par0_go_out;
wire _guard17542 = early_reset_static_par0_go_out;
wire _guard17543 = early_reset_static_par0_go_out;
wire _guard17544 = early_reset_static_par0_go_out;
wire _guard17545 = ~_guard0;
wire _guard17546 = early_reset_static_par0_go_out;
wire _guard17547 = _guard17545 & _guard17546;
wire _guard17548 = early_reset_static_par0_go_out;
wire _guard17549 = ~_guard0;
wire _guard17550 = early_reset_static_par0_go_out;
wire _guard17551 = _guard17549 & _guard17550;
wire _guard17552 = early_reset_static_par0_go_out;
wire _guard17553 = ~_guard0;
wire _guard17554 = early_reset_static_par0_go_out;
wire _guard17555 = _guard17553 & _guard17554;
wire _guard17556 = early_reset_static_par0_go_out;
wire _guard17557 = early_reset_static_par0_go_out;
wire _guard17558 = early_reset_static_par0_go_out;
wire _guard17559 = early_reset_static_par0_go_out;
wire _guard17560 = ~_guard0;
wire _guard17561 = early_reset_static_par0_go_out;
wire _guard17562 = _guard17560 & _guard17561;
wire _guard17563 = ~_guard0;
wire _guard17564 = early_reset_static_par0_go_out;
wire _guard17565 = _guard17563 & _guard17564;
wire _guard17566 = early_reset_static_par0_go_out;
wire _guard17567 = early_reset_static_par0_go_out;
wire _guard17568 = early_reset_static_par0_go_out;
wire _guard17569 = early_reset_static_par0_go_out;
wire _guard17570 = early_reset_static_par0_go_out;
wire _guard17571 = early_reset_static_par0_go_out;
wire _guard17572 = early_reset_static_par0_go_out;
wire _guard17573 = ~_guard0;
wire _guard17574 = early_reset_static_par0_go_out;
wire _guard17575 = _guard17573 & _guard17574;
wire _guard17576 = early_reset_static_par0_go_out;
wire _guard17577 = early_reset_static_par0_go_out;
wire _guard17578 = ~_guard0;
wire _guard17579 = early_reset_static_par0_go_out;
wire _guard17580 = _guard17578 & _guard17579;
wire _guard17581 = early_reset_static_par0_go_out;
wire _guard17582 = ~_guard0;
wire _guard17583 = early_reset_static_par0_go_out;
wire _guard17584 = _guard17582 & _guard17583;
wire _guard17585 = early_reset_static_par0_go_out;
wire _guard17586 = early_reset_static_par0_go_out;
wire _guard17587 = early_reset_static_par0_go_out;
wire _guard17588 = ~_guard0;
wire _guard17589 = early_reset_static_par0_go_out;
wire _guard17590 = _guard17588 & _guard17589;
wire _guard17591 = early_reset_static_par0_go_out;
wire _guard17592 = early_reset_static_par0_go_out;
wire _guard17593 = early_reset_static_par0_go_out;
wire _guard17594 = early_reset_static_par0_go_out;
wire _guard17595 = early_reset_static_par0_go_out;
wire _guard17596 = ~_guard0;
wire _guard17597 = early_reset_static_par0_go_out;
wire _guard17598 = _guard17596 & _guard17597;
wire _guard17599 = early_reset_static_par0_go_out;
wire _guard17600 = early_reset_static_par0_go_out;
wire _guard17601 = early_reset_static_par0_go_out;
wire _guard17602 = early_reset_static_par0_go_out;
wire _guard17603 = ~_guard0;
wire _guard17604 = early_reset_static_par0_go_out;
wire _guard17605 = _guard17603 & _guard17604;
wire _guard17606 = early_reset_static_par0_go_out;
wire _guard17607 = early_reset_static_par0_go_out;
wire _guard17608 = early_reset_static_par0_go_out;
wire _guard17609 = early_reset_static_par0_go_out;
wire _guard17610 = early_reset_static_par0_go_out;
wire _guard17611 = ~_guard0;
wire _guard17612 = early_reset_static_par0_go_out;
wire _guard17613 = _guard17611 & _guard17612;
wire _guard17614 = early_reset_static_par0_go_out;
wire _guard17615 = ~_guard0;
wire _guard17616 = early_reset_static_par0_go_out;
wire _guard17617 = _guard17615 & _guard17616;
wire _guard17618 = early_reset_static_par0_go_out;
wire _guard17619 = ~_guard0;
wire _guard17620 = early_reset_static_par0_go_out;
wire _guard17621 = _guard17619 & _guard17620;
wire _guard17622 = early_reset_static_par0_go_out;
wire _guard17623 = early_reset_static_par0_go_out;
wire _guard17624 = early_reset_static_par0_go_out;
wire _guard17625 = early_reset_static_par0_go_out;
wire _guard17626 = early_reset_static_par0_go_out;
wire _guard17627 = early_reset_static_par0_go_out;
wire _guard17628 = early_reset_static_par0_go_out;
wire _guard17629 = early_reset_static_par0_go_out;
wire _guard17630 = early_reset_static_par0_go_out;
wire _guard17631 = early_reset_static_par0_go_out;
wire _guard17632 = ~_guard0;
wire _guard17633 = early_reset_static_par0_go_out;
wire _guard17634 = _guard17632 & _guard17633;
wire _guard17635 = early_reset_static_par0_go_out;
wire _guard17636 = early_reset_static_par0_go_out;
wire _guard17637 = ~_guard0;
wire _guard17638 = early_reset_static_par0_go_out;
wire _guard17639 = _guard17637 & _guard17638;
wire _guard17640 = early_reset_static_par0_go_out;
wire _guard17641 = early_reset_static_par0_go_out;
wire _guard17642 = early_reset_static_par0_go_out;
wire _guard17643 = early_reset_static_par0_go_out;
wire _guard17644 = early_reset_static_par0_go_out;
wire _guard17645 = ~_guard0;
wire _guard17646 = early_reset_static_par0_go_out;
wire _guard17647 = _guard17645 & _guard17646;
wire _guard17648 = early_reset_static_par0_go_out;
wire _guard17649 = early_reset_static_par0_go_out;
wire _guard17650 = ~_guard0;
wire _guard17651 = early_reset_static_par0_go_out;
wire _guard17652 = _guard17650 & _guard17651;
wire _guard17653 = early_reset_static_par0_go_out;
wire _guard17654 = early_reset_static_par0_go_out;
wire _guard17655 = early_reset_static_par0_go_out;
wire _guard17656 = ~_guard0;
wire _guard17657 = early_reset_static_par0_go_out;
wire _guard17658 = _guard17656 & _guard17657;
wire _guard17659 = early_reset_static_par0_go_out;
wire _guard17660 = ~_guard0;
wire _guard17661 = early_reset_static_par0_go_out;
wire _guard17662 = _guard17660 & _guard17661;
wire _guard17663 = early_reset_static_par0_go_out;
wire _guard17664 = ~_guard0;
wire _guard17665 = early_reset_static_par0_go_out;
wire _guard17666 = _guard17664 & _guard17665;
wire _guard17667 = ~_guard0;
wire _guard17668 = early_reset_static_par0_go_out;
wire _guard17669 = _guard17667 & _guard17668;
wire _guard17670 = early_reset_static_par0_go_out;
wire _guard17671 = early_reset_static_par0_go_out;
wire _guard17672 = early_reset_static_par0_go_out;
wire _guard17673 = early_reset_static_par0_go_out;
wire _guard17674 = ~_guard0;
wire _guard17675 = early_reset_static_par0_go_out;
wire _guard17676 = _guard17674 & _guard17675;
wire _guard17677 = early_reset_static_par0_go_out;
wire _guard17678 = early_reset_static_par0_go_out;
wire _guard17679 = early_reset_static_par0_go_out;
wire _guard17680 = early_reset_static_par0_go_out;
wire _guard17681 = early_reset_static_par0_go_out;
wire _guard17682 = ~_guard0;
wire _guard17683 = early_reset_static_par0_go_out;
wire _guard17684 = _guard17682 & _guard17683;
wire _guard17685 = early_reset_static_par0_go_out;
wire _guard17686 = ~_guard0;
wire _guard17687 = early_reset_static_par0_go_out;
wire _guard17688 = _guard17686 & _guard17687;
wire _guard17689 = early_reset_static_par0_go_out;
wire _guard17690 = early_reset_static_par0_go_out;
wire _guard17691 = ~_guard0;
wire _guard17692 = early_reset_static_par0_go_out;
wire _guard17693 = _guard17691 & _guard17692;
wire _guard17694 = early_reset_static_par0_go_out;
wire _guard17695 = ~_guard0;
wire _guard17696 = early_reset_static_par0_go_out;
wire _guard17697 = _guard17695 & _guard17696;
wire _guard17698 = early_reset_static_par0_go_out;
wire _guard17699 = early_reset_static_par0_go_out;
wire _guard17700 = early_reset_static_par0_go_out;
wire _guard17701 = ~_guard0;
wire _guard17702 = early_reset_static_par0_go_out;
wire _guard17703 = _guard17701 & _guard17702;
wire _guard17704 = early_reset_static_par0_go_out;
wire _guard17705 = early_reset_static_par0_go_out;
wire _guard17706 = early_reset_static_par0_go_out;
wire _guard17707 = early_reset_static_par0_go_out;
wire _guard17708 = ~_guard0;
wire _guard17709 = early_reset_static_par0_go_out;
wire _guard17710 = _guard17708 & _guard17709;
wire _guard17711 = early_reset_static_par0_go_out;
wire _guard17712 = early_reset_static_par0_go_out;
wire _guard17713 = wrapper_early_reset_static_seq_go_out;
wire _guard17714 = cond_wire9_out;
wire _guard17715 = early_reset_static_par0_go_out;
wire _guard17716 = _guard17714 & _guard17715;
wire _guard17717 = cond_wire9_out;
wire _guard17718 = early_reset_static_par0_go_out;
wire _guard17719 = _guard17717 & _guard17718;
wire _guard17720 = cond_wire36_out;
wire _guard17721 = early_reset_static_par0_go_out;
wire _guard17722 = _guard17720 & _guard17721;
wire _guard17723 = cond_wire36_out;
wire _guard17724 = early_reset_static_par0_go_out;
wire _guard17725 = _guard17723 & _guard17724;
wire _guard17726 = cond_wire57_out;
wire _guard17727 = early_reset_static_par0_go_out;
wire _guard17728 = _guard17726 & _guard17727;
wire _guard17729 = cond_wire55_out;
wire _guard17730 = early_reset_static_par0_go_out;
wire _guard17731 = _guard17729 & _guard17730;
wire _guard17732 = fsm_out == 1'd0;
wire _guard17733 = cond_wire55_out;
wire _guard17734 = _guard17732 & _guard17733;
wire _guard17735 = fsm_out == 1'd0;
wire _guard17736 = _guard17734 & _guard17735;
wire _guard17737 = fsm_out == 1'd0;
wire _guard17738 = cond_wire57_out;
wire _guard17739 = _guard17737 & _guard17738;
wire _guard17740 = fsm_out == 1'd0;
wire _guard17741 = _guard17739 & _guard17740;
wire _guard17742 = _guard17736 | _guard17741;
wire _guard17743 = early_reset_static_par0_go_out;
wire _guard17744 = _guard17742 & _guard17743;
wire _guard17745 = fsm_out == 1'd0;
wire _guard17746 = cond_wire55_out;
wire _guard17747 = _guard17745 & _guard17746;
wire _guard17748 = fsm_out == 1'd0;
wire _guard17749 = _guard17747 & _guard17748;
wire _guard17750 = fsm_out == 1'd0;
wire _guard17751 = cond_wire57_out;
wire _guard17752 = _guard17750 & _guard17751;
wire _guard17753 = fsm_out == 1'd0;
wire _guard17754 = _guard17752 & _guard17753;
wire _guard17755 = _guard17749 | _guard17754;
wire _guard17756 = early_reset_static_par0_go_out;
wire _guard17757 = _guard17755 & _guard17756;
wire _guard17758 = fsm_out == 1'd0;
wire _guard17759 = cond_wire55_out;
wire _guard17760 = _guard17758 & _guard17759;
wire _guard17761 = fsm_out == 1'd0;
wire _guard17762 = _guard17760 & _guard17761;
wire _guard17763 = fsm_out == 1'd0;
wire _guard17764 = cond_wire57_out;
wire _guard17765 = _guard17763 & _guard17764;
wire _guard17766 = fsm_out == 1'd0;
wire _guard17767 = _guard17765 & _guard17766;
wire _guard17768 = _guard17762 | _guard17767;
wire _guard17769 = early_reset_static_par0_go_out;
wire _guard17770 = _guard17768 & _guard17769;
wire _guard17771 = cond_wire66_out;
wire _guard17772 = early_reset_static_par0_go_out;
wire _guard17773 = _guard17771 & _guard17772;
wire _guard17774 = cond_wire66_out;
wire _guard17775 = early_reset_static_par0_go_out;
wire _guard17776 = _guard17774 & _guard17775;
wire _guard17777 = cond_wire6_out;
wire _guard17778 = early_reset_static_par0_go_out;
wire _guard17779 = _guard17777 & _guard17778;
wire _guard17780 = cond_wire6_out;
wire _guard17781 = early_reset_static_par0_go_out;
wire _guard17782 = _guard17780 & _guard17781;
wire _guard17783 = cond_wire215_out;
wire _guard17784 = early_reset_static_par0_go_out;
wire _guard17785 = _guard17783 & _guard17784;
wire _guard17786 = cond_wire215_out;
wire _guard17787 = early_reset_static_par0_go_out;
wire _guard17788 = _guard17786 & _guard17787;
wire _guard17789 = cond_wire223_out;
wire _guard17790 = early_reset_static_par0_go_out;
wire _guard17791 = _guard17789 & _guard17790;
wire _guard17792 = cond_wire223_out;
wire _guard17793 = early_reset_static_par0_go_out;
wire _guard17794 = _guard17792 & _guard17793;
wire _guard17795 = cond_wire215_out;
wire _guard17796 = early_reset_static_par0_go_out;
wire _guard17797 = _guard17795 & _guard17796;
wire _guard17798 = cond_wire215_out;
wire _guard17799 = early_reset_static_par0_go_out;
wire _guard17800 = _guard17798 & _guard17799;
wire _guard17801 = cond_wire219_out;
wire _guard17802 = early_reset_static_par0_go_out;
wire _guard17803 = _guard17801 & _guard17802;
wire _guard17804 = cond_wire219_out;
wire _guard17805 = early_reset_static_par0_go_out;
wire _guard17806 = _guard17804 & _guard17805;
wire _guard17807 = cond_wire332_out;
wire _guard17808 = early_reset_static_par0_go_out;
wire _guard17809 = _guard17807 & _guard17808;
wire _guard17810 = cond_wire332_out;
wire _guard17811 = early_reset_static_par0_go_out;
wire _guard17812 = _guard17810 & _guard17811;
wire _guard17813 = cond_wire312_out;
wire _guard17814 = early_reset_static_par0_go_out;
wire _guard17815 = _guard17813 & _guard17814;
wire _guard17816 = cond_wire312_out;
wire _guard17817 = early_reset_static_par0_go_out;
wire _guard17818 = _guard17816 & _guard17817;
wire _guard17819 = cond_wire320_out;
wire _guard17820 = early_reset_static_par0_go_out;
wire _guard17821 = _guard17819 & _guard17820;
wire _guard17822 = cond_wire320_out;
wire _guard17823 = early_reset_static_par0_go_out;
wire _guard17824 = _guard17822 & _guard17823;
wire _guard17825 = cond_wire357_out;
wire _guard17826 = early_reset_static_par0_go_out;
wire _guard17827 = _guard17825 & _guard17826;
wire _guard17828 = cond_wire357_out;
wire _guard17829 = early_reset_static_par0_go_out;
wire _guard17830 = _guard17828 & _guard17829;
wire _guard17831 = cond_wire361_out;
wire _guard17832 = early_reset_static_par0_go_out;
wire _guard17833 = _guard17831 & _guard17832;
wire _guard17834 = cond_wire361_out;
wire _guard17835 = early_reset_static_par0_go_out;
wire _guard17836 = _guard17834 & _guard17835;
wire _guard17837 = cond_wire426_out;
wire _guard17838 = early_reset_static_par0_go_out;
wire _guard17839 = _guard17837 & _guard17838;
wire _guard17840 = cond_wire426_out;
wire _guard17841 = early_reset_static_par0_go_out;
wire _guard17842 = _guard17840 & _guard17841;
wire _guard17843 = cond_wire475_out;
wire _guard17844 = early_reset_static_par0_go_out;
wire _guard17845 = _guard17843 & _guard17844;
wire _guard17846 = cond_wire475_out;
wire _guard17847 = early_reset_static_par0_go_out;
wire _guard17848 = _guard17846 & _guard17847;
wire _guard17849 = cond_wire492_out;
wire _guard17850 = early_reset_static_par0_go_out;
wire _guard17851 = _guard17849 & _guard17850;
wire _guard17852 = cond_wire490_out;
wire _guard17853 = early_reset_static_par0_go_out;
wire _guard17854 = _guard17852 & _guard17853;
wire _guard17855 = fsm_out == 1'd0;
wire _guard17856 = cond_wire490_out;
wire _guard17857 = _guard17855 & _guard17856;
wire _guard17858 = fsm_out == 1'd0;
wire _guard17859 = _guard17857 & _guard17858;
wire _guard17860 = fsm_out == 1'd0;
wire _guard17861 = cond_wire492_out;
wire _guard17862 = _guard17860 & _guard17861;
wire _guard17863 = fsm_out == 1'd0;
wire _guard17864 = _guard17862 & _guard17863;
wire _guard17865 = _guard17859 | _guard17864;
wire _guard17866 = early_reset_static_par0_go_out;
wire _guard17867 = _guard17865 & _guard17866;
wire _guard17868 = fsm_out == 1'd0;
wire _guard17869 = cond_wire490_out;
wire _guard17870 = _guard17868 & _guard17869;
wire _guard17871 = fsm_out == 1'd0;
wire _guard17872 = _guard17870 & _guard17871;
wire _guard17873 = fsm_out == 1'd0;
wire _guard17874 = cond_wire492_out;
wire _guard17875 = _guard17873 & _guard17874;
wire _guard17876 = fsm_out == 1'd0;
wire _guard17877 = _guard17875 & _guard17876;
wire _guard17878 = _guard17872 | _guard17877;
wire _guard17879 = early_reset_static_par0_go_out;
wire _guard17880 = _guard17878 & _guard17879;
wire _guard17881 = fsm_out == 1'd0;
wire _guard17882 = cond_wire490_out;
wire _guard17883 = _guard17881 & _guard17882;
wire _guard17884 = fsm_out == 1'd0;
wire _guard17885 = _guard17883 & _guard17884;
wire _guard17886 = fsm_out == 1'd0;
wire _guard17887 = cond_wire492_out;
wire _guard17888 = _guard17886 & _guard17887;
wire _guard17889 = fsm_out == 1'd0;
wire _guard17890 = _guard17888 & _guard17889;
wire _guard17891 = _guard17885 | _guard17890;
wire _guard17892 = early_reset_static_par0_go_out;
wire _guard17893 = _guard17891 & _guard17892;
wire _guard17894 = cond_wire496_out;
wire _guard17895 = early_reset_static_par0_go_out;
wire _guard17896 = _guard17894 & _guard17895;
wire _guard17897 = cond_wire494_out;
wire _guard17898 = early_reset_static_par0_go_out;
wire _guard17899 = _guard17897 & _guard17898;
wire _guard17900 = fsm_out == 1'd0;
wire _guard17901 = cond_wire494_out;
wire _guard17902 = _guard17900 & _guard17901;
wire _guard17903 = fsm_out == 1'd0;
wire _guard17904 = _guard17902 & _guard17903;
wire _guard17905 = fsm_out == 1'd0;
wire _guard17906 = cond_wire496_out;
wire _guard17907 = _guard17905 & _guard17906;
wire _guard17908 = fsm_out == 1'd0;
wire _guard17909 = _guard17907 & _guard17908;
wire _guard17910 = _guard17904 | _guard17909;
wire _guard17911 = early_reset_static_par0_go_out;
wire _guard17912 = _guard17910 & _guard17911;
wire _guard17913 = fsm_out == 1'd0;
wire _guard17914 = cond_wire494_out;
wire _guard17915 = _guard17913 & _guard17914;
wire _guard17916 = fsm_out == 1'd0;
wire _guard17917 = _guard17915 & _guard17916;
wire _guard17918 = fsm_out == 1'd0;
wire _guard17919 = cond_wire496_out;
wire _guard17920 = _guard17918 & _guard17919;
wire _guard17921 = fsm_out == 1'd0;
wire _guard17922 = _guard17920 & _guard17921;
wire _guard17923 = _guard17917 | _guard17922;
wire _guard17924 = early_reset_static_par0_go_out;
wire _guard17925 = _guard17923 & _guard17924;
wire _guard17926 = fsm_out == 1'd0;
wire _guard17927 = cond_wire494_out;
wire _guard17928 = _guard17926 & _guard17927;
wire _guard17929 = fsm_out == 1'd0;
wire _guard17930 = _guard17928 & _guard17929;
wire _guard17931 = fsm_out == 1'd0;
wire _guard17932 = cond_wire496_out;
wire _guard17933 = _guard17931 & _guard17932;
wire _guard17934 = fsm_out == 1'd0;
wire _guard17935 = _guard17933 & _guard17934;
wire _guard17936 = _guard17930 | _guard17935;
wire _guard17937 = early_reset_static_par0_go_out;
wire _guard17938 = _guard17936 & _guard17937;
wire _guard17939 = cond_wire438_out;
wire _guard17940 = early_reset_static_par0_go_out;
wire _guard17941 = _guard17939 & _guard17940;
wire _guard17942 = cond_wire438_out;
wire _guard17943 = early_reset_static_par0_go_out;
wire _guard17944 = _guard17942 & _guard17943;
wire _guard17945 = cond_wire528_out;
wire _guard17946 = early_reset_static_par0_go_out;
wire _guard17947 = _guard17945 & _guard17946;
wire _guard17948 = cond_wire526_out;
wire _guard17949 = early_reset_static_par0_go_out;
wire _guard17950 = _guard17948 & _guard17949;
wire _guard17951 = fsm_out == 1'd0;
wire _guard17952 = cond_wire526_out;
wire _guard17953 = _guard17951 & _guard17952;
wire _guard17954 = fsm_out == 1'd0;
wire _guard17955 = _guard17953 & _guard17954;
wire _guard17956 = fsm_out == 1'd0;
wire _guard17957 = cond_wire528_out;
wire _guard17958 = _guard17956 & _guard17957;
wire _guard17959 = fsm_out == 1'd0;
wire _guard17960 = _guard17958 & _guard17959;
wire _guard17961 = _guard17955 | _guard17960;
wire _guard17962 = early_reset_static_par0_go_out;
wire _guard17963 = _guard17961 & _guard17962;
wire _guard17964 = fsm_out == 1'd0;
wire _guard17965 = cond_wire526_out;
wire _guard17966 = _guard17964 & _guard17965;
wire _guard17967 = fsm_out == 1'd0;
wire _guard17968 = _guard17966 & _guard17967;
wire _guard17969 = fsm_out == 1'd0;
wire _guard17970 = cond_wire528_out;
wire _guard17971 = _guard17969 & _guard17970;
wire _guard17972 = fsm_out == 1'd0;
wire _guard17973 = _guard17971 & _guard17972;
wire _guard17974 = _guard17968 | _guard17973;
wire _guard17975 = early_reset_static_par0_go_out;
wire _guard17976 = _guard17974 & _guard17975;
wire _guard17977 = fsm_out == 1'd0;
wire _guard17978 = cond_wire526_out;
wire _guard17979 = _guard17977 & _guard17978;
wire _guard17980 = fsm_out == 1'd0;
wire _guard17981 = _guard17979 & _guard17980;
wire _guard17982 = fsm_out == 1'd0;
wire _guard17983 = cond_wire528_out;
wire _guard17984 = _guard17982 & _guard17983;
wire _guard17985 = fsm_out == 1'd0;
wire _guard17986 = _guard17984 & _guard17985;
wire _guard17987 = _guard17981 | _guard17986;
wire _guard17988 = early_reset_static_par0_go_out;
wire _guard17989 = _guard17987 & _guard17988;
wire _guard17990 = cond_wire581_out;
wire _guard17991 = early_reset_static_par0_go_out;
wire _guard17992 = _guard17990 & _guard17991;
wire _guard17993 = cond_wire579_out;
wire _guard17994 = early_reset_static_par0_go_out;
wire _guard17995 = _guard17993 & _guard17994;
wire _guard17996 = fsm_out == 1'd0;
wire _guard17997 = cond_wire579_out;
wire _guard17998 = _guard17996 & _guard17997;
wire _guard17999 = fsm_out == 1'd0;
wire _guard18000 = _guard17998 & _guard17999;
wire _guard18001 = fsm_out == 1'd0;
wire _guard18002 = cond_wire581_out;
wire _guard18003 = _guard18001 & _guard18002;
wire _guard18004 = fsm_out == 1'd0;
wire _guard18005 = _guard18003 & _guard18004;
wire _guard18006 = _guard18000 | _guard18005;
wire _guard18007 = early_reset_static_par0_go_out;
wire _guard18008 = _guard18006 & _guard18007;
wire _guard18009 = fsm_out == 1'd0;
wire _guard18010 = cond_wire579_out;
wire _guard18011 = _guard18009 & _guard18010;
wire _guard18012 = fsm_out == 1'd0;
wire _guard18013 = _guard18011 & _guard18012;
wire _guard18014 = fsm_out == 1'd0;
wire _guard18015 = cond_wire581_out;
wire _guard18016 = _guard18014 & _guard18015;
wire _guard18017 = fsm_out == 1'd0;
wire _guard18018 = _guard18016 & _guard18017;
wire _guard18019 = _guard18013 | _guard18018;
wire _guard18020 = early_reset_static_par0_go_out;
wire _guard18021 = _guard18019 & _guard18020;
wire _guard18022 = fsm_out == 1'd0;
wire _guard18023 = cond_wire579_out;
wire _guard18024 = _guard18022 & _guard18023;
wire _guard18025 = fsm_out == 1'd0;
wire _guard18026 = _guard18024 & _guard18025;
wire _guard18027 = fsm_out == 1'd0;
wire _guard18028 = cond_wire581_out;
wire _guard18029 = _guard18027 & _guard18028;
wire _guard18030 = fsm_out == 1'd0;
wire _guard18031 = _guard18029 & _guard18030;
wire _guard18032 = _guard18026 | _guard18031;
wire _guard18033 = early_reset_static_par0_go_out;
wire _guard18034 = _guard18032 & _guard18033;
wire _guard18035 = cond_wire531_out;
wire _guard18036 = early_reset_static_par0_go_out;
wire _guard18037 = _guard18035 & _guard18036;
wire _guard18038 = cond_wire531_out;
wire _guard18039 = early_reset_static_par0_go_out;
wire _guard18040 = _guard18038 & _guard18039;
wire _guard18041 = cond_wire622_out;
wire _guard18042 = early_reset_static_par0_go_out;
wire _guard18043 = _guard18041 & _guard18042;
wire _guard18044 = cond_wire620_out;
wire _guard18045 = early_reset_static_par0_go_out;
wire _guard18046 = _guard18044 & _guard18045;
wire _guard18047 = fsm_out == 1'd0;
wire _guard18048 = cond_wire620_out;
wire _guard18049 = _guard18047 & _guard18048;
wire _guard18050 = fsm_out == 1'd0;
wire _guard18051 = _guard18049 & _guard18050;
wire _guard18052 = fsm_out == 1'd0;
wire _guard18053 = cond_wire622_out;
wire _guard18054 = _guard18052 & _guard18053;
wire _guard18055 = fsm_out == 1'd0;
wire _guard18056 = _guard18054 & _guard18055;
wire _guard18057 = _guard18051 | _guard18056;
wire _guard18058 = early_reset_static_par0_go_out;
wire _guard18059 = _guard18057 & _guard18058;
wire _guard18060 = fsm_out == 1'd0;
wire _guard18061 = cond_wire620_out;
wire _guard18062 = _guard18060 & _guard18061;
wire _guard18063 = fsm_out == 1'd0;
wire _guard18064 = _guard18062 & _guard18063;
wire _guard18065 = fsm_out == 1'd0;
wire _guard18066 = cond_wire622_out;
wire _guard18067 = _guard18065 & _guard18066;
wire _guard18068 = fsm_out == 1'd0;
wire _guard18069 = _guard18067 & _guard18068;
wire _guard18070 = _guard18064 | _guard18069;
wire _guard18071 = early_reset_static_par0_go_out;
wire _guard18072 = _guard18070 & _guard18071;
wire _guard18073 = fsm_out == 1'd0;
wire _guard18074 = cond_wire620_out;
wire _guard18075 = _guard18073 & _guard18074;
wire _guard18076 = fsm_out == 1'd0;
wire _guard18077 = _guard18075 & _guard18076;
wire _guard18078 = fsm_out == 1'd0;
wire _guard18079 = cond_wire622_out;
wire _guard18080 = _guard18078 & _guard18079;
wire _guard18081 = fsm_out == 1'd0;
wire _guard18082 = _guard18080 & _guard18081;
wire _guard18083 = _guard18077 | _guard18082;
wire _guard18084 = early_reset_static_par0_go_out;
wire _guard18085 = _guard18083 & _guard18084;
wire _guard18086 = cond_wire629_out;
wire _guard18087 = early_reset_static_par0_go_out;
wire _guard18088 = _guard18086 & _guard18087;
wire _guard18089 = cond_wire629_out;
wire _guard18090 = early_reset_static_par0_go_out;
wire _guard18091 = _guard18089 & _guard18090;
wire _guard18092 = cond_wire675_out;
wire _guard18093 = early_reset_static_par0_go_out;
wire _guard18094 = _guard18092 & _guard18093;
wire _guard18095 = cond_wire673_out;
wire _guard18096 = early_reset_static_par0_go_out;
wire _guard18097 = _guard18095 & _guard18096;
wire _guard18098 = fsm_out == 1'd0;
wire _guard18099 = cond_wire673_out;
wire _guard18100 = _guard18098 & _guard18099;
wire _guard18101 = fsm_out == 1'd0;
wire _guard18102 = _guard18100 & _guard18101;
wire _guard18103 = fsm_out == 1'd0;
wire _guard18104 = cond_wire675_out;
wire _guard18105 = _guard18103 & _guard18104;
wire _guard18106 = fsm_out == 1'd0;
wire _guard18107 = _guard18105 & _guard18106;
wire _guard18108 = _guard18102 | _guard18107;
wire _guard18109 = early_reset_static_par0_go_out;
wire _guard18110 = _guard18108 & _guard18109;
wire _guard18111 = fsm_out == 1'd0;
wire _guard18112 = cond_wire673_out;
wire _guard18113 = _guard18111 & _guard18112;
wire _guard18114 = fsm_out == 1'd0;
wire _guard18115 = _guard18113 & _guard18114;
wire _guard18116 = fsm_out == 1'd0;
wire _guard18117 = cond_wire675_out;
wire _guard18118 = _guard18116 & _guard18117;
wire _guard18119 = fsm_out == 1'd0;
wire _guard18120 = _guard18118 & _guard18119;
wire _guard18121 = _guard18115 | _guard18120;
wire _guard18122 = early_reset_static_par0_go_out;
wire _guard18123 = _guard18121 & _guard18122;
wire _guard18124 = fsm_out == 1'd0;
wire _guard18125 = cond_wire673_out;
wire _guard18126 = _guard18124 & _guard18125;
wire _guard18127 = fsm_out == 1'd0;
wire _guard18128 = _guard18126 & _guard18127;
wire _guard18129 = fsm_out == 1'd0;
wire _guard18130 = cond_wire675_out;
wire _guard18131 = _guard18129 & _guard18130;
wire _guard18132 = fsm_out == 1'd0;
wire _guard18133 = _guard18131 & _guard18132;
wire _guard18134 = _guard18128 | _guard18133;
wire _guard18135 = early_reset_static_par0_go_out;
wire _guard18136 = _guard18134 & _guard18135;
wire _guard18137 = cond_wire690_out;
wire _guard18138 = early_reset_static_par0_go_out;
wire _guard18139 = _guard18137 & _guard18138;
wire _guard18140 = cond_wire690_out;
wire _guard18141 = early_reset_static_par0_go_out;
wire _guard18142 = _guard18140 & _guard18141;
wire _guard18143 = cond_wire736_out;
wire _guard18144 = early_reset_static_par0_go_out;
wire _guard18145 = _guard18143 & _guard18144;
wire _guard18146 = cond_wire734_out;
wire _guard18147 = early_reset_static_par0_go_out;
wire _guard18148 = _guard18146 & _guard18147;
wire _guard18149 = fsm_out == 1'd0;
wire _guard18150 = cond_wire734_out;
wire _guard18151 = _guard18149 & _guard18150;
wire _guard18152 = fsm_out == 1'd0;
wire _guard18153 = _guard18151 & _guard18152;
wire _guard18154 = fsm_out == 1'd0;
wire _guard18155 = cond_wire736_out;
wire _guard18156 = _guard18154 & _guard18155;
wire _guard18157 = fsm_out == 1'd0;
wire _guard18158 = _guard18156 & _guard18157;
wire _guard18159 = _guard18153 | _guard18158;
wire _guard18160 = early_reset_static_par0_go_out;
wire _guard18161 = _guard18159 & _guard18160;
wire _guard18162 = fsm_out == 1'd0;
wire _guard18163 = cond_wire734_out;
wire _guard18164 = _guard18162 & _guard18163;
wire _guard18165 = fsm_out == 1'd0;
wire _guard18166 = _guard18164 & _guard18165;
wire _guard18167 = fsm_out == 1'd0;
wire _guard18168 = cond_wire736_out;
wire _guard18169 = _guard18167 & _guard18168;
wire _guard18170 = fsm_out == 1'd0;
wire _guard18171 = _guard18169 & _guard18170;
wire _guard18172 = _guard18166 | _guard18171;
wire _guard18173 = early_reset_static_par0_go_out;
wire _guard18174 = _guard18172 & _guard18173;
wire _guard18175 = fsm_out == 1'd0;
wire _guard18176 = cond_wire734_out;
wire _guard18177 = _guard18175 & _guard18176;
wire _guard18178 = fsm_out == 1'd0;
wire _guard18179 = _guard18177 & _guard18178;
wire _guard18180 = fsm_out == 1'd0;
wire _guard18181 = cond_wire736_out;
wire _guard18182 = _guard18180 & _guard18181;
wire _guard18183 = fsm_out == 1'd0;
wire _guard18184 = _guard18182 & _guard18183;
wire _guard18185 = _guard18179 | _guard18184;
wire _guard18186 = early_reset_static_par0_go_out;
wire _guard18187 = _guard18185 & _guard18186;
wire _guard18188 = cond_wire718_out;
wire _guard18189 = early_reset_static_par0_go_out;
wire _guard18190 = _guard18188 & _guard18189;
wire _guard18191 = cond_wire718_out;
wire _guard18192 = early_reset_static_par0_go_out;
wire _guard18193 = _guard18191 & _guard18192;
wire _guard18194 = cond_wire783_out;
wire _guard18195 = early_reset_static_par0_go_out;
wire _guard18196 = _guard18194 & _guard18195;
wire _guard18197 = cond_wire783_out;
wire _guard18198 = early_reset_static_par0_go_out;
wire _guard18199 = _guard18197 & _guard18198;
wire _guard18200 = cond_wire821_out;
wire _guard18201 = early_reset_static_par0_go_out;
wire _guard18202 = _guard18200 & _guard18201;
wire _guard18203 = cond_wire819_out;
wire _guard18204 = early_reset_static_par0_go_out;
wire _guard18205 = _guard18203 & _guard18204;
wire _guard18206 = fsm_out == 1'd0;
wire _guard18207 = cond_wire819_out;
wire _guard18208 = _guard18206 & _guard18207;
wire _guard18209 = fsm_out == 1'd0;
wire _guard18210 = _guard18208 & _guard18209;
wire _guard18211 = fsm_out == 1'd0;
wire _guard18212 = cond_wire821_out;
wire _guard18213 = _guard18211 & _guard18212;
wire _guard18214 = fsm_out == 1'd0;
wire _guard18215 = _guard18213 & _guard18214;
wire _guard18216 = _guard18210 | _guard18215;
wire _guard18217 = early_reset_static_par0_go_out;
wire _guard18218 = _guard18216 & _guard18217;
wire _guard18219 = fsm_out == 1'd0;
wire _guard18220 = cond_wire819_out;
wire _guard18221 = _guard18219 & _guard18220;
wire _guard18222 = fsm_out == 1'd0;
wire _guard18223 = _guard18221 & _guard18222;
wire _guard18224 = fsm_out == 1'd0;
wire _guard18225 = cond_wire821_out;
wire _guard18226 = _guard18224 & _guard18225;
wire _guard18227 = fsm_out == 1'd0;
wire _guard18228 = _guard18226 & _guard18227;
wire _guard18229 = _guard18223 | _guard18228;
wire _guard18230 = early_reset_static_par0_go_out;
wire _guard18231 = _guard18229 & _guard18230;
wire _guard18232 = fsm_out == 1'd0;
wire _guard18233 = cond_wire819_out;
wire _guard18234 = _guard18232 & _guard18233;
wire _guard18235 = fsm_out == 1'd0;
wire _guard18236 = _guard18234 & _guard18235;
wire _guard18237 = fsm_out == 1'd0;
wire _guard18238 = cond_wire821_out;
wire _guard18239 = _guard18237 & _guard18238;
wire _guard18240 = fsm_out == 1'd0;
wire _guard18241 = _guard18239 & _guard18240;
wire _guard18242 = _guard18236 | _guard18241;
wire _guard18243 = early_reset_static_par0_go_out;
wire _guard18244 = _guard18242 & _guard18243;
wire _guard18245 = cond_wire755_out;
wire _guard18246 = early_reset_static_par0_go_out;
wire _guard18247 = _guard18245 & _guard18246;
wire _guard18248 = cond_wire755_out;
wire _guard18249 = early_reset_static_par0_go_out;
wire _guard18250 = _guard18248 & _guard18249;
wire _guard18251 = cond_wire763_out;
wire _guard18252 = early_reset_static_par0_go_out;
wire _guard18253 = _guard18251 & _guard18252;
wire _guard18254 = cond_wire763_out;
wire _guard18255 = early_reset_static_par0_go_out;
wire _guard18256 = _guard18254 & _guard18255;
wire _guard18257 = cond_wire852_out;
wire _guard18258 = early_reset_static_par0_go_out;
wire _guard18259 = _guard18257 & _guard18258;
wire _guard18260 = cond_wire852_out;
wire _guard18261 = early_reset_static_par0_go_out;
wire _guard18262 = _guard18260 & _guard18261;
wire _guard18263 = cond_wire878_out;
wire _guard18264 = early_reset_static_par0_go_out;
wire _guard18265 = _guard18263 & _guard18264;
wire _guard18266 = cond_wire876_out;
wire _guard18267 = early_reset_static_par0_go_out;
wire _guard18268 = _guard18266 & _guard18267;
wire _guard18269 = fsm_out == 1'd0;
wire _guard18270 = cond_wire876_out;
wire _guard18271 = _guard18269 & _guard18270;
wire _guard18272 = fsm_out == 1'd0;
wire _guard18273 = _guard18271 & _guard18272;
wire _guard18274 = fsm_out == 1'd0;
wire _guard18275 = cond_wire878_out;
wire _guard18276 = _guard18274 & _guard18275;
wire _guard18277 = fsm_out == 1'd0;
wire _guard18278 = _guard18276 & _guard18277;
wire _guard18279 = _guard18273 | _guard18278;
wire _guard18280 = early_reset_static_par0_go_out;
wire _guard18281 = _guard18279 & _guard18280;
wire _guard18282 = fsm_out == 1'd0;
wire _guard18283 = cond_wire876_out;
wire _guard18284 = _guard18282 & _guard18283;
wire _guard18285 = fsm_out == 1'd0;
wire _guard18286 = _guard18284 & _guard18285;
wire _guard18287 = fsm_out == 1'd0;
wire _guard18288 = cond_wire878_out;
wire _guard18289 = _guard18287 & _guard18288;
wire _guard18290 = fsm_out == 1'd0;
wire _guard18291 = _guard18289 & _guard18290;
wire _guard18292 = _guard18286 | _guard18291;
wire _guard18293 = early_reset_static_par0_go_out;
wire _guard18294 = _guard18292 & _guard18293;
wire _guard18295 = fsm_out == 1'd0;
wire _guard18296 = cond_wire876_out;
wire _guard18297 = _guard18295 & _guard18296;
wire _guard18298 = fsm_out == 1'd0;
wire _guard18299 = _guard18297 & _guard18298;
wire _guard18300 = fsm_out == 1'd0;
wire _guard18301 = cond_wire878_out;
wire _guard18302 = _guard18300 & _guard18301;
wire _guard18303 = fsm_out == 1'd0;
wire _guard18304 = _guard18302 & _guard18303;
wire _guard18305 = _guard18299 | _guard18304;
wire _guard18306 = early_reset_static_par0_go_out;
wire _guard18307 = _guard18305 & _guard18306;
wire _guard18308 = cond_wire840_out;
wire _guard18309 = early_reset_static_par0_go_out;
wire _guard18310 = _guard18308 & _guard18309;
wire _guard18311 = cond_wire840_out;
wire _guard18312 = early_reset_static_par0_go_out;
wire _guard18313 = _guard18311 & _guard18312;
wire _guard18314 = cond_wire848_out;
wire _guard18315 = early_reset_static_par0_go_out;
wire _guard18316 = _guard18314 & _guard18315;
wire _guard18317 = cond_wire848_out;
wire _guard18318 = early_reset_static_par0_go_out;
wire _guard18319 = _guard18317 & _guard18318;
wire _guard18320 = cond_wire951_out;
wire _guard18321 = early_reset_static_par0_go_out;
wire _guard18322 = _guard18320 & _guard18321;
wire _guard18323 = cond_wire949_out;
wire _guard18324 = early_reset_static_par0_go_out;
wire _guard18325 = _guard18323 & _guard18324;
wire _guard18326 = fsm_out == 1'd0;
wire _guard18327 = cond_wire949_out;
wire _guard18328 = _guard18326 & _guard18327;
wire _guard18329 = fsm_out == 1'd0;
wire _guard18330 = _guard18328 & _guard18329;
wire _guard18331 = fsm_out == 1'd0;
wire _guard18332 = cond_wire951_out;
wire _guard18333 = _guard18331 & _guard18332;
wire _guard18334 = fsm_out == 1'd0;
wire _guard18335 = _guard18333 & _guard18334;
wire _guard18336 = _guard18330 | _guard18335;
wire _guard18337 = early_reset_static_par0_go_out;
wire _guard18338 = _guard18336 & _guard18337;
wire _guard18339 = fsm_out == 1'd0;
wire _guard18340 = cond_wire949_out;
wire _guard18341 = _guard18339 & _guard18340;
wire _guard18342 = fsm_out == 1'd0;
wire _guard18343 = _guard18341 & _guard18342;
wire _guard18344 = fsm_out == 1'd0;
wire _guard18345 = cond_wire951_out;
wire _guard18346 = _guard18344 & _guard18345;
wire _guard18347 = fsm_out == 1'd0;
wire _guard18348 = _guard18346 & _guard18347;
wire _guard18349 = _guard18343 | _guard18348;
wire _guard18350 = early_reset_static_par0_go_out;
wire _guard18351 = _guard18349 & _guard18350;
wire _guard18352 = fsm_out == 1'd0;
wire _guard18353 = cond_wire949_out;
wire _guard18354 = _guard18352 & _guard18353;
wire _guard18355 = fsm_out == 1'd0;
wire _guard18356 = _guard18354 & _guard18355;
wire _guard18357 = fsm_out == 1'd0;
wire _guard18358 = cond_wire951_out;
wire _guard18359 = _guard18357 & _guard18358;
wire _guard18360 = fsm_out == 1'd0;
wire _guard18361 = _guard18359 & _guard18360;
wire _guard18362 = _guard18356 | _guard18361;
wire _guard18363 = early_reset_static_par0_go_out;
wire _guard18364 = _guard18362 & _guard18363;
wire _guard18365 = cond_wire1008_out;
wire _guard18366 = early_reset_static_par0_go_out;
wire _guard18367 = _guard18365 & _guard18366;
wire _guard18368 = cond_wire1006_out;
wire _guard18369 = early_reset_static_par0_go_out;
wire _guard18370 = _guard18368 & _guard18369;
wire _guard18371 = fsm_out == 1'd0;
wire _guard18372 = cond_wire1006_out;
wire _guard18373 = _guard18371 & _guard18372;
wire _guard18374 = fsm_out == 1'd0;
wire _guard18375 = _guard18373 & _guard18374;
wire _guard18376 = fsm_out == 1'd0;
wire _guard18377 = cond_wire1008_out;
wire _guard18378 = _guard18376 & _guard18377;
wire _guard18379 = fsm_out == 1'd0;
wire _guard18380 = _guard18378 & _guard18379;
wire _guard18381 = _guard18375 | _guard18380;
wire _guard18382 = early_reset_static_par0_go_out;
wire _guard18383 = _guard18381 & _guard18382;
wire _guard18384 = fsm_out == 1'd0;
wire _guard18385 = cond_wire1006_out;
wire _guard18386 = _guard18384 & _guard18385;
wire _guard18387 = fsm_out == 1'd0;
wire _guard18388 = _guard18386 & _guard18387;
wire _guard18389 = fsm_out == 1'd0;
wire _guard18390 = cond_wire1008_out;
wire _guard18391 = _guard18389 & _guard18390;
wire _guard18392 = fsm_out == 1'd0;
wire _guard18393 = _guard18391 & _guard18392;
wire _guard18394 = _guard18388 | _guard18393;
wire _guard18395 = early_reset_static_par0_go_out;
wire _guard18396 = _guard18394 & _guard18395;
wire _guard18397 = fsm_out == 1'd0;
wire _guard18398 = cond_wire1006_out;
wire _guard18399 = _guard18397 & _guard18398;
wire _guard18400 = fsm_out == 1'd0;
wire _guard18401 = _guard18399 & _guard18400;
wire _guard18402 = fsm_out == 1'd0;
wire _guard18403 = cond_wire1008_out;
wire _guard18404 = _guard18402 & _guard18403;
wire _guard18405 = fsm_out == 1'd0;
wire _guard18406 = _guard18404 & _guard18405;
wire _guard18407 = _guard18401 | _guard18406;
wire _guard18408 = early_reset_static_par0_go_out;
wire _guard18409 = _guard18407 & _guard18408;
wire _guard18410 = cond_wire1011_out;
wire _guard18411 = early_reset_static_par0_go_out;
wire _guard18412 = _guard18410 & _guard18411;
wire _guard18413 = cond_wire1011_out;
wire _guard18414 = early_reset_static_par0_go_out;
wire _guard18415 = _guard18413 & _guard18414;
wire _guard18416 = cond_wire982_out;
wire _guard18417 = early_reset_static_par0_go_out;
wire _guard18418 = _guard18416 & _guard18417;
wire _guard18419 = cond_wire982_out;
wire _guard18420 = early_reset_static_par0_go_out;
wire _guard18421 = _guard18419 & _guard18420;
wire _guard18422 = cond_wire_out;
wire _guard18423 = early_reset_static_par0_go_out;
wire _guard18424 = _guard18422 & _guard18423;
wire _guard18425 = cond_wire_out;
wire _guard18426 = early_reset_static_par0_go_out;
wire _guard18427 = _guard18425 & _guard18426;
wire _guard18428 = cond_wire_out;
wire _guard18429 = early_reset_static_par0_go_out;
wire _guard18430 = _guard18428 & _guard18429;
wire _guard18431 = cond_wire_out;
wire _guard18432 = early_reset_static_par0_go_out;
wire _guard18433 = _guard18431 & _guard18432;
wire _guard18434 = early_reset_static_par0_go_out;
wire _guard18435 = early_reset_static_par0_go_out;
wire _guard18436 = early_reset_static_par0_go_out;
wire _guard18437 = early_reset_static_par0_go_out;
wire _guard18438 = early_reset_static_par0_go_out;
wire _guard18439 = early_reset_static_par0_go_out;
wire _guard18440 = fsm0_out == 6'd0;
wire _guard18441 = early_reset_static_seq_go_out;
wire _guard18442 = _guard18440 & _guard18441;
wire _guard18443 = early_reset_static_par0_go_out;
wire _guard18444 = _guard18442 | _guard18443;
wire _guard18445 = early_reset_static_par0_go_out;
wire _guard18446 = fsm0_out == 6'd0;
wire _guard18447 = early_reset_static_seq_go_out;
wire _guard18448 = _guard18446 & _guard18447;
wire _guard18449 = early_reset_static_par0_go_out;
wire _guard18450 = early_reset_static_par0_go_out;
wire _guard18451 = early_reset_static_par0_go_out;
wire _guard18452 = early_reset_static_par0_go_out;
wire _guard18453 = fsm0_out == 6'd0;
wire _guard18454 = early_reset_static_seq_go_out;
wire _guard18455 = _guard18453 & _guard18454;
wire _guard18456 = early_reset_static_par0_go_out;
wire _guard18457 = _guard18455 | _guard18456;
wire _guard18458 = early_reset_static_par0_go_out;
wire _guard18459 = fsm0_out == 6'd0;
wire _guard18460 = early_reset_static_seq_go_out;
wire _guard18461 = _guard18459 & _guard18460;
wire _guard18462 = early_reset_static_par0_go_out;
wire _guard18463 = early_reset_static_par0_go_out;
wire _guard18464 = fsm0_out == 6'd0;
wire _guard18465 = early_reset_static_seq_go_out;
wire _guard18466 = _guard18464 & _guard18465;
wire _guard18467 = early_reset_static_par0_go_out;
wire _guard18468 = _guard18466 | _guard18467;
wire _guard18469 = early_reset_static_par0_go_out;
wire _guard18470 = fsm0_out == 6'd0;
wire _guard18471 = early_reset_static_seq_go_out;
wire _guard18472 = _guard18470 & _guard18471;
wire _guard18473 = early_reset_static_par0_go_out;
wire _guard18474 = early_reset_static_par0_go_out;
wire _guard18475 = early_reset_static_par0_go_out;
wire _guard18476 = early_reset_static_par0_go_out;
wire _guard18477 = early_reset_static_par0_go_out;
wire _guard18478 = early_reset_static_par0_go_out;
wire _guard18479 = early_reset_static_par0_go_out;
wire _guard18480 = early_reset_static_par0_go_out;
wire _guard18481 = fsm0_out == 6'd0;
wire _guard18482 = early_reset_static_seq_go_out;
wire _guard18483 = _guard18481 & _guard18482;
wire _guard18484 = early_reset_static_par0_go_out;
wire _guard18485 = _guard18483 | _guard18484;
wire _guard18486 = fsm0_out == 6'd0;
wire _guard18487 = early_reset_static_seq_go_out;
wire _guard18488 = _guard18486 & _guard18487;
wire _guard18489 = early_reset_static_par0_go_out;
wire _guard18490 = early_reset_static_par0_go_out;
wire _guard18491 = early_reset_static_par0_go_out;
wire _guard18492 = early_reset_static_par0_go_out;
wire _guard18493 = early_reset_static_par0_go_out;
wire _guard18494 = early_reset_static_par0_go_out;
wire _guard18495 = early_reset_static_par0_go_out;
wire _guard18496 = early_reset_static_par0_go_out;
wire _guard18497 = early_reset_static_par0_go_out;
wire _guard18498 = early_reset_static_par0_go_out;
wire _guard18499 = ~_guard0;
wire _guard18500 = early_reset_static_par0_go_out;
wire _guard18501 = _guard18499 & _guard18500;
wire _guard18502 = early_reset_static_par0_go_out;
wire _guard18503 = ~_guard0;
wire _guard18504 = early_reset_static_par0_go_out;
wire _guard18505 = _guard18503 & _guard18504;
wire _guard18506 = early_reset_static_par0_go_out;
wire _guard18507 = early_reset_static_par0_go_out;
wire _guard18508 = ~_guard0;
wire _guard18509 = early_reset_static_par0_go_out;
wire _guard18510 = _guard18508 & _guard18509;
wire _guard18511 = early_reset_static_par0_go_out;
wire _guard18512 = early_reset_static_par0_go_out;
wire _guard18513 = early_reset_static_par0_go_out;
wire _guard18514 = early_reset_static_par0_go_out;
wire _guard18515 = early_reset_static_par0_go_out;
wire _guard18516 = early_reset_static_par0_go_out;
wire _guard18517 = early_reset_static_par0_go_out;
wire _guard18518 = early_reset_static_par0_go_out;
wire _guard18519 = early_reset_static_par0_go_out;
wire _guard18520 = ~_guard0;
wire _guard18521 = early_reset_static_par0_go_out;
wire _guard18522 = _guard18520 & _guard18521;
wire _guard18523 = early_reset_static_par0_go_out;
wire _guard18524 = ~_guard0;
wire _guard18525 = early_reset_static_par0_go_out;
wire _guard18526 = _guard18524 & _guard18525;
wire _guard18527 = early_reset_static_par0_go_out;
wire _guard18528 = early_reset_static_par0_go_out;
wire _guard18529 = early_reset_static_par0_go_out;
wire _guard18530 = early_reset_static_par0_go_out;
wire _guard18531 = ~_guard0;
wire _guard18532 = early_reset_static_par0_go_out;
wire _guard18533 = _guard18531 & _guard18532;
wire _guard18534 = early_reset_static_par0_go_out;
wire _guard18535 = ~_guard0;
wire _guard18536 = early_reset_static_par0_go_out;
wire _guard18537 = _guard18535 & _guard18536;
wire _guard18538 = early_reset_static_par0_go_out;
wire _guard18539 = early_reset_static_par0_go_out;
wire _guard18540 = early_reset_static_par0_go_out;
wire _guard18541 = early_reset_static_par0_go_out;
wire _guard18542 = ~_guard0;
wire _guard18543 = early_reset_static_par0_go_out;
wire _guard18544 = _guard18542 & _guard18543;
wire _guard18545 = early_reset_static_par0_go_out;
wire _guard18546 = early_reset_static_par0_go_out;
wire _guard18547 = early_reset_static_par0_go_out;
wire _guard18548 = early_reset_static_par0_go_out;
wire _guard18549 = early_reset_static_par0_go_out;
wire _guard18550 = ~_guard0;
wire _guard18551 = early_reset_static_par0_go_out;
wire _guard18552 = _guard18550 & _guard18551;
wire _guard18553 = early_reset_static_par0_go_out;
wire _guard18554 = early_reset_static_par0_go_out;
wire _guard18555 = early_reset_static_par0_go_out;
wire _guard18556 = early_reset_static_par0_go_out;
wire _guard18557 = early_reset_static_par0_go_out;
wire _guard18558 = early_reset_static_par0_go_out;
wire _guard18559 = ~_guard0;
wire _guard18560 = early_reset_static_par0_go_out;
wire _guard18561 = _guard18559 & _guard18560;
wire _guard18562 = early_reset_static_par0_go_out;
wire _guard18563 = ~_guard0;
wire _guard18564 = early_reset_static_par0_go_out;
wire _guard18565 = _guard18563 & _guard18564;
wire _guard18566 = early_reset_static_par0_go_out;
wire _guard18567 = ~_guard0;
wire _guard18568 = early_reset_static_par0_go_out;
wire _guard18569 = _guard18567 & _guard18568;
wire _guard18570 = early_reset_static_par0_go_out;
wire _guard18571 = early_reset_static_par0_go_out;
wire _guard18572 = early_reset_static_par0_go_out;
wire _guard18573 = ~_guard0;
wire _guard18574 = early_reset_static_par0_go_out;
wire _guard18575 = _guard18573 & _guard18574;
wire _guard18576 = ~_guard0;
wire _guard18577 = early_reset_static_par0_go_out;
wire _guard18578 = _guard18576 & _guard18577;
wire _guard18579 = early_reset_static_par0_go_out;
wire _guard18580 = early_reset_static_par0_go_out;
wire _guard18581 = early_reset_static_par0_go_out;
wire _guard18582 = early_reset_static_par0_go_out;
wire _guard18583 = ~_guard0;
wire _guard18584 = early_reset_static_par0_go_out;
wire _guard18585 = _guard18583 & _guard18584;
wire _guard18586 = early_reset_static_par0_go_out;
wire _guard18587 = early_reset_static_par0_go_out;
wire _guard18588 = ~_guard0;
wire _guard18589 = early_reset_static_par0_go_out;
wire _guard18590 = _guard18588 & _guard18589;
wire _guard18591 = early_reset_static_par0_go_out;
wire _guard18592 = early_reset_static_par0_go_out;
wire _guard18593 = early_reset_static_par0_go_out;
wire _guard18594 = ~_guard0;
wire _guard18595 = early_reset_static_par0_go_out;
wire _guard18596 = _guard18594 & _guard18595;
wire _guard18597 = early_reset_static_par0_go_out;
wire _guard18598 = early_reset_static_par0_go_out;
wire _guard18599 = ~_guard0;
wire _guard18600 = early_reset_static_par0_go_out;
wire _guard18601 = _guard18599 & _guard18600;
wire _guard18602 = early_reset_static_par0_go_out;
wire _guard18603 = early_reset_static_par0_go_out;
wire _guard18604 = ~_guard0;
wire _guard18605 = early_reset_static_par0_go_out;
wire _guard18606 = _guard18604 & _guard18605;
wire _guard18607 = early_reset_static_par0_go_out;
wire _guard18608 = early_reset_static_par0_go_out;
wire _guard18609 = ~_guard0;
wire _guard18610 = early_reset_static_par0_go_out;
wire _guard18611 = _guard18609 & _guard18610;
wire _guard18612 = ~_guard0;
wire _guard18613 = early_reset_static_par0_go_out;
wire _guard18614 = _guard18612 & _guard18613;
wire _guard18615 = early_reset_static_par0_go_out;
wire _guard18616 = early_reset_static_par0_go_out;
wire _guard18617 = early_reset_static_par0_go_out;
wire _guard18618 = early_reset_static_par0_go_out;
wire _guard18619 = early_reset_static_par0_go_out;
wire _guard18620 = early_reset_static_par0_go_out;
wire _guard18621 = early_reset_static_par0_go_out;
wire _guard18622 = ~_guard0;
wire _guard18623 = early_reset_static_par0_go_out;
wire _guard18624 = _guard18622 & _guard18623;
wire _guard18625 = early_reset_static_par0_go_out;
wire _guard18626 = early_reset_static_par0_go_out;
wire _guard18627 = early_reset_static_par0_go_out;
wire _guard18628 = early_reset_static_par0_go_out;
wire _guard18629 = ~_guard0;
wire _guard18630 = early_reset_static_par0_go_out;
wire _guard18631 = _guard18629 & _guard18630;
wire _guard18632 = ~_guard0;
wire _guard18633 = early_reset_static_par0_go_out;
wire _guard18634 = _guard18632 & _guard18633;
wire _guard18635 = early_reset_static_par0_go_out;
wire _guard18636 = early_reset_static_par0_go_out;
wire _guard18637 = early_reset_static_par0_go_out;
wire _guard18638 = early_reset_static_par0_go_out;
wire _guard18639 = early_reset_static_par0_go_out;
wire _guard18640 = early_reset_static_par0_go_out;
wire _guard18641 = early_reset_static_par0_go_out;
wire _guard18642 = early_reset_static_par0_go_out;
wire _guard18643 = early_reset_static_par0_go_out;
wire _guard18644 = early_reset_static_par0_go_out;
wire _guard18645 = ~_guard0;
wire _guard18646 = early_reset_static_par0_go_out;
wire _guard18647 = _guard18645 & _guard18646;
wire _guard18648 = ~_guard0;
wire _guard18649 = early_reset_static_par0_go_out;
wire _guard18650 = _guard18648 & _guard18649;
wire _guard18651 = early_reset_static_par0_go_out;
wire _guard18652 = early_reset_static_par0_go_out;
wire _guard18653 = ~_guard0;
wire _guard18654 = early_reset_static_par0_go_out;
wire _guard18655 = _guard18653 & _guard18654;
wire _guard18656 = early_reset_static_par0_go_out;
wire _guard18657 = early_reset_static_par0_go_out;
wire _guard18658 = early_reset_static_par0_go_out;
wire _guard18659 = early_reset_static_par0_go_out;
wire _guard18660 = early_reset_static_par0_go_out;
wire _guard18661 = ~_guard0;
wire _guard18662 = early_reset_static_par0_go_out;
wire _guard18663 = _guard18661 & _guard18662;
wire _guard18664 = ~_guard0;
wire _guard18665 = early_reset_static_par0_go_out;
wire _guard18666 = _guard18664 & _guard18665;
wire _guard18667 = early_reset_static_par0_go_out;
wire _guard18668 = early_reset_static_par0_go_out;
wire _guard18669 = early_reset_static_par0_go_out;
wire _guard18670 = early_reset_static_par0_go_out;
wire _guard18671 = early_reset_static_par0_go_out;
wire _guard18672 = early_reset_static_par0_go_out;
wire _guard18673 = early_reset_static_par0_go_out;
wire _guard18674 = ~_guard0;
wire _guard18675 = early_reset_static_par0_go_out;
wire _guard18676 = _guard18674 & _guard18675;
wire _guard18677 = early_reset_static_par0_go_out;
wire _guard18678 = early_reset_static_par0_go_out;
wire _guard18679 = early_reset_static_par0_go_out;
wire _guard18680 = ~_guard0;
wire _guard18681 = early_reset_static_par0_go_out;
wire _guard18682 = _guard18680 & _guard18681;
wire _guard18683 = early_reset_static_par0_go_out;
wire _guard18684 = early_reset_static_par0_go_out;
wire _guard18685 = early_reset_static_par0_go_out;
wire _guard18686 = early_reset_static_par0_go_out;
wire _guard18687 = early_reset_static_par0_go_out;
wire _guard18688 = early_reset_static_par0_go_out;
wire _guard18689 = early_reset_static_par0_go_out;
wire _guard18690 = early_reset_static_par0_go_out;
wire _guard18691 = early_reset_static_par0_go_out;
wire _guard18692 = early_reset_static_par0_go_out;
wire _guard18693 = ~_guard0;
wire _guard18694 = early_reset_static_par0_go_out;
wire _guard18695 = _guard18693 & _guard18694;
wire _guard18696 = early_reset_static_par0_go_out;
wire _guard18697 = early_reset_static_par0_go_out;
wire _guard18698 = early_reset_static_par0_go_out;
wire _guard18699 = early_reset_static_par0_go_out;
wire _guard18700 = early_reset_static_par0_go_out;
wire _guard18701 = early_reset_static_par0_go_out;
wire _guard18702 = early_reset_static_par0_go_out;
wire _guard18703 = early_reset_static_par0_go_out;
wire _guard18704 = early_reset_static_par0_go_out;
wire _guard18705 = early_reset_static_par0_go_out;
wire _guard18706 = ~_guard0;
wire _guard18707 = early_reset_static_par0_go_out;
wire _guard18708 = _guard18706 & _guard18707;
wire _guard18709 = early_reset_static_par0_go_out;
wire _guard18710 = early_reset_static_par0_go_out;
wire _guard18711 = early_reset_static_par0_go_out;
wire _guard18712 = ~_guard0;
wire _guard18713 = early_reset_static_par0_go_out;
wire _guard18714 = _guard18712 & _guard18713;
wire _guard18715 = early_reset_static_par0_go_out;
wire _guard18716 = early_reset_static_par0_go_out;
wire _guard18717 = early_reset_static_par0_go_out;
wire _guard18718 = early_reset_static_par0_go_out;
wire _guard18719 = early_reset_static_par0_go_out;
wire _guard18720 = early_reset_static_par0_go_out;
wire _guard18721 = early_reset_static_par0_go_out;
wire _guard18722 = early_reset_static_par0_go_out;
wire _guard18723 = ~_guard0;
wire _guard18724 = early_reset_static_par0_go_out;
wire _guard18725 = _guard18723 & _guard18724;
wire _guard18726 = early_reset_static_par0_go_out;
wire _guard18727 = early_reset_static_par0_go_out;
wire _guard18728 = early_reset_static_par0_go_out;
wire _guard18729 = early_reset_static_par0_go_out;
wire _guard18730 = ~_guard0;
wire _guard18731 = early_reset_static_par0_go_out;
wire _guard18732 = _guard18730 & _guard18731;
wire _guard18733 = early_reset_static_par0_go_out;
wire _guard18734 = early_reset_static_par0_go_out;
wire _guard18735 = early_reset_static_par0_go_out;
wire _guard18736 = early_reset_static_par0_go_out;
wire _guard18737 = early_reset_static_par0_go_out;
wire _guard18738 = early_reset_static_par0_go_out;
wire _guard18739 = early_reset_static_par0_go_out;
wire _guard18740 = ~_guard0;
wire _guard18741 = early_reset_static_par0_go_out;
wire _guard18742 = _guard18740 & _guard18741;
wire _guard18743 = early_reset_static_par0_go_out;
wire _guard18744 = ~_guard0;
wire _guard18745 = early_reset_static_par0_go_out;
wire _guard18746 = _guard18744 & _guard18745;
wire _guard18747 = early_reset_static_par0_go_out;
wire _guard18748 = early_reset_static_par0_go_out;
wire _guard18749 = ~_guard0;
wire _guard18750 = early_reset_static_par0_go_out;
wire _guard18751 = _guard18749 & _guard18750;
wire _guard18752 = ~_guard0;
wire _guard18753 = early_reset_static_par0_go_out;
wire _guard18754 = _guard18752 & _guard18753;
wire _guard18755 = early_reset_static_par0_go_out;
wire _guard18756 = ~_guard0;
wire _guard18757 = early_reset_static_par0_go_out;
wire _guard18758 = _guard18756 & _guard18757;
wire _guard18759 = early_reset_static_par0_go_out;
wire _guard18760 = ~_guard0;
wire _guard18761 = early_reset_static_par0_go_out;
wire _guard18762 = _guard18760 & _guard18761;
wire _guard18763 = early_reset_static_par0_go_out;
wire _guard18764 = early_reset_static_par0_go_out;
wire _guard18765 = ~_guard0;
wire _guard18766 = early_reset_static_par0_go_out;
wire _guard18767 = _guard18765 & _guard18766;
wire _guard18768 = ~_guard0;
wire _guard18769 = early_reset_static_par0_go_out;
wire _guard18770 = _guard18768 & _guard18769;
wire _guard18771 = early_reset_static_par0_go_out;
wire _guard18772 = early_reset_static_par0_go_out;
wire _guard18773 = early_reset_static_par0_go_out;
wire _guard18774 = ~_guard0;
wire _guard18775 = early_reset_static_par0_go_out;
wire _guard18776 = _guard18774 & _guard18775;
wire _guard18777 = early_reset_static_par0_go_out;
wire _guard18778 = early_reset_static_par0_go_out;
wire _guard18779 = early_reset_static_par0_go_out;
wire _guard18780 = ~_guard0;
wire _guard18781 = early_reset_static_par0_go_out;
wire _guard18782 = _guard18780 & _guard18781;
wire _guard18783 = early_reset_static_par0_go_out;
wire _guard18784 = early_reset_static_par0_go_out;
wire _guard18785 = ~_guard0;
wire _guard18786 = early_reset_static_par0_go_out;
wire _guard18787 = _guard18785 & _guard18786;
wire _guard18788 = ~_guard0;
wire _guard18789 = early_reset_static_par0_go_out;
wire _guard18790 = _guard18788 & _guard18789;
wire _guard18791 = early_reset_static_par0_go_out;
wire _guard18792 = early_reset_static_par0_go_out;
wire _guard18793 = ~_guard0;
wire _guard18794 = early_reset_static_par0_go_out;
wire _guard18795 = _guard18793 & _guard18794;
wire _guard18796 = early_reset_static_par0_go_out;
wire _guard18797 = early_reset_static_par0_go_out;
wire _guard18798 = early_reset_static_par0_go_out;
wire _guard18799 = early_reset_static_par0_go_out;
wire _guard18800 = early_reset_static_par0_go_out;
wire _guard18801 = early_reset_static_par0_go_out;
wire _guard18802 = early_reset_static_par0_go_out;
wire _guard18803 = ~_guard0;
wire _guard18804 = early_reset_static_par0_go_out;
wire _guard18805 = _guard18803 & _guard18804;
wire _guard18806 = early_reset_static_par0_go_out;
wire _guard18807 = early_reset_static_par0_go_out;
wire _guard18808 = early_reset_static_par0_go_out;
wire _guard18809 = ~_guard0;
wire _guard18810 = early_reset_static_par0_go_out;
wire _guard18811 = _guard18809 & _guard18810;
wire _guard18812 = early_reset_static_par0_go_out;
wire _guard18813 = early_reset_static_par0_go_out;
wire _guard18814 = early_reset_static_par0_go_out;
wire _guard18815 = ~_guard0;
wire _guard18816 = early_reset_static_par0_go_out;
wire _guard18817 = _guard18815 & _guard18816;
wire _guard18818 = ~_guard0;
wire _guard18819 = early_reset_static_par0_go_out;
wire _guard18820 = _guard18818 & _guard18819;
wire _guard18821 = early_reset_static_par0_go_out;
wire _guard18822 = early_reset_static_par0_go_out;
wire _guard18823 = ~_guard0;
wire _guard18824 = early_reset_static_par0_go_out;
wire _guard18825 = _guard18823 & _guard18824;
wire _guard18826 = early_reset_static_par0_go_out;
wire _guard18827 = early_reset_static_par0_go_out;
wire _guard18828 = early_reset_static_par0_go_out;
wire _guard18829 = early_reset_static_par0_go_out;
wire _guard18830 = early_reset_static_par0_go_out;
wire _guard18831 = early_reset_static_par0_go_out;
wire _guard18832 = early_reset_static_par0_go_out;
wire _guard18833 = early_reset_static_par0_go_out;
wire _guard18834 = ~_guard0;
wire _guard18835 = early_reset_static_par0_go_out;
wire _guard18836 = _guard18834 & _guard18835;
wire _guard18837 = early_reset_static_par0_go_out;
wire _guard18838 = ~_guard0;
wire _guard18839 = early_reset_static_par0_go_out;
wire _guard18840 = _guard18838 & _guard18839;
wire _guard18841 = early_reset_static_par0_go_out;
wire _guard18842 = early_reset_static_par0_go_out;
wire _guard18843 = ~_guard0;
wire _guard18844 = early_reset_static_par0_go_out;
wire _guard18845 = _guard18843 & _guard18844;
wire _guard18846 = early_reset_static_par0_go_out;
wire _guard18847 = early_reset_static_par0_go_out;
wire _guard18848 = ~_guard0;
wire _guard18849 = early_reset_static_par0_go_out;
wire _guard18850 = _guard18848 & _guard18849;
wire _guard18851 = early_reset_static_par0_go_out;
wire _guard18852 = early_reset_static_par0_go_out;
wire _guard18853 = ~_guard0;
wire _guard18854 = early_reset_static_par0_go_out;
wire _guard18855 = _guard18853 & _guard18854;
wire _guard18856 = early_reset_static_par0_go_out;
wire _guard18857 = ~_guard0;
wire _guard18858 = early_reset_static_par0_go_out;
wire _guard18859 = _guard18857 & _guard18858;
wire _guard18860 = early_reset_static_par0_go_out;
wire _guard18861 = early_reset_static_par0_go_out;
wire _guard18862 = ~_guard0;
wire _guard18863 = early_reset_static_par0_go_out;
wire _guard18864 = _guard18862 & _guard18863;
wire _guard18865 = early_reset_static_par0_go_out;
wire _guard18866 = ~_guard0;
wire _guard18867 = early_reset_static_par0_go_out;
wire _guard18868 = _guard18866 & _guard18867;
wire _guard18869 = early_reset_static_par0_go_out;
wire _guard18870 = early_reset_static_par0_go_out;
wire _guard18871 = ~_guard0;
wire _guard18872 = early_reset_static_par0_go_out;
wire _guard18873 = _guard18871 & _guard18872;
wire _guard18874 = ~_guard0;
wire _guard18875 = early_reset_static_par0_go_out;
wire _guard18876 = _guard18874 & _guard18875;
wire _guard18877 = early_reset_static_par0_go_out;
wire _guard18878 = early_reset_static_par0_go_out;
wire _guard18879 = ~_guard0;
wire _guard18880 = early_reset_static_par0_go_out;
wire _guard18881 = _guard18879 & _guard18880;
wire _guard18882 = ~_guard0;
wire _guard18883 = early_reset_static_par0_go_out;
wire _guard18884 = _guard18882 & _guard18883;
wire _guard18885 = early_reset_static_par0_go_out;
wire _guard18886 = ~_guard0;
wire _guard18887 = early_reset_static_par0_go_out;
wire _guard18888 = _guard18886 & _guard18887;
wire _guard18889 = early_reset_static_par0_go_out;
wire _guard18890 = early_reset_static_par0_go_out;
wire _guard18891 = early_reset_static_par0_go_out;
wire _guard18892 = early_reset_static_par0_go_out;
wire _guard18893 = early_reset_static_par0_go_out;
wire _guard18894 = ~_guard0;
wire _guard18895 = early_reset_static_par0_go_out;
wire _guard18896 = _guard18894 & _guard18895;
wire _guard18897 = early_reset_static_par0_go_out;
wire _guard18898 = early_reset_static_par0_go_out;
wire _guard18899 = ~_guard0;
wire _guard18900 = early_reset_static_par0_go_out;
wire _guard18901 = _guard18899 & _guard18900;
wire _guard18902 = early_reset_static_par0_go_out;
wire _guard18903 = early_reset_static_par0_go_out;
wire _guard18904 = fsm0_out == 6'd0;
wire _guard18905 = signal_reg_out;
wire _guard18906 = _guard18904 & _guard18905;
wire _guard18907 = fsm0_out == 6'd0;
wire _guard18908 = signal_reg_out;
wire _guard18909 = ~_guard18908;
wire _guard18910 = _guard18907 & _guard18909;
wire _guard18911 = wrapper_early_reset_static_seq_go_out;
wire _guard18912 = _guard18910 & _guard18911;
wire _guard18913 = _guard18906 | _guard18912;
wire _guard18914 = fsm0_out == 6'd0;
wire _guard18915 = signal_reg_out;
wire _guard18916 = ~_guard18915;
wire _guard18917 = _guard18914 & _guard18916;
wire _guard18918 = wrapper_early_reset_static_seq_go_out;
wire _guard18919 = _guard18917 & _guard18918;
wire _guard18920 = fsm0_out == 6'd0;
wire _guard18921 = signal_reg_out;
wire _guard18922 = _guard18920 & _guard18921;
wire _guard18923 = cond_wire19_out;
wire _guard18924 = early_reset_static_par0_go_out;
wire _guard18925 = _guard18923 & _guard18924;
wire _guard18926 = cond_wire19_out;
wire _guard18927 = early_reset_static_par0_go_out;
wire _guard18928 = _guard18926 & _guard18927;
wire _guard18929 = cond_wire21_out;
wire _guard18930 = early_reset_static_par0_go_out;
wire _guard18931 = _guard18929 & _guard18930;
wire _guard18932 = cond_wire21_out;
wire _guard18933 = early_reset_static_par0_go_out;
wire _guard18934 = _guard18932 & _guard18933;
wire _guard18935 = cond_wire49_out;
wire _guard18936 = early_reset_static_par0_go_out;
wire _guard18937 = _guard18935 & _guard18936;
wire _guard18938 = cond_wire49_out;
wire _guard18939 = early_reset_static_par0_go_out;
wire _guard18940 = _guard18938 & _guard18939;
wire _guard18941 = cond_wire126_out;
wire _guard18942 = early_reset_static_par0_go_out;
wire _guard18943 = _guard18941 & _guard18942;
wire _guard18944 = cond_wire124_out;
wire _guard18945 = early_reset_static_par0_go_out;
wire _guard18946 = _guard18944 & _guard18945;
wire _guard18947 = fsm_out == 1'd0;
wire _guard18948 = cond_wire124_out;
wire _guard18949 = _guard18947 & _guard18948;
wire _guard18950 = fsm_out == 1'd0;
wire _guard18951 = _guard18949 & _guard18950;
wire _guard18952 = fsm_out == 1'd0;
wire _guard18953 = cond_wire126_out;
wire _guard18954 = _guard18952 & _guard18953;
wire _guard18955 = fsm_out == 1'd0;
wire _guard18956 = _guard18954 & _guard18955;
wire _guard18957 = _guard18951 | _guard18956;
wire _guard18958 = early_reset_static_par0_go_out;
wire _guard18959 = _guard18957 & _guard18958;
wire _guard18960 = fsm_out == 1'd0;
wire _guard18961 = cond_wire124_out;
wire _guard18962 = _guard18960 & _guard18961;
wire _guard18963 = fsm_out == 1'd0;
wire _guard18964 = _guard18962 & _guard18963;
wire _guard18965 = fsm_out == 1'd0;
wire _guard18966 = cond_wire126_out;
wire _guard18967 = _guard18965 & _guard18966;
wire _guard18968 = fsm_out == 1'd0;
wire _guard18969 = _guard18967 & _guard18968;
wire _guard18970 = _guard18964 | _guard18969;
wire _guard18971 = early_reset_static_par0_go_out;
wire _guard18972 = _guard18970 & _guard18971;
wire _guard18973 = fsm_out == 1'd0;
wire _guard18974 = cond_wire124_out;
wire _guard18975 = _guard18973 & _guard18974;
wire _guard18976 = fsm_out == 1'd0;
wire _guard18977 = _guard18975 & _guard18976;
wire _guard18978 = fsm_out == 1'd0;
wire _guard18979 = cond_wire126_out;
wire _guard18980 = _guard18978 & _guard18979;
wire _guard18981 = fsm_out == 1'd0;
wire _guard18982 = _guard18980 & _guard18981;
wire _guard18983 = _guard18977 | _guard18982;
wire _guard18984 = early_reset_static_par0_go_out;
wire _guard18985 = _guard18983 & _guard18984;
wire _guard18986 = cond_wire125_out;
wire _guard18987 = early_reset_static_par0_go_out;
wire _guard18988 = _guard18986 & _guard18987;
wire _guard18989 = cond_wire125_out;
wire _guard18990 = early_reset_static_par0_go_out;
wire _guard18991 = _guard18989 & _guard18990;
wire _guard18992 = cond_wire147_out;
wire _guard18993 = early_reset_static_par0_go_out;
wire _guard18994 = _guard18992 & _guard18993;
wire _guard18995 = cond_wire145_out;
wire _guard18996 = early_reset_static_par0_go_out;
wire _guard18997 = _guard18995 & _guard18996;
wire _guard18998 = fsm_out == 1'd0;
wire _guard18999 = cond_wire145_out;
wire _guard19000 = _guard18998 & _guard18999;
wire _guard19001 = fsm_out == 1'd0;
wire _guard19002 = _guard19000 & _guard19001;
wire _guard19003 = fsm_out == 1'd0;
wire _guard19004 = cond_wire147_out;
wire _guard19005 = _guard19003 & _guard19004;
wire _guard19006 = fsm_out == 1'd0;
wire _guard19007 = _guard19005 & _guard19006;
wire _guard19008 = _guard19002 | _guard19007;
wire _guard19009 = early_reset_static_par0_go_out;
wire _guard19010 = _guard19008 & _guard19009;
wire _guard19011 = fsm_out == 1'd0;
wire _guard19012 = cond_wire145_out;
wire _guard19013 = _guard19011 & _guard19012;
wire _guard19014 = fsm_out == 1'd0;
wire _guard19015 = _guard19013 & _guard19014;
wire _guard19016 = fsm_out == 1'd0;
wire _guard19017 = cond_wire147_out;
wire _guard19018 = _guard19016 & _guard19017;
wire _guard19019 = fsm_out == 1'd0;
wire _guard19020 = _guard19018 & _guard19019;
wire _guard19021 = _guard19015 | _guard19020;
wire _guard19022 = early_reset_static_par0_go_out;
wire _guard19023 = _guard19021 & _guard19022;
wire _guard19024 = fsm_out == 1'd0;
wire _guard19025 = cond_wire145_out;
wire _guard19026 = _guard19024 & _guard19025;
wire _guard19027 = fsm_out == 1'd0;
wire _guard19028 = _guard19026 & _guard19027;
wire _guard19029 = fsm_out == 1'd0;
wire _guard19030 = cond_wire147_out;
wire _guard19031 = _guard19029 & _guard19030;
wire _guard19032 = fsm_out == 1'd0;
wire _guard19033 = _guard19031 & _guard19032;
wire _guard19034 = _guard19028 | _guard19033;
wire _guard19035 = early_reset_static_par0_go_out;
wire _guard19036 = _guard19034 & _guard19035;
wire _guard19037 = cond_wire146_out;
wire _guard19038 = early_reset_static_par0_go_out;
wire _guard19039 = _guard19037 & _guard19038;
wire _guard19040 = cond_wire146_out;
wire _guard19041 = early_reset_static_par0_go_out;
wire _guard19042 = _guard19040 & _guard19041;
wire _guard19043 = cond_wire89_out;
wire _guard19044 = early_reset_static_par0_go_out;
wire _guard19045 = _guard19043 & _guard19044;
wire _guard19046 = cond_wire89_out;
wire _guard19047 = early_reset_static_par0_go_out;
wire _guard19048 = _guard19046 & _guard19047;
wire _guard19049 = cond_wire162_out;
wire _guard19050 = early_reset_static_par0_go_out;
wire _guard19051 = _guard19049 & _guard19050;
wire _guard19052 = cond_wire162_out;
wire _guard19053 = early_reset_static_par0_go_out;
wire _guard19054 = _guard19052 & _guard19053;
wire _guard19055 = cond_wire231_out;
wire _guard19056 = early_reset_static_par0_go_out;
wire _guard19057 = _guard19055 & _guard19056;
wire _guard19058 = cond_wire231_out;
wire _guard19059 = early_reset_static_par0_go_out;
wire _guard19060 = _guard19058 & _guard19059;
wire _guard19061 = cond_wire239_out;
wire _guard19062 = early_reset_static_par0_go_out;
wire _guard19063 = _guard19061 & _guard19062;
wire _guard19064 = cond_wire239_out;
wire _guard19065 = early_reset_static_par0_go_out;
wire _guard19066 = _guard19064 & _guard19065;
wire _guard19067 = cond_wire260_out;
wire _guard19068 = early_reset_static_par0_go_out;
wire _guard19069 = _guard19067 & _guard19068;
wire _guard19070 = cond_wire258_out;
wire _guard19071 = early_reset_static_par0_go_out;
wire _guard19072 = _guard19070 & _guard19071;
wire _guard19073 = fsm_out == 1'd0;
wire _guard19074 = cond_wire258_out;
wire _guard19075 = _guard19073 & _guard19074;
wire _guard19076 = fsm_out == 1'd0;
wire _guard19077 = _guard19075 & _guard19076;
wire _guard19078 = fsm_out == 1'd0;
wire _guard19079 = cond_wire260_out;
wire _guard19080 = _guard19078 & _guard19079;
wire _guard19081 = fsm_out == 1'd0;
wire _guard19082 = _guard19080 & _guard19081;
wire _guard19083 = _guard19077 | _guard19082;
wire _guard19084 = early_reset_static_par0_go_out;
wire _guard19085 = _guard19083 & _guard19084;
wire _guard19086 = fsm_out == 1'd0;
wire _guard19087 = cond_wire258_out;
wire _guard19088 = _guard19086 & _guard19087;
wire _guard19089 = fsm_out == 1'd0;
wire _guard19090 = _guard19088 & _guard19089;
wire _guard19091 = fsm_out == 1'd0;
wire _guard19092 = cond_wire260_out;
wire _guard19093 = _guard19091 & _guard19092;
wire _guard19094 = fsm_out == 1'd0;
wire _guard19095 = _guard19093 & _guard19094;
wire _guard19096 = _guard19090 | _guard19095;
wire _guard19097 = early_reset_static_par0_go_out;
wire _guard19098 = _guard19096 & _guard19097;
wire _guard19099 = fsm_out == 1'd0;
wire _guard19100 = cond_wire258_out;
wire _guard19101 = _guard19099 & _guard19100;
wire _guard19102 = fsm_out == 1'd0;
wire _guard19103 = _guard19101 & _guard19102;
wire _guard19104 = fsm_out == 1'd0;
wire _guard19105 = cond_wire260_out;
wire _guard19106 = _guard19104 & _guard19105;
wire _guard19107 = fsm_out == 1'd0;
wire _guard19108 = _guard19106 & _guard19107;
wire _guard19109 = _guard19103 | _guard19108;
wire _guard19110 = early_reset_static_par0_go_out;
wire _guard19111 = _guard19109 & _guard19110;
wire _guard19112 = cond_wire194_out;
wire _guard19113 = early_reset_static_par0_go_out;
wire _guard19114 = _guard19112 & _guard19113;
wire _guard19115 = cond_wire194_out;
wire _guard19116 = early_reset_static_par0_go_out;
wire _guard19117 = _guard19115 & _guard19116;
wire _guard19118 = cond_wire267_out;
wire _guard19119 = early_reset_static_par0_go_out;
wire _guard19120 = _guard19118 & _guard19119;
wire _guard19121 = cond_wire267_out;
wire _guard19122 = early_reset_static_par0_go_out;
wire _guard19123 = _guard19121 & _guard19122;
wire _guard19124 = cond_wire293_out;
wire _guard19125 = early_reset_static_par0_go_out;
wire _guard19126 = _guard19124 & _guard19125;
wire _guard19127 = cond_wire291_out;
wire _guard19128 = early_reset_static_par0_go_out;
wire _guard19129 = _guard19127 & _guard19128;
wire _guard19130 = fsm_out == 1'd0;
wire _guard19131 = cond_wire291_out;
wire _guard19132 = _guard19130 & _guard19131;
wire _guard19133 = fsm_out == 1'd0;
wire _guard19134 = _guard19132 & _guard19133;
wire _guard19135 = fsm_out == 1'd0;
wire _guard19136 = cond_wire293_out;
wire _guard19137 = _guard19135 & _guard19136;
wire _guard19138 = fsm_out == 1'd0;
wire _guard19139 = _guard19137 & _guard19138;
wire _guard19140 = _guard19134 | _guard19139;
wire _guard19141 = early_reset_static_par0_go_out;
wire _guard19142 = _guard19140 & _guard19141;
wire _guard19143 = fsm_out == 1'd0;
wire _guard19144 = cond_wire291_out;
wire _guard19145 = _guard19143 & _guard19144;
wire _guard19146 = fsm_out == 1'd0;
wire _guard19147 = _guard19145 & _guard19146;
wire _guard19148 = fsm_out == 1'd0;
wire _guard19149 = cond_wire293_out;
wire _guard19150 = _guard19148 & _guard19149;
wire _guard19151 = fsm_out == 1'd0;
wire _guard19152 = _guard19150 & _guard19151;
wire _guard19153 = _guard19147 | _guard19152;
wire _guard19154 = early_reset_static_par0_go_out;
wire _guard19155 = _guard19153 & _guard19154;
wire _guard19156 = fsm_out == 1'd0;
wire _guard19157 = cond_wire291_out;
wire _guard19158 = _guard19156 & _guard19157;
wire _guard19159 = fsm_out == 1'd0;
wire _guard19160 = _guard19158 & _guard19159;
wire _guard19161 = fsm_out == 1'd0;
wire _guard19162 = cond_wire293_out;
wire _guard19163 = _guard19161 & _guard19162;
wire _guard19164 = fsm_out == 1'd0;
wire _guard19165 = _guard19163 & _guard19164;
wire _guard19166 = _guard19160 | _guard19165;
wire _guard19167 = early_reset_static_par0_go_out;
wire _guard19168 = _guard19166 & _guard19167;
wire _guard19169 = cond_wire288_out;
wire _guard19170 = early_reset_static_par0_go_out;
wire _guard19171 = _guard19169 & _guard19170;
wire _guard19172 = cond_wire288_out;
wire _guard19173 = early_reset_static_par0_go_out;
wire _guard19174 = _guard19172 & _guard19173;
wire _guard19175 = cond_wire305_out;
wire _guard19176 = early_reset_static_par0_go_out;
wire _guard19177 = _guard19175 & _guard19176;
wire _guard19178 = cond_wire303_out;
wire _guard19179 = early_reset_static_par0_go_out;
wire _guard19180 = _guard19178 & _guard19179;
wire _guard19181 = fsm_out == 1'd0;
wire _guard19182 = cond_wire303_out;
wire _guard19183 = _guard19181 & _guard19182;
wire _guard19184 = fsm_out == 1'd0;
wire _guard19185 = _guard19183 & _guard19184;
wire _guard19186 = fsm_out == 1'd0;
wire _guard19187 = cond_wire305_out;
wire _guard19188 = _guard19186 & _guard19187;
wire _guard19189 = fsm_out == 1'd0;
wire _guard19190 = _guard19188 & _guard19189;
wire _guard19191 = _guard19185 | _guard19190;
wire _guard19192 = early_reset_static_par0_go_out;
wire _guard19193 = _guard19191 & _guard19192;
wire _guard19194 = fsm_out == 1'd0;
wire _guard19195 = cond_wire303_out;
wire _guard19196 = _guard19194 & _guard19195;
wire _guard19197 = fsm_out == 1'd0;
wire _guard19198 = _guard19196 & _guard19197;
wire _guard19199 = fsm_out == 1'd0;
wire _guard19200 = cond_wire305_out;
wire _guard19201 = _guard19199 & _guard19200;
wire _guard19202 = fsm_out == 1'd0;
wire _guard19203 = _guard19201 & _guard19202;
wire _guard19204 = _guard19198 | _guard19203;
wire _guard19205 = early_reset_static_par0_go_out;
wire _guard19206 = _guard19204 & _guard19205;
wire _guard19207 = fsm_out == 1'd0;
wire _guard19208 = cond_wire303_out;
wire _guard19209 = _guard19207 & _guard19208;
wire _guard19210 = fsm_out == 1'd0;
wire _guard19211 = _guard19209 & _guard19210;
wire _guard19212 = fsm_out == 1'd0;
wire _guard19213 = cond_wire305_out;
wire _guard19214 = _guard19212 & _guard19213;
wire _guard19215 = fsm_out == 1'd0;
wire _guard19216 = _guard19214 & _guard19215;
wire _guard19217 = _guard19211 | _guard19216;
wire _guard19218 = early_reset_static_par0_go_out;
wire _guard19219 = _guard19217 & _guard19218;
wire _guard19220 = cond_wire255_out;
wire _guard19221 = early_reset_static_par0_go_out;
wire _guard19222 = _guard19220 & _guard19221;
wire _guard19223 = cond_wire255_out;
wire _guard19224 = early_reset_static_par0_go_out;
wire _guard19225 = _guard19223 & _guard19224;
wire _guard19226 = cond_wire259_out;
wire _guard19227 = early_reset_static_par0_go_out;
wire _guard19228 = _guard19226 & _guard19227;
wire _guard19229 = cond_wire259_out;
wire _guard19230 = early_reset_static_par0_go_out;
wire _guard19231 = _guard19229 & _guard19230;
wire _guard19232 = cond_wire329_out;
wire _guard19233 = early_reset_static_par0_go_out;
wire _guard19234 = _guard19232 & _guard19233;
wire _guard19235 = cond_wire327_out;
wire _guard19236 = early_reset_static_par0_go_out;
wire _guard19237 = _guard19235 & _guard19236;
wire _guard19238 = fsm_out == 1'd0;
wire _guard19239 = cond_wire327_out;
wire _guard19240 = _guard19238 & _guard19239;
wire _guard19241 = fsm_out == 1'd0;
wire _guard19242 = _guard19240 & _guard19241;
wire _guard19243 = fsm_out == 1'd0;
wire _guard19244 = cond_wire329_out;
wire _guard19245 = _guard19243 & _guard19244;
wire _guard19246 = fsm_out == 1'd0;
wire _guard19247 = _guard19245 & _guard19246;
wire _guard19248 = _guard19242 | _guard19247;
wire _guard19249 = early_reset_static_par0_go_out;
wire _guard19250 = _guard19248 & _guard19249;
wire _guard19251 = fsm_out == 1'd0;
wire _guard19252 = cond_wire327_out;
wire _guard19253 = _guard19251 & _guard19252;
wire _guard19254 = fsm_out == 1'd0;
wire _guard19255 = _guard19253 & _guard19254;
wire _guard19256 = fsm_out == 1'd0;
wire _guard19257 = cond_wire329_out;
wire _guard19258 = _guard19256 & _guard19257;
wire _guard19259 = fsm_out == 1'd0;
wire _guard19260 = _guard19258 & _guard19259;
wire _guard19261 = _guard19255 | _guard19260;
wire _guard19262 = early_reset_static_par0_go_out;
wire _guard19263 = _guard19261 & _guard19262;
wire _guard19264 = fsm_out == 1'd0;
wire _guard19265 = cond_wire327_out;
wire _guard19266 = _guard19264 & _guard19265;
wire _guard19267 = fsm_out == 1'd0;
wire _guard19268 = _guard19266 & _guard19267;
wire _guard19269 = fsm_out == 1'd0;
wire _guard19270 = cond_wire329_out;
wire _guard19271 = _guard19269 & _guard19270;
wire _guard19272 = fsm_out == 1'd0;
wire _guard19273 = _guard19271 & _guard19272;
wire _guard19274 = _guard19268 | _guard19273;
wire _guard19275 = early_reset_static_par0_go_out;
wire _guard19276 = _guard19274 & _guard19275;
wire _guard19277 = cond_wire357_out;
wire _guard19278 = early_reset_static_par0_go_out;
wire _guard19279 = _guard19277 & _guard19278;
wire _guard19280 = cond_wire357_out;
wire _guard19281 = early_reset_static_par0_go_out;
wire _guard19282 = _guard19280 & _guard19281;
wire _guard19283 = cond_wire373_out;
wire _guard19284 = early_reset_static_par0_go_out;
wire _guard19285 = _guard19283 & _guard19284;
wire _guard19286 = cond_wire373_out;
wire _guard19287 = early_reset_static_par0_go_out;
wire _guard19288 = _guard19286 & _guard19287;
wire _guard19289 = cond_wire316_out;
wire _guard19290 = early_reset_static_par0_go_out;
wire _guard19291 = _guard19289 & _guard19290;
wire _guard19292 = cond_wire316_out;
wire _guard19293 = early_reset_static_par0_go_out;
wire _guard19294 = _guard19292 & _guard19293;
wire _guard19295 = cond_wire398_out;
wire _guard19296 = early_reset_static_par0_go_out;
wire _guard19297 = _guard19295 & _guard19296;
wire _guard19298 = cond_wire396_out;
wire _guard19299 = early_reset_static_par0_go_out;
wire _guard19300 = _guard19298 & _guard19299;
wire _guard19301 = fsm_out == 1'd0;
wire _guard19302 = cond_wire396_out;
wire _guard19303 = _guard19301 & _guard19302;
wire _guard19304 = fsm_out == 1'd0;
wire _guard19305 = _guard19303 & _guard19304;
wire _guard19306 = fsm_out == 1'd0;
wire _guard19307 = cond_wire398_out;
wire _guard19308 = _guard19306 & _guard19307;
wire _guard19309 = fsm_out == 1'd0;
wire _guard19310 = _guard19308 & _guard19309;
wire _guard19311 = _guard19305 | _guard19310;
wire _guard19312 = early_reset_static_par0_go_out;
wire _guard19313 = _guard19311 & _guard19312;
wire _guard19314 = fsm_out == 1'd0;
wire _guard19315 = cond_wire396_out;
wire _guard19316 = _guard19314 & _guard19315;
wire _guard19317 = fsm_out == 1'd0;
wire _guard19318 = _guard19316 & _guard19317;
wire _guard19319 = fsm_out == 1'd0;
wire _guard19320 = cond_wire398_out;
wire _guard19321 = _guard19319 & _guard19320;
wire _guard19322 = fsm_out == 1'd0;
wire _guard19323 = _guard19321 & _guard19322;
wire _guard19324 = _guard19318 | _guard19323;
wire _guard19325 = early_reset_static_par0_go_out;
wire _guard19326 = _guard19324 & _guard19325;
wire _guard19327 = fsm_out == 1'd0;
wire _guard19328 = cond_wire396_out;
wire _guard19329 = _guard19327 & _guard19328;
wire _guard19330 = fsm_out == 1'd0;
wire _guard19331 = _guard19329 & _guard19330;
wire _guard19332 = fsm_out == 1'd0;
wire _guard19333 = cond_wire398_out;
wire _guard19334 = _guard19332 & _guard19333;
wire _guard19335 = fsm_out == 1'd0;
wire _guard19336 = _guard19334 & _guard19335;
wire _guard19337 = _guard19331 | _guard19336;
wire _guard19338 = early_reset_static_par0_go_out;
wire _guard19339 = _guard19337 & _guard19338;
wire _guard19340 = cond_wire397_out;
wire _guard19341 = early_reset_static_par0_go_out;
wire _guard19342 = _guard19340 & _guard19341;
wire _guard19343 = cond_wire397_out;
wire _guard19344 = early_reset_static_par0_go_out;
wire _guard19345 = _guard19343 & _guard19344;
wire _guard19346 = cond_wire442_out;
wire _guard19347 = early_reset_static_par0_go_out;
wire _guard19348 = _guard19346 & _guard19347;
wire _guard19349 = cond_wire442_out;
wire _guard19350 = early_reset_static_par0_go_out;
wire _guard19351 = _guard19349 & _guard19350;
wire _guard19352 = cond_wire469_out;
wire _guard19353 = early_reset_static_par0_go_out;
wire _guard19354 = _guard19352 & _guard19353;
wire _guard19355 = cond_wire469_out;
wire _guard19356 = early_reset_static_par0_go_out;
wire _guard19357 = _guard19355 & _guard19356;
wire _guard19358 = cond_wire418_out;
wire _guard19359 = early_reset_static_par0_go_out;
wire _guard19360 = _guard19358 & _guard19359;
wire _guard19361 = cond_wire418_out;
wire _guard19362 = early_reset_static_par0_go_out;
wire _guard19363 = _guard19361 & _guard19362;
wire _guard19364 = cond_wire430_out;
wire _guard19365 = early_reset_static_par0_go_out;
wire _guard19366 = _guard19364 & _guard19365;
wire _guard19367 = cond_wire430_out;
wire _guard19368 = early_reset_static_par0_go_out;
wire _guard19369 = _guard19367 & _guard19368;
wire _guard19370 = cond_wire507_out;
wire _guard19371 = early_reset_static_par0_go_out;
wire _guard19372 = _guard19370 & _guard19371;
wire _guard19373 = cond_wire507_out;
wire _guard19374 = early_reset_static_par0_go_out;
wire _guard19375 = _guard19373 & _guard19374;
wire _guard19376 = cond_wire534_out;
wire _guard19377 = early_reset_static_par0_go_out;
wire _guard19378 = _guard19376 & _guard19377;
wire _guard19379 = cond_wire534_out;
wire _guard19380 = early_reset_static_par0_go_out;
wire _guard19381 = _guard19379 & _guard19380;
wire _guard19382 = cond_wire556_out;
wire _guard19383 = early_reset_static_par0_go_out;
wire _guard19384 = _guard19382 & _guard19383;
wire _guard19385 = cond_wire556_out;
wire _guard19386 = early_reset_static_par0_go_out;
wire _guard19387 = _guard19385 & _guard19386;
wire _guard19388 = cond_wire606_out;
wire _guard19389 = early_reset_static_par0_go_out;
wire _guard19390 = _guard19388 & _guard19389;
wire _guard19391 = cond_wire604_out;
wire _guard19392 = early_reset_static_par0_go_out;
wire _guard19393 = _guard19391 & _guard19392;
wire _guard19394 = fsm_out == 1'd0;
wire _guard19395 = cond_wire604_out;
wire _guard19396 = _guard19394 & _guard19395;
wire _guard19397 = fsm_out == 1'd0;
wire _guard19398 = _guard19396 & _guard19397;
wire _guard19399 = fsm_out == 1'd0;
wire _guard19400 = cond_wire606_out;
wire _guard19401 = _guard19399 & _guard19400;
wire _guard19402 = fsm_out == 1'd0;
wire _guard19403 = _guard19401 & _guard19402;
wire _guard19404 = _guard19398 | _guard19403;
wire _guard19405 = early_reset_static_par0_go_out;
wire _guard19406 = _guard19404 & _guard19405;
wire _guard19407 = fsm_out == 1'd0;
wire _guard19408 = cond_wire604_out;
wire _guard19409 = _guard19407 & _guard19408;
wire _guard19410 = fsm_out == 1'd0;
wire _guard19411 = _guard19409 & _guard19410;
wire _guard19412 = fsm_out == 1'd0;
wire _guard19413 = cond_wire606_out;
wire _guard19414 = _guard19412 & _guard19413;
wire _guard19415 = fsm_out == 1'd0;
wire _guard19416 = _guard19414 & _guard19415;
wire _guard19417 = _guard19411 | _guard19416;
wire _guard19418 = early_reset_static_par0_go_out;
wire _guard19419 = _guard19417 & _guard19418;
wire _guard19420 = fsm_out == 1'd0;
wire _guard19421 = cond_wire604_out;
wire _guard19422 = _guard19420 & _guard19421;
wire _guard19423 = fsm_out == 1'd0;
wire _guard19424 = _guard19422 & _guard19423;
wire _guard19425 = fsm_out == 1'd0;
wire _guard19426 = cond_wire606_out;
wire _guard19427 = _guard19425 & _guard19426;
wire _guard19428 = fsm_out == 1'd0;
wire _guard19429 = _guard19427 & _guard19428;
wire _guard19430 = _guard19424 | _guard19429;
wire _guard19431 = early_reset_static_par0_go_out;
wire _guard19432 = _guard19430 & _guard19431;
wire _guard19433 = cond_wire548_out;
wire _guard19434 = early_reset_static_par0_go_out;
wire _guard19435 = _guard19433 & _guard19434;
wire _guard19436 = cond_wire548_out;
wire _guard19437 = early_reset_static_par0_go_out;
wire _guard19438 = _guard19436 & _guard19437;
wire _guard19439 = cond_wire625_out;
wire _guard19440 = early_reset_static_par0_go_out;
wire _guard19441 = _guard19439 & _guard19440;
wire _guard19442 = cond_wire625_out;
wire _guard19443 = early_reset_static_par0_go_out;
wire _guard19444 = _guard19442 & _guard19443;
wire _guard19445 = cond_wire634_out;
wire _guard19446 = early_reset_static_par0_go_out;
wire _guard19447 = _guard19445 & _guard19446;
wire _guard19448 = cond_wire632_out;
wire _guard19449 = early_reset_static_par0_go_out;
wire _guard19450 = _guard19448 & _guard19449;
wire _guard19451 = fsm_out == 1'd0;
wire _guard19452 = cond_wire632_out;
wire _guard19453 = _guard19451 & _guard19452;
wire _guard19454 = fsm_out == 1'd0;
wire _guard19455 = _guard19453 & _guard19454;
wire _guard19456 = fsm_out == 1'd0;
wire _guard19457 = cond_wire634_out;
wire _guard19458 = _guard19456 & _guard19457;
wire _guard19459 = fsm_out == 1'd0;
wire _guard19460 = _guard19458 & _guard19459;
wire _guard19461 = _guard19455 | _guard19460;
wire _guard19462 = early_reset_static_par0_go_out;
wire _guard19463 = _guard19461 & _guard19462;
wire _guard19464 = fsm_out == 1'd0;
wire _guard19465 = cond_wire632_out;
wire _guard19466 = _guard19464 & _guard19465;
wire _guard19467 = fsm_out == 1'd0;
wire _guard19468 = _guard19466 & _guard19467;
wire _guard19469 = fsm_out == 1'd0;
wire _guard19470 = cond_wire634_out;
wire _guard19471 = _guard19469 & _guard19470;
wire _guard19472 = fsm_out == 1'd0;
wire _guard19473 = _guard19471 & _guard19472;
wire _guard19474 = _guard19468 | _guard19473;
wire _guard19475 = early_reset_static_par0_go_out;
wire _guard19476 = _guard19474 & _guard19475;
wire _guard19477 = fsm_out == 1'd0;
wire _guard19478 = cond_wire632_out;
wire _guard19479 = _guard19477 & _guard19478;
wire _guard19480 = fsm_out == 1'd0;
wire _guard19481 = _guard19479 & _guard19480;
wire _guard19482 = fsm_out == 1'd0;
wire _guard19483 = cond_wire634_out;
wire _guard19484 = _guard19482 & _guard19483;
wire _guard19485 = fsm_out == 1'd0;
wire _guard19486 = _guard19484 & _guard19485;
wire _guard19487 = _guard19481 | _guard19486;
wire _guard19488 = early_reset_static_par0_go_out;
wire _guard19489 = _guard19487 & _guard19488;
wire _guard19490 = cond_wire679_out;
wire _guard19491 = early_reset_static_par0_go_out;
wire _guard19492 = _guard19490 & _guard19491;
wire _guard19493 = cond_wire677_out;
wire _guard19494 = early_reset_static_par0_go_out;
wire _guard19495 = _guard19493 & _guard19494;
wire _guard19496 = fsm_out == 1'd0;
wire _guard19497 = cond_wire677_out;
wire _guard19498 = _guard19496 & _guard19497;
wire _guard19499 = fsm_out == 1'd0;
wire _guard19500 = _guard19498 & _guard19499;
wire _guard19501 = fsm_out == 1'd0;
wire _guard19502 = cond_wire679_out;
wire _guard19503 = _guard19501 & _guard19502;
wire _guard19504 = fsm_out == 1'd0;
wire _guard19505 = _guard19503 & _guard19504;
wire _guard19506 = _guard19500 | _guard19505;
wire _guard19507 = early_reset_static_par0_go_out;
wire _guard19508 = _guard19506 & _guard19507;
wire _guard19509 = fsm_out == 1'd0;
wire _guard19510 = cond_wire677_out;
wire _guard19511 = _guard19509 & _guard19510;
wire _guard19512 = fsm_out == 1'd0;
wire _guard19513 = _guard19511 & _guard19512;
wire _guard19514 = fsm_out == 1'd0;
wire _guard19515 = cond_wire679_out;
wire _guard19516 = _guard19514 & _guard19515;
wire _guard19517 = fsm_out == 1'd0;
wire _guard19518 = _guard19516 & _guard19517;
wire _guard19519 = _guard19513 | _guard19518;
wire _guard19520 = early_reset_static_par0_go_out;
wire _guard19521 = _guard19519 & _guard19520;
wire _guard19522 = fsm_out == 1'd0;
wire _guard19523 = cond_wire677_out;
wire _guard19524 = _guard19522 & _guard19523;
wire _guard19525 = fsm_out == 1'd0;
wire _guard19526 = _guard19524 & _guard19525;
wire _guard19527 = fsm_out == 1'd0;
wire _guard19528 = cond_wire679_out;
wire _guard19529 = _guard19527 & _guard19528;
wire _guard19530 = fsm_out == 1'd0;
wire _guard19531 = _guard19529 & _guard19530;
wire _guard19532 = _guard19526 | _guard19531;
wire _guard19533 = early_reset_static_par0_go_out;
wire _guard19534 = _guard19532 & _guard19533;
wire _guard19535 = cond_wire682_out;
wire _guard19536 = early_reset_static_par0_go_out;
wire _guard19537 = _guard19535 & _guard19536;
wire _guard19538 = cond_wire682_out;
wire _guard19539 = early_reset_static_par0_go_out;
wire _guard19540 = _guard19538 & _guard19539;
wire _guard19541 = cond_wire637_out;
wire _guard19542 = early_reset_static_par0_go_out;
wire _guard19543 = _guard19541 & _guard19542;
wire _guard19544 = cond_wire637_out;
wire _guard19545 = early_reset_static_par0_go_out;
wire _guard19546 = _guard19544 & _guard19545;
wire _guard19547 = cond_wire694_out;
wire _guard19548 = early_reset_static_par0_go_out;
wire _guard19549 = _guard19547 & _guard19548;
wire _guard19550 = cond_wire694_out;
wire _guard19551 = early_reset_static_par0_go_out;
wire _guard19552 = _guard19550 & _guard19551;
wire _guard19553 = cond_wire869_out;
wire _guard19554 = early_reset_static_par0_go_out;
wire _guard19555 = _guard19553 & _guard19554;
wire _guard19556 = cond_wire869_out;
wire _guard19557 = early_reset_static_par0_go_out;
wire _guard19558 = _guard19556 & _guard19557;
wire _guard19559 = cond_wire820_out;
wire _guard19560 = early_reset_static_par0_go_out;
wire _guard19561 = _guard19559 & _guard19560;
wire _guard19562 = cond_wire820_out;
wire _guard19563 = early_reset_static_par0_go_out;
wire _guard19564 = _guard19562 & _guard19563;
wire _guard19565 = cond_wire938_out;
wire _guard19566 = early_reset_static_par0_go_out;
wire _guard19567 = _guard19565 & _guard19566;
wire _guard19568 = cond_wire938_out;
wire _guard19569 = early_reset_static_par0_go_out;
wire _guard19570 = _guard19568 & _guard19569;
wire _guard19571 = cond_wire958_out;
wire _guard19572 = early_reset_static_par0_go_out;
wire _guard19573 = _guard19571 & _guard19572;
wire _guard19574 = cond_wire958_out;
wire _guard19575 = early_reset_static_par0_go_out;
wire _guard19576 = _guard19574 & _guard19575;
wire _guard19577 = cond_wire4_out;
wire _guard19578 = early_reset_static_par0_go_out;
wire _guard19579 = _guard19577 & _guard19578;
wire _guard19580 = cond_wire4_out;
wire _guard19581 = early_reset_static_par0_go_out;
wire _guard19582 = _guard19580 & _guard19581;
wire _guard19583 = fsm0_out == 6'd0;
wire _guard19584 = early_reset_static_seq_go_out;
wire _guard19585 = _guard19583 & _guard19584;
wire _guard19586 = cond_wire14_out;
wire _guard19587 = early_reset_static_par0_go_out;
wire _guard19588 = _guard19586 & _guard19587;
wire _guard19589 = _guard19585 | _guard19588;
wire _guard19590 = cond_wire14_out;
wire _guard19591 = early_reset_static_par0_go_out;
wire _guard19592 = _guard19590 & _guard19591;
wire _guard19593 = fsm0_out == 6'd0;
wire _guard19594 = early_reset_static_seq_go_out;
wire _guard19595 = _guard19593 & _guard19594;
wire _guard19596 = cond_wire59_out;
wire _guard19597 = early_reset_static_par0_go_out;
wire _guard19598 = _guard19596 & _guard19597;
wire _guard19599 = cond_wire59_out;
wire _guard19600 = early_reset_static_par0_go_out;
wire _guard19601 = _guard19599 & _guard19600;
wire _guard19602 = cond_wire274_out;
wire _guard19603 = early_reset_static_par0_go_out;
wire _guard19604 = _guard19602 & _guard19603;
wire _guard19605 = cond_wire274_out;
wire _guard19606 = early_reset_static_par0_go_out;
wire _guard19607 = _guard19605 & _guard19606;
wire _guard19608 = early_reset_static_par0_go_out;
wire _guard19609 = early_reset_static_par0_go_out;
wire _guard19610 = early_reset_static_par0_go_out;
wire _guard19611 = early_reset_static_par0_go_out;
wire _guard19612 = early_reset_static_par0_go_out;
wire _guard19613 = early_reset_static_par0_go_out;
wire _guard19614 = fsm0_out == 6'd0;
wire _guard19615 = early_reset_static_seq_go_out;
wire _guard19616 = _guard19614 & _guard19615;
wire _guard19617 = early_reset_static_par0_go_out;
wire _guard19618 = _guard19616 | _guard19617;
wire _guard19619 = early_reset_static_par0_go_out;
wire _guard19620 = fsm0_out == 6'd0;
wire _guard19621 = early_reset_static_seq_go_out;
wire _guard19622 = _guard19620 & _guard19621;
wire _guard19623 = fsm0_out == 6'd0;
wire _guard19624 = early_reset_static_seq_go_out;
wire _guard19625 = _guard19623 & _guard19624;
wire _guard19626 = early_reset_static_par0_go_out;
wire _guard19627 = _guard19625 | _guard19626;
wire _guard19628 = early_reset_static_par0_go_out;
wire _guard19629 = fsm0_out == 6'd0;
wire _guard19630 = early_reset_static_seq_go_out;
wire _guard19631 = _guard19629 & _guard19630;
wire _guard19632 = fsm0_out == 6'd0;
wire _guard19633 = early_reset_static_seq_go_out;
wire _guard19634 = _guard19632 & _guard19633;
wire _guard19635 = early_reset_static_par0_go_out;
wire _guard19636 = _guard19634 | _guard19635;
wire _guard19637 = early_reset_static_par0_go_out;
wire _guard19638 = fsm0_out == 6'd0;
wire _guard19639 = early_reset_static_seq_go_out;
wire _guard19640 = _guard19638 & _guard19639;
wire _guard19641 = fsm0_out == 6'd0;
wire _guard19642 = early_reset_static_seq_go_out;
wire _guard19643 = _guard19641 & _guard19642;
wire _guard19644 = early_reset_static_par0_go_out;
wire _guard19645 = _guard19643 | _guard19644;
wire _guard19646 = fsm0_out == 6'd0;
wire _guard19647 = early_reset_static_seq_go_out;
wire _guard19648 = _guard19646 & _guard19647;
wire _guard19649 = early_reset_static_par0_go_out;
wire _guard19650 = early_reset_static_par0_go_out;
wire _guard19651 = early_reset_static_par0_go_out;
wire _guard19652 = early_reset_static_par0_go_out;
wire _guard19653 = early_reset_static_par0_go_out;
wire _guard19654 = early_reset_static_par0_go_out;
wire _guard19655 = early_reset_static_par0_go_out;
wire _guard19656 = early_reset_static_par0_go_out;
wire _guard19657 = early_reset_static_par0_go_out;
wire _guard19658 = fsm0_out == 6'd0;
wire _guard19659 = early_reset_static_seq_go_out;
wire _guard19660 = _guard19658 & _guard19659;
wire _guard19661 = early_reset_static_par0_go_out;
wire _guard19662 = _guard19660 | _guard19661;
wire _guard19663 = early_reset_static_par0_go_out;
wire _guard19664 = fsm0_out == 6'd0;
wire _guard19665 = early_reset_static_seq_go_out;
wire _guard19666 = _guard19664 & _guard19665;
wire _guard19667 = early_reset_static_par0_go_out;
wire _guard19668 = early_reset_static_par0_go_out;
wire _guard19669 = early_reset_static_par0_go_out;
wire _guard19670 = early_reset_static_par0_go_out;
wire _guard19671 = early_reset_static_par0_go_out;
wire _guard19672 = early_reset_static_par0_go_out;
wire _guard19673 = early_reset_static_par0_go_out;
wire _guard19674 = early_reset_static_par0_go_out;
wire _guard19675 = early_reset_static_par0_go_out;
wire _guard19676 = early_reset_static_par0_go_out;
wire _guard19677 = fsm0_out == 6'd0;
wire _guard19678 = early_reset_static_seq_go_out;
wire _guard19679 = _guard19677 & _guard19678;
wire _guard19680 = early_reset_static_par0_go_out;
wire _guard19681 = _guard19679 | _guard19680;
wire _guard19682 = fsm0_out == 6'd0;
wire _guard19683 = early_reset_static_seq_go_out;
wire _guard19684 = _guard19682 & _guard19683;
wire _guard19685 = early_reset_static_par0_go_out;
wire _guard19686 = fsm0_out == 6'd0;
wire _guard19687 = early_reset_static_seq_go_out;
wire _guard19688 = _guard19686 & _guard19687;
wire _guard19689 = early_reset_static_par0_go_out;
wire _guard19690 = _guard19688 | _guard19689;
wire _guard19691 = early_reset_static_par0_go_out;
wire _guard19692 = fsm0_out == 6'd0;
wire _guard19693 = early_reset_static_seq_go_out;
wire _guard19694 = _guard19692 & _guard19693;
wire _guard19695 = fsm0_out == 6'd0;
wire _guard19696 = early_reset_static_seq_go_out;
wire _guard19697 = _guard19695 & _guard19696;
wire _guard19698 = early_reset_static_par0_go_out;
wire _guard19699 = _guard19697 | _guard19698;
wire _guard19700 = early_reset_static_par0_go_out;
wire _guard19701 = fsm0_out == 6'd0;
wire _guard19702 = early_reset_static_seq_go_out;
wire _guard19703 = _guard19701 & _guard19702;
wire _guard19704 = early_reset_static_par0_go_out;
wire _guard19705 = early_reset_static_par0_go_out;
wire _guard19706 = ~_guard0;
wire _guard19707 = early_reset_static_par0_go_out;
wire _guard19708 = _guard19706 & _guard19707;
wire _guard19709 = early_reset_static_par0_go_out;
wire _guard19710 = ~_guard0;
wire _guard19711 = early_reset_static_par0_go_out;
wire _guard19712 = _guard19710 & _guard19711;
wire _guard19713 = early_reset_static_par0_go_out;
wire _guard19714 = early_reset_static_par0_go_out;
wire _guard19715 = early_reset_static_par0_go_out;
wire _guard19716 = early_reset_static_par0_go_out;
wire _guard19717 = early_reset_static_par0_go_out;
wire _guard19718 = early_reset_static_par0_go_out;
wire _guard19719 = ~_guard0;
wire _guard19720 = early_reset_static_par0_go_out;
wire _guard19721 = _guard19719 & _guard19720;
wire _guard19722 = early_reset_static_par0_go_out;
wire _guard19723 = ~_guard0;
wire _guard19724 = early_reset_static_par0_go_out;
wire _guard19725 = _guard19723 & _guard19724;
wire _guard19726 = early_reset_static_par0_go_out;
wire _guard19727 = ~_guard0;
wire _guard19728 = early_reset_static_par0_go_out;
wire _guard19729 = _guard19727 & _guard19728;
wire _guard19730 = early_reset_static_par0_go_out;
wire _guard19731 = ~_guard0;
wire _guard19732 = early_reset_static_par0_go_out;
wire _guard19733 = _guard19731 & _guard19732;
wire _guard19734 = early_reset_static_par0_go_out;
wire _guard19735 = ~_guard0;
wire _guard19736 = early_reset_static_par0_go_out;
wire _guard19737 = _guard19735 & _guard19736;
wire _guard19738 = early_reset_static_par0_go_out;
wire _guard19739 = ~_guard0;
wire _guard19740 = early_reset_static_par0_go_out;
wire _guard19741 = _guard19739 & _guard19740;
wire _guard19742 = early_reset_static_par0_go_out;
wire _guard19743 = early_reset_static_par0_go_out;
wire _guard19744 = early_reset_static_par0_go_out;
wire _guard19745 = early_reset_static_par0_go_out;
wire _guard19746 = ~_guard0;
wire _guard19747 = early_reset_static_par0_go_out;
wire _guard19748 = _guard19746 & _guard19747;
wire _guard19749 = early_reset_static_par0_go_out;
wire _guard19750 = ~_guard0;
wire _guard19751 = early_reset_static_par0_go_out;
wire _guard19752 = _guard19750 & _guard19751;
wire _guard19753 = early_reset_static_par0_go_out;
wire _guard19754 = early_reset_static_par0_go_out;
wire _guard19755 = early_reset_static_par0_go_out;
wire _guard19756 = early_reset_static_par0_go_out;
wire _guard19757 = early_reset_static_par0_go_out;
wire _guard19758 = ~_guard0;
wire _guard19759 = early_reset_static_par0_go_out;
wire _guard19760 = _guard19758 & _guard19759;
wire _guard19761 = early_reset_static_par0_go_out;
wire _guard19762 = early_reset_static_par0_go_out;
wire _guard19763 = early_reset_static_par0_go_out;
wire _guard19764 = ~_guard0;
wire _guard19765 = early_reset_static_par0_go_out;
wire _guard19766 = _guard19764 & _guard19765;
wire _guard19767 = early_reset_static_par0_go_out;
wire _guard19768 = early_reset_static_par0_go_out;
wire _guard19769 = early_reset_static_par0_go_out;
wire _guard19770 = early_reset_static_par0_go_out;
wire _guard19771 = early_reset_static_par0_go_out;
wire _guard19772 = early_reset_static_par0_go_out;
wire _guard19773 = early_reset_static_par0_go_out;
wire _guard19774 = early_reset_static_par0_go_out;
wire _guard19775 = early_reset_static_par0_go_out;
wire _guard19776 = ~_guard0;
wire _guard19777 = early_reset_static_par0_go_out;
wire _guard19778 = _guard19776 & _guard19777;
wire _guard19779 = early_reset_static_par0_go_out;
wire _guard19780 = ~_guard0;
wire _guard19781 = early_reset_static_par0_go_out;
wire _guard19782 = _guard19780 & _guard19781;
wire _guard19783 = early_reset_static_par0_go_out;
wire _guard19784 = early_reset_static_par0_go_out;
wire _guard19785 = early_reset_static_par0_go_out;
wire _guard19786 = early_reset_static_par0_go_out;
wire _guard19787 = early_reset_static_par0_go_out;
wire _guard19788 = early_reset_static_par0_go_out;
wire _guard19789 = early_reset_static_par0_go_out;
wire _guard19790 = early_reset_static_par0_go_out;
wire _guard19791 = early_reset_static_par0_go_out;
wire _guard19792 = early_reset_static_par0_go_out;
wire _guard19793 = early_reset_static_par0_go_out;
wire _guard19794 = early_reset_static_par0_go_out;
wire _guard19795 = ~_guard0;
wire _guard19796 = early_reset_static_par0_go_out;
wire _guard19797 = _guard19795 & _guard19796;
wire _guard19798 = early_reset_static_par0_go_out;
wire _guard19799 = ~_guard0;
wire _guard19800 = early_reset_static_par0_go_out;
wire _guard19801 = _guard19799 & _guard19800;
wire _guard19802 = ~_guard0;
wire _guard19803 = early_reset_static_par0_go_out;
wire _guard19804 = _guard19802 & _guard19803;
wire _guard19805 = early_reset_static_par0_go_out;
wire _guard19806 = early_reset_static_par0_go_out;
wire _guard19807 = early_reset_static_par0_go_out;
wire _guard19808 = early_reset_static_par0_go_out;
wire _guard19809 = ~_guard0;
wire _guard19810 = early_reset_static_par0_go_out;
wire _guard19811 = _guard19809 & _guard19810;
wire _guard19812 = early_reset_static_par0_go_out;
wire _guard19813 = early_reset_static_par0_go_out;
wire _guard19814 = ~_guard0;
wire _guard19815 = early_reset_static_par0_go_out;
wire _guard19816 = _guard19814 & _guard19815;
wire _guard19817 = early_reset_static_par0_go_out;
wire _guard19818 = early_reset_static_par0_go_out;
wire _guard19819 = ~_guard0;
wire _guard19820 = early_reset_static_par0_go_out;
wire _guard19821 = _guard19819 & _guard19820;
wire _guard19822 = early_reset_static_par0_go_out;
wire _guard19823 = early_reset_static_par0_go_out;
wire _guard19824 = early_reset_static_par0_go_out;
wire _guard19825 = early_reset_static_par0_go_out;
wire _guard19826 = early_reset_static_par0_go_out;
wire _guard19827 = early_reset_static_par0_go_out;
wire _guard19828 = early_reset_static_par0_go_out;
wire _guard19829 = early_reset_static_par0_go_out;
wire _guard19830 = ~_guard0;
wire _guard19831 = early_reset_static_par0_go_out;
wire _guard19832 = _guard19830 & _guard19831;
wire _guard19833 = early_reset_static_par0_go_out;
wire _guard19834 = ~_guard0;
wire _guard19835 = early_reset_static_par0_go_out;
wire _guard19836 = _guard19834 & _guard19835;
wire _guard19837 = early_reset_static_par0_go_out;
wire _guard19838 = early_reset_static_par0_go_out;
wire _guard19839 = early_reset_static_par0_go_out;
wire _guard19840 = early_reset_static_par0_go_out;
wire _guard19841 = ~_guard0;
wire _guard19842 = early_reset_static_par0_go_out;
wire _guard19843 = _guard19841 & _guard19842;
wire _guard19844 = early_reset_static_par0_go_out;
wire _guard19845 = ~_guard0;
wire _guard19846 = early_reset_static_par0_go_out;
wire _guard19847 = _guard19845 & _guard19846;
wire _guard19848 = early_reset_static_par0_go_out;
wire _guard19849 = early_reset_static_par0_go_out;
wire _guard19850 = ~_guard0;
wire _guard19851 = early_reset_static_par0_go_out;
wire _guard19852 = _guard19850 & _guard19851;
wire _guard19853 = early_reset_static_par0_go_out;
wire _guard19854 = early_reset_static_par0_go_out;
wire _guard19855 = early_reset_static_par0_go_out;
wire _guard19856 = ~_guard0;
wire _guard19857 = early_reset_static_par0_go_out;
wire _guard19858 = _guard19856 & _guard19857;
wire _guard19859 = early_reset_static_par0_go_out;
wire _guard19860 = early_reset_static_par0_go_out;
wire _guard19861 = ~_guard0;
wire _guard19862 = early_reset_static_par0_go_out;
wire _guard19863 = _guard19861 & _guard19862;
wire _guard19864 = early_reset_static_par0_go_out;
wire _guard19865 = early_reset_static_par0_go_out;
wire _guard19866 = early_reset_static_par0_go_out;
wire _guard19867 = early_reset_static_par0_go_out;
wire _guard19868 = early_reset_static_par0_go_out;
wire _guard19869 = early_reset_static_par0_go_out;
wire _guard19870 = early_reset_static_par0_go_out;
wire _guard19871 = early_reset_static_par0_go_out;
wire _guard19872 = early_reset_static_par0_go_out;
wire _guard19873 = early_reset_static_par0_go_out;
wire _guard19874 = early_reset_static_par0_go_out;
wire _guard19875 = early_reset_static_par0_go_out;
wire _guard19876 = ~_guard0;
wire _guard19877 = early_reset_static_par0_go_out;
wire _guard19878 = _guard19876 & _guard19877;
wire _guard19879 = early_reset_static_par0_go_out;
wire _guard19880 = early_reset_static_par0_go_out;
wire _guard19881 = early_reset_static_par0_go_out;
wire _guard19882 = early_reset_static_par0_go_out;
wire _guard19883 = early_reset_static_par0_go_out;
wire _guard19884 = early_reset_static_par0_go_out;
wire _guard19885 = ~_guard0;
wire _guard19886 = early_reset_static_par0_go_out;
wire _guard19887 = _guard19885 & _guard19886;
wire _guard19888 = ~_guard0;
wire _guard19889 = early_reset_static_par0_go_out;
wire _guard19890 = _guard19888 & _guard19889;
wire _guard19891 = early_reset_static_par0_go_out;
wire _guard19892 = early_reset_static_par0_go_out;
wire _guard19893 = early_reset_static_par0_go_out;
wire _guard19894 = ~_guard0;
wire _guard19895 = early_reset_static_par0_go_out;
wire _guard19896 = _guard19894 & _guard19895;
wire _guard19897 = early_reset_static_par0_go_out;
wire _guard19898 = ~_guard0;
wire _guard19899 = early_reset_static_par0_go_out;
wire _guard19900 = _guard19898 & _guard19899;
wire _guard19901 = early_reset_static_par0_go_out;
wire _guard19902 = ~_guard0;
wire _guard19903 = early_reset_static_par0_go_out;
wire _guard19904 = _guard19902 & _guard19903;
wire _guard19905 = early_reset_static_par0_go_out;
wire _guard19906 = early_reset_static_par0_go_out;
wire _guard19907 = ~_guard0;
wire _guard19908 = early_reset_static_par0_go_out;
wire _guard19909 = _guard19907 & _guard19908;
wire _guard19910 = early_reset_static_par0_go_out;
wire _guard19911 = early_reset_static_par0_go_out;
wire _guard19912 = early_reset_static_par0_go_out;
wire _guard19913 = ~_guard0;
wire _guard19914 = early_reset_static_par0_go_out;
wire _guard19915 = _guard19913 & _guard19914;
wire _guard19916 = early_reset_static_par0_go_out;
wire _guard19917 = early_reset_static_par0_go_out;
wire _guard19918 = early_reset_static_par0_go_out;
wire _guard19919 = early_reset_static_par0_go_out;
wire _guard19920 = ~_guard0;
wire _guard19921 = early_reset_static_par0_go_out;
wire _guard19922 = _guard19920 & _guard19921;
wire _guard19923 = early_reset_static_par0_go_out;
wire _guard19924 = early_reset_static_par0_go_out;
wire _guard19925 = ~_guard0;
wire _guard19926 = early_reset_static_par0_go_out;
wire _guard19927 = _guard19925 & _guard19926;
wire _guard19928 = early_reset_static_par0_go_out;
wire _guard19929 = early_reset_static_par0_go_out;
wire _guard19930 = early_reset_static_par0_go_out;
wire _guard19931 = ~_guard0;
wire _guard19932 = early_reset_static_par0_go_out;
wire _guard19933 = _guard19931 & _guard19932;
wire _guard19934 = early_reset_static_par0_go_out;
wire _guard19935 = early_reset_static_par0_go_out;
wire _guard19936 = early_reset_static_par0_go_out;
wire _guard19937 = early_reset_static_par0_go_out;
wire _guard19938 = early_reset_static_par0_go_out;
wire _guard19939 = ~_guard0;
wire _guard19940 = early_reset_static_par0_go_out;
wire _guard19941 = _guard19939 & _guard19940;
wire _guard19942 = early_reset_static_par0_go_out;
wire _guard19943 = ~_guard0;
wire _guard19944 = early_reset_static_par0_go_out;
wire _guard19945 = _guard19943 & _guard19944;
wire _guard19946 = early_reset_static_par0_go_out;
wire _guard19947 = early_reset_static_par0_go_out;
wire _guard19948 = early_reset_static_par0_go_out;
wire _guard19949 = early_reset_static_par0_go_out;
wire _guard19950 = early_reset_static_par0_go_out;
wire _guard19951 = ~_guard0;
wire _guard19952 = early_reset_static_par0_go_out;
wire _guard19953 = _guard19951 & _guard19952;
wire _guard19954 = early_reset_static_par0_go_out;
wire _guard19955 = early_reset_static_par0_go_out;
wire _guard19956 = early_reset_static_par0_go_out;
wire _guard19957 = ~_guard0;
wire _guard19958 = early_reset_static_par0_go_out;
wire _guard19959 = _guard19957 & _guard19958;
wire _guard19960 = ~_guard0;
wire _guard19961 = early_reset_static_par0_go_out;
wire _guard19962 = _guard19960 & _guard19961;
wire _guard19963 = early_reset_static_par0_go_out;
wire _guard19964 = early_reset_static_par0_go_out;
wire _guard19965 = early_reset_static_par0_go_out;
wire _guard19966 = early_reset_static_par0_go_out;
wire _guard19967 = ~_guard0;
wire _guard19968 = early_reset_static_par0_go_out;
wire _guard19969 = _guard19967 & _guard19968;
wire _guard19970 = early_reset_static_par0_go_out;
wire _guard19971 = ~_guard0;
wire _guard19972 = early_reset_static_par0_go_out;
wire _guard19973 = _guard19971 & _guard19972;
wire _guard19974 = early_reset_static_par0_go_out;
wire _guard19975 = early_reset_static_par0_go_out;
wire _guard19976 = early_reset_static_par0_go_out;
wire _guard19977 = early_reset_static_par0_go_out;
wire _guard19978 = early_reset_static_par0_go_out;
wire _guard19979 = ~_guard0;
wire _guard19980 = early_reset_static_par0_go_out;
wire _guard19981 = _guard19979 & _guard19980;
wire _guard19982 = early_reset_static_par0_go_out;
wire _guard19983 = early_reset_static_par0_go_out;
wire _guard19984 = early_reset_static_par0_go_out;
wire _guard19985 = ~_guard0;
wire _guard19986 = early_reset_static_par0_go_out;
wire _guard19987 = _guard19985 & _guard19986;
wire _guard19988 = early_reset_static_par0_go_out;
wire _guard19989 = ~_guard0;
wire _guard19990 = early_reset_static_par0_go_out;
wire _guard19991 = _guard19989 & _guard19990;
wire _guard19992 = early_reset_static_par0_go_out;
wire _guard19993 = early_reset_static_par0_go_out;
wire _guard19994 = early_reset_static_par0_go_out;
wire _guard19995 = early_reset_static_par0_go_out;
wire _guard19996 = early_reset_static_par0_go_out;
wire _guard19997 = early_reset_static_par0_go_out;
wire _guard19998 = early_reset_static_par0_go_out;
wire _guard19999 = early_reset_static_par0_go_out;
wire _guard20000 = ~_guard0;
wire _guard20001 = early_reset_static_par0_go_out;
wire _guard20002 = _guard20000 & _guard20001;
wire _guard20003 = early_reset_static_par0_go_out;
wire _guard20004 = early_reset_static_par0_go_out;
wire _guard20005 = early_reset_static_par0_go_out;
wire _guard20006 = early_reset_static_par0_go_out;
wire _guard20007 = ~_guard0;
wire _guard20008 = early_reset_static_par0_go_out;
wire _guard20009 = _guard20007 & _guard20008;
wire _guard20010 = early_reset_static_par0_go_out;
wire _guard20011 = early_reset_static_par0_go_out;
wire _guard20012 = early_reset_static_par0_go_out;
wire _guard20013 = early_reset_static_par0_go_out;
wire _guard20014 = early_reset_static_par0_go_out;
wire _guard20015 = ~_guard0;
wire _guard20016 = early_reset_static_par0_go_out;
wire _guard20017 = _guard20015 & _guard20016;
wire _guard20018 = early_reset_static_par0_go_out;
wire _guard20019 = early_reset_static_par0_go_out;
wire _guard20020 = early_reset_static_par0_go_out;
wire _guard20021 = ~_guard0;
wire _guard20022 = early_reset_static_par0_go_out;
wire _guard20023 = _guard20021 & _guard20022;
wire _guard20024 = early_reset_static_par0_go_out;
wire _guard20025 = early_reset_static_par0_go_out;
wire _guard20026 = early_reset_static_par0_go_out;
wire _guard20027 = early_reset_static_par0_go_out;
wire _guard20028 = ~_guard0;
wire _guard20029 = early_reset_static_par0_go_out;
wire _guard20030 = _guard20028 & _guard20029;
wire _guard20031 = early_reset_static_par0_go_out;
wire _guard20032 = early_reset_static_par0_go_out;
wire _guard20033 = early_reset_static_par0_go_out;
wire _guard20034 = ~_guard0;
wire _guard20035 = early_reset_static_par0_go_out;
wire _guard20036 = _guard20034 & _guard20035;
wire _guard20037 = early_reset_static_par0_go_out;
wire _guard20038 = early_reset_static_par0_go_out;
wire _guard20039 = early_reset_static_par0_go_out;
wire _guard20040 = ~_guard0;
wire _guard20041 = early_reset_static_par0_go_out;
wire _guard20042 = _guard20040 & _guard20041;
wire _guard20043 = early_reset_static_par0_go_out;
wire _guard20044 = early_reset_static_par0_go_out;
wire _guard20045 = ~_guard0;
wire _guard20046 = early_reset_static_par0_go_out;
wire _guard20047 = _guard20045 & _guard20046;
wire _guard20048 = early_reset_static_par0_go_out;
wire _guard20049 = early_reset_static_par0_go_out;
wire _guard20050 = ~_guard0;
wire _guard20051 = early_reset_static_par0_go_out;
wire _guard20052 = _guard20050 & _guard20051;
wire _guard20053 = early_reset_static_par0_go_out;
wire _guard20054 = early_reset_static_par0_go_out;
wire _guard20055 = early_reset_static_par0_go_out;
wire _guard20056 = early_reset_static_par0_go_out;
wire _guard20057 = ~_guard0;
wire _guard20058 = early_reset_static_par0_go_out;
wire _guard20059 = _guard20057 & _guard20058;
wire _guard20060 = early_reset_static_par0_go_out;
wire _guard20061 = early_reset_static_par0_go_out;
wire _guard20062 = early_reset_static_par0_go_out;
wire _guard20063 = early_reset_static_par0_go_out;
wire _guard20064 = ~_guard0;
wire _guard20065 = early_reset_static_par0_go_out;
wire _guard20066 = _guard20064 & _guard20065;
wire _guard20067 = early_reset_static_par0_go_out;
wire _guard20068 = early_reset_static_par0_go_out;
wire _guard20069 = early_reset_static_par0_go_out;
wire _guard20070 = early_reset_static_par0_go_out;
wire _guard20071 = early_reset_static_par0_go_out;
wire _guard20072 = early_reset_static_par0_go_out;
wire _guard20073 = ~_guard0;
wire _guard20074 = early_reset_static_par0_go_out;
wire _guard20075 = _guard20073 & _guard20074;
wire _guard20076 = early_reset_static_par0_go_out;
wire _guard20077 = early_reset_static_par0_go_out;
wire _guard20078 = ~_guard0;
wire _guard20079 = early_reset_static_par0_go_out;
wire _guard20080 = _guard20078 & _guard20079;
wire _guard20081 = early_reset_static_par0_go_out;
wire _guard20082 = early_reset_static_par0_go_out;
wire _guard20083 = early_reset_static_par0_go_out;
wire _guard20084 = early_reset_static_par0_go_out;
wire _guard20085 = early_reset_static_par0_go_out;
wire _guard20086 = early_reset_static_par0_go_out;
wire _guard20087 = early_reset_static_par0_go_out;
wire _guard20088 = ~_guard0;
wire _guard20089 = early_reset_static_par0_go_out;
wire _guard20090 = _guard20088 & _guard20089;
wire _guard20091 = early_reset_static_par0_go_out;
wire _guard20092 = ~_guard0;
wire _guard20093 = early_reset_static_par0_go_out;
wire _guard20094 = _guard20092 & _guard20093;
wire _guard20095 = early_reset_static_par0_go_out;
wire _guard20096 = early_reset_static_par0_go_out;
wire _guard20097 = early_reset_static_par0_go_out;
wire _guard20098 = early_reset_static_par0_go_out;
wire _guard20099 = early_reset_static_par0_go_out;
wire _guard20100 = cond_wire2_out;
wire _guard20101 = early_reset_static_par0_go_out;
wire _guard20102 = _guard20100 & _guard20101;
wire _guard20103 = cond_wire0_out;
wire _guard20104 = early_reset_static_par0_go_out;
wire _guard20105 = _guard20103 & _guard20104;
wire _guard20106 = fsm_out == 1'd0;
wire _guard20107 = cond_wire0_out;
wire _guard20108 = _guard20106 & _guard20107;
wire _guard20109 = fsm_out == 1'd0;
wire _guard20110 = _guard20108 & _guard20109;
wire _guard20111 = fsm_out == 1'd0;
wire _guard20112 = cond_wire2_out;
wire _guard20113 = _guard20111 & _guard20112;
wire _guard20114 = fsm_out == 1'd0;
wire _guard20115 = _guard20113 & _guard20114;
wire _guard20116 = _guard20110 | _guard20115;
wire _guard20117 = early_reset_static_par0_go_out;
wire _guard20118 = _guard20116 & _guard20117;
wire _guard20119 = fsm_out == 1'd0;
wire _guard20120 = cond_wire0_out;
wire _guard20121 = _guard20119 & _guard20120;
wire _guard20122 = fsm_out == 1'd0;
wire _guard20123 = _guard20121 & _guard20122;
wire _guard20124 = fsm_out == 1'd0;
wire _guard20125 = cond_wire2_out;
wire _guard20126 = _guard20124 & _guard20125;
wire _guard20127 = fsm_out == 1'd0;
wire _guard20128 = _guard20126 & _guard20127;
wire _guard20129 = _guard20123 | _guard20128;
wire _guard20130 = early_reset_static_par0_go_out;
wire _guard20131 = _guard20129 & _guard20130;
wire _guard20132 = fsm_out == 1'd0;
wire _guard20133 = cond_wire0_out;
wire _guard20134 = _guard20132 & _guard20133;
wire _guard20135 = fsm_out == 1'd0;
wire _guard20136 = _guard20134 & _guard20135;
wire _guard20137 = fsm_out == 1'd0;
wire _guard20138 = cond_wire2_out;
wire _guard20139 = _guard20137 & _guard20138;
wire _guard20140 = fsm_out == 1'd0;
wire _guard20141 = _guard20139 & _guard20140;
wire _guard20142 = _guard20136 | _guard20141;
wire _guard20143 = early_reset_static_par0_go_out;
wire _guard20144 = _guard20142 & _guard20143;
wire _guard20145 = cond_wire61_out;
wire _guard20146 = early_reset_static_par0_go_out;
wire _guard20147 = _guard20145 & _guard20146;
wire _guard20148 = cond_wire61_out;
wire _guard20149 = early_reset_static_par0_go_out;
wire _guard20150 = _guard20148 & _guard20149;
wire _guard20151 = cond_wire101_out;
wire _guard20152 = early_reset_static_par0_go_out;
wire _guard20153 = _guard20151 & _guard20152;
wire _guard20154 = cond_wire101_out;
wire _guard20155 = early_reset_static_par0_go_out;
wire _guard20156 = _guard20154 & _guard20155;
wire _guard20157 = cond_wire109_out;
wire _guard20158 = early_reset_static_par0_go_out;
wire _guard20159 = _guard20157 & _guard20158;
wire _guard20160 = cond_wire109_out;
wire _guard20161 = early_reset_static_par0_go_out;
wire _guard20162 = _guard20160 & _guard20161;
wire _guard20163 = cond_wire71_out;
wire _guard20164 = early_reset_static_par0_go_out;
wire _guard20165 = _guard20163 & _guard20164;
wire _guard20166 = cond_wire71_out;
wire _guard20167 = early_reset_static_par0_go_out;
wire _guard20168 = _guard20166 & _guard20167;
wire _guard20169 = cond_wire113_out;
wire _guard20170 = early_reset_static_par0_go_out;
wire _guard20171 = _guard20169 & _guard20170;
wire _guard20172 = cond_wire113_out;
wire _guard20173 = early_reset_static_par0_go_out;
wire _guard20174 = _guard20172 & _guard20173;
wire _guard20175 = cond_wire182_out;
wire _guard20176 = early_reset_static_par0_go_out;
wire _guard20177 = _guard20175 & _guard20176;
wire _guard20178 = cond_wire182_out;
wire _guard20179 = early_reset_static_par0_go_out;
wire _guard20180 = _guard20178 & _guard20179;
wire _guard20181 = cond_wire224_out;
wire _guard20182 = early_reset_static_par0_go_out;
wire _guard20183 = _guard20181 & _guard20182;
wire _guard20184 = cond_wire222_out;
wire _guard20185 = early_reset_static_par0_go_out;
wire _guard20186 = _guard20184 & _guard20185;
wire _guard20187 = fsm_out == 1'd0;
wire _guard20188 = cond_wire222_out;
wire _guard20189 = _guard20187 & _guard20188;
wire _guard20190 = fsm_out == 1'd0;
wire _guard20191 = _guard20189 & _guard20190;
wire _guard20192 = fsm_out == 1'd0;
wire _guard20193 = cond_wire224_out;
wire _guard20194 = _guard20192 & _guard20193;
wire _guard20195 = fsm_out == 1'd0;
wire _guard20196 = _guard20194 & _guard20195;
wire _guard20197 = _guard20191 | _guard20196;
wire _guard20198 = early_reset_static_par0_go_out;
wire _guard20199 = _guard20197 & _guard20198;
wire _guard20200 = fsm_out == 1'd0;
wire _guard20201 = cond_wire222_out;
wire _guard20202 = _guard20200 & _guard20201;
wire _guard20203 = fsm_out == 1'd0;
wire _guard20204 = _guard20202 & _guard20203;
wire _guard20205 = fsm_out == 1'd0;
wire _guard20206 = cond_wire224_out;
wire _guard20207 = _guard20205 & _guard20206;
wire _guard20208 = fsm_out == 1'd0;
wire _guard20209 = _guard20207 & _guard20208;
wire _guard20210 = _guard20204 | _guard20209;
wire _guard20211 = early_reset_static_par0_go_out;
wire _guard20212 = _guard20210 & _guard20211;
wire _guard20213 = fsm_out == 1'd0;
wire _guard20214 = cond_wire222_out;
wire _guard20215 = _guard20213 & _guard20214;
wire _guard20216 = fsm_out == 1'd0;
wire _guard20217 = _guard20215 & _guard20216;
wire _guard20218 = fsm_out == 1'd0;
wire _guard20219 = cond_wire224_out;
wire _guard20220 = _guard20218 & _guard20219;
wire _guard20221 = fsm_out == 1'd0;
wire _guard20222 = _guard20220 & _guard20221;
wire _guard20223 = _guard20217 | _guard20222;
wire _guard20224 = early_reset_static_par0_go_out;
wire _guard20225 = _guard20223 & _guard20224;
wire _guard20226 = cond_wire158_out;
wire _guard20227 = early_reset_static_par0_go_out;
wire _guard20228 = _guard20226 & _guard20227;
wire _guard20229 = cond_wire158_out;
wire _guard20230 = early_reset_static_par0_go_out;
wire _guard20231 = _guard20229 & _guard20230;
wire _guard20232 = cond_wire247_out;
wire _guard20233 = early_reset_static_par0_go_out;
wire _guard20234 = _guard20232 & _guard20233;
wire _guard20235 = cond_wire247_out;
wire _guard20236 = early_reset_static_par0_go_out;
wire _guard20237 = _guard20235 & _guard20236;
wire _guard20238 = cond_wire263_out;
wire _guard20239 = early_reset_static_par0_go_out;
wire _guard20240 = _guard20238 & _guard20239;
wire _guard20241 = cond_wire263_out;
wire _guard20242 = early_reset_static_par0_go_out;
wire _guard20243 = _guard20241 & _guard20242;
wire _guard20244 = cond_wire223_out;
wire _guard20245 = early_reset_static_par0_go_out;
wire _guard20246 = _guard20244 & _guard20245;
wire _guard20247 = cond_wire223_out;
wire _guard20248 = early_reset_static_par0_go_out;
wire _guard20249 = _guard20247 & _guard20248;
wire _guard20250 = cond_wire235_out;
wire _guard20251 = early_reset_static_par0_go_out;
wire _guard20252 = _guard20250 & _guard20251;
wire _guard20253 = cond_wire235_out;
wire _guard20254 = early_reset_static_par0_go_out;
wire _guard20255 = _guard20253 & _guard20254;
wire _guard20256 = cond_wire366_out;
wire _guard20257 = early_reset_static_par0_go_out;
wire _guard20258 = _guard20256 & _guard20257;
wire _guard20259 = cond_wire364_out;
wire _guard20260 = early_reset_static_par0_go_out;
wire _guard20261 = _guard20259 & _guard20260;
wire _guard20262 = fsm_out == 1'd0;
wire _guard20263 = cond_wire364_out;
wire _guard20264 = _guard20262 & _guard20263;
wire _guard20265 = fsm_out == 1'd0;
wire _guard20266 = _guard20264 & _guard20265;
wire _guard20267 = fsm_out == 1'd0;
wire _guard20268 = cond_wire366_out;
wire _guard20269 = _guard20267 & _guard20268;
wire _guard20270 = fsm_out == 1'd0;
wire _guard20271 = _guard20269 & _guard20270;
wire _guard20272 = _guard20266 | _guard20271;
wire _guard20273 = early_reset_static_par0_go_out;
wire _guard20274 = _guard20272 & _guard20273;
wire _guard20275 = fsm_out == 1'd0;
wire _guard20276 = cond_wire364_out;
wire _guard20277 = _guard20275 & _guard20276;
wire _guard20278 = fsm_out == 1'd0;
wire _guard20279 = _guard20277 & _guard20278;
wire _guard20280 = fsm_out == 1'd0;
wire _guard20281 = cond_wire366_out;
wire _guard20282 = _guard20280 & _guard20281;
wire _guard20283 = fsm_out == 1'd0;
wire _guard20284 = _guard20282 & _guard20283;
wire _guard20285 = _guard20279 | _guard20284;
wire _guard20286 = early_reset_static_par0_go_out;
wire _guard20287 = _guard20285 & _guard20286;
wire _guard20288 = fsm_out == 1'd0;
wire _guard20289 = cond_wire364_out;
wire _guard20290 = _guard20288 & _guard20289;
wire _guard20291 = fsm_out == 1'd0;
wire _guard20292 = _guard20290 & _guard20291;
wire _guard20293 = fsm_out == 1'd0;
wire _guard20294 = cond_wire366_out;
wire _guard20295 = _guard20293 & _guard20294;
wire _guard20296 = fsm_out == 1'd0;
wire _guard20297 = _guard20295 & _guard20296;
wire _guard20298 = _guard20292 | _guard20297;
wire _guard20299 = early_reset_static_par0_go_out;
wire _guard20300 = _guard20298 & _guard20299;
wire _guard20301 = cond_wire300_out;
wire _guard20302 = early_reset_static_par0_go_out;
wire _guard20303 = _guard20301 & _guard20302;
wire _guard20304 = cond_wire300_out;
wire _guard20305 = early_reset_static_par0_go_out;
wire _guard20306 = _guard20304 & _guard20305;
wire _guard20307 = cond_wire349_out;
wire _guard20308 = early_reset_static_par0_go_out;
wire _guard20309 = _guard20307 & _guard20308;
wire _guard20310 = cond_wire349_out;
wire _guard20311 = early_reset_static_par0_go_out;
wire _guard20312 = _guard20310 & _guard20311;
wire _guard20313 = cond_wire438_out;
wire _guard20314 = early_reset_static_par0_go_out;
wire _guard20315 = _guard20313 & _guard20314;
wire _guard20316 = cond_wire438_out;
wire _guard20317 = early_reset_static_par0_go_out;
wire _guard20318 = _guard20316 & _guard20317;
wire _guard20319 = cond_wire401_out;
wire _guard20320 = early_reset_static_par0_go_out;
wire _guard20321 = _guard20319 & _guard20320;
wire _guard20322 = cond_wire401_out;
wire _guard20323 = early_reset_static_par0_go_out;
wire _guard20324 = _guard20322 & _guard20323;
wire _guard20325 = cond_wire476_out;
wire _guard20326 = early_reset_static_par0_go_out;
wire _guard20327 = _guard20325 & _guard20326;
wire _guard20328 = cond_wire474_out;
wire _guard20329 = early_reset_static_par0_go_out;
wire _guard20330 = _guard20328 & _guard20329;
wire _guard20331 = fsm_out == 1'd0;
wire _guard20332 = cond_wire474_out;
wire _guard20333 = _guard20331 & _guard20332;
wire _guard20334 = fsm_out == 1'd0;
wire _guard20335 = _guard20333 & _guard20334;
wire _guard20336 = fsm_out == 1'd0;
wire _guard20337 = cond_wire476_out;
wire _guard20338 = _guard20336 & _guard20337;
wire _guard20339 = fsm_out == 1'd0;
wire _guard20340 = _guard20338 & _guard20339;
wire _guard20341 = _guard20335 | _guard20340;
wire _guard20342 = early_reset_static_par0_go_out;
wire _guard20343 = _guard20341 & _guard20342;
wire _guard20344 = fsm_out == 1'd0;
wire _guard20345 = cond_wire474_out;
wire _guard20346 = _guard20344 & _guard20345;
wire _guard20347 = fsm_out == 1'd0;
wire _guard20348 = _guard20346 & _guard20347;
wire _guard20349 = fsm_out == 1'd0;
wire _guard20350 = cond_wire476_out;
wire _guard20351 = _guard20349 & _guard20350;
wire _guard20352 = fsm_out == 1'd0;
wire _guard20353 = _guard20351 & _guard20352;
wire _guard20354 = _guard20348 | _guard20353;
wire _guard20355 = early_reset_static_par0_go_out;
wire _guard20356 = _guard20354 & _guard20355;
wire _guard20357 = fsm_out == 1'd0;
wire _guard20358 = cond_wire474_out;
wire _guard20359 = _guard20357 & _guard20358;
wire _guard20360 = fsm_out == 1'd0;
wire _guard20361 = _guard20359 & _guard20360;
wire _guard20362 = fsm_out == 1'd0;
wire _guard20363 = cond_wire476_out;
wire _guard20364 = _guard20362 & _guard20363;
wire _guard20365 = fsm_out == 1'd0;
wire _guard20366 = _guard20364 & _guard20365;
wire _guard20367 = _guard20361 | _guard20366;
wire _guard20368 = early_reset_static_par0_go_out;
wire _guard20369 = _guard20367 & _guard20368;
wire _guard20370 = cond_wire520_out;
wire _guard20371 = early_reset_static_par0_go_out;
wire _guard20372 = _guard20370 & _guard20371;
wire _guard20373 = cond_wire518_out;
wire _guard20374 = early_reset_static_par0_go_out;
wire _guard20375 = _guard20373 & _guard20374;
wire _guard20376 = fsm_out == 1'd0;
wire _guard20377 = cond_wire518_out;
wire _guard20378 = _guard20376 & _guard20377;
wire _guard20379 = fsm_out == 1'd0;
wire _guard20380 = _guard20378 & _guard20379;
wire _guard20381 = fsm_out == 1'd0;
wire _guard20382 = cond_wire520_out;
wire _guard20383 = _guard20381 & _guard20382;
wire _guard20384 = fsm_out == 1'd0;
wire _guard20385 = _guard20383 & _guard20384;
wire _guard20386 = _guard20380 | _guard20385;
wire _guard20387 = early_reset_static_par0_go_out;
wire _guard20388 = _guard20386 & _guard20387;
wire _guard20389 = fsm_out == 1'd0;
wire _guard20390 = cond_wire518_out;
wire _guard20391 = _guard20389 & _guard20390;
wire _guard20392 = fsm_out == 1'd0;
wire _guard20393 = _guard20391 & _guard20392;
wire _guard20394 = fsm_out == 1'd0;
wire _guard20395 = cond_wire520_out;
wire _guard20396 = _guard20394 & _guard20395;
wire _guard20397 = fsm_out == 1'd0;
wire _guard20398 = _guard20396 & _guard20397;
wire _guard20399 = _guard20393 | _guard20398;
wire _guard20400 = early_reset_static_par0_go_out;
wire _guard20401 = _guard20399 & _guard20400;
wire _guard20402 = fsm_out == 1'd0;
wire _guard20403 = cond_wire518_out;
wire _guard20404 = _guard20402 & _guard20403;
wire _guard20405 = fsm_out == 1'd0;
wire _guard20406 = _guard20404 & _guard20405;
wire _guard20407 = fsm_out == 1'd0;
wire _guard20408 = cond_wire520_out;
wire _guard20409 = _guard20407 & _guard20408;
wire _guard20410 = fsm_out == 1'd0;
wire _guard20411 = _guard20409 & _guard20410;
wire _guard20412 = _guard20406 | _guard20411;
wire _guard20413 = early_reset_static_par0_go_out;
wire _guard20414 = _guard20412 & _guard20413;
wire _guard20415 = cond_wire519_out;
wire _guard20416 = early_reset_static_par0_go_out;
wire _guard20417 = _guard20415 & _guard20416;
wire _guard20418 = cond_wire519_out;
wire _guard20419 = early_reset_static_par0_go_out;
wire _guard20420 = _guard20418 & _guard20419;
wire _guard20421 = cond_wire549_out;
wire _guard20422 = early_reset_static_par0_go_out;
wire _guard20423 = _guard20421 & _guard20422;
wire _guard20424 = cond_wire547_out;
wire _guard20425 = early_reset_static_par0_go_out;
wire _guard20426 = _guard20424 & _guard20425;
wire _guard20427 = fsm_out == 1'd0;
wire _guard20428 = cond_wire547_out;
wire _guard20429 = _guard20427 & _guard20428;
wire _guard20430 = fsm_out == 1'd0;
wire _guard20431 = _guard20429 & _guard20430;
wire _guard20432 = fsm_out == 1'd0;
wire _guard20433 = cond_wire549_out;
wire _guard20434 = _guard20432 & _guard20433;
wire _guard20435 = fsm_out == 1'd0;
wire _guard20436 = _guard20434 & _guard20435;
wire _guard20437 = _guard20431 | _guard20436;
wire _guard20438 = early_reset_static_par0_go_out;
wire _guard20439 = _guard20437 & _guard20438;
wire _guard20440 = fsm_out == 1'd0;
wire _guard20441 = cond_wire547_out;
wire _guard20442 = _guard20440 & _guard20441;
wire _guard20443 = fsm_out == 1'd0;
wire _guard20444 = _guard20442 & _guard20443;
wire _guard20445 = fsm_out == 1'd0;
wire _guard20446 = cond_wire549_out;
wire _guard20447 = _guard20445 & _guard20446;
wire _guard20448 = fsm_out == 1'd0;
wire _guard20449 = _guard20447 & _guard20448;
wire _guard20450 = _guard20444 | _guard20449;
wire _guard20451 = early_reset_static_par0_go_out;
wire _guard20452 = _guard20450 & _guard20451;
wire _guard20453 = fsm_out == 1'd0;
wire _guard20454 = cond_wire547_out;
wire _guard20455 = _guard20453 & _guard20454;
wire _guard20456 = fsm_out == 1'd0;
wire _guard20457 = _guard20455 & _guard20456;
wire _guard20458 = fsm_out == 1'd0;
wire _guard20459 = cond_wire549_out;
wire _guard20460 = _guard20458 & _guard20459;
wire _guard20461 = fsm_out == 1'd0;
wire _guard20462 = _guard20460 & _guard20461;
wire _guard20463 = _guard20457 | _guard20462;
wire _guard20464 = early_reset_static_par0_go_out;
wire _guard20465 = _guard20463 & _guard20464;
wire _guard20466 = cond_wire585_out;
wire _guard20467 = early_reset_static_par0_go_out;
wire _guard20468 = _guard20466 & _guard20467;
wire _guard20469 = cond_wire583_out;
wire _guard20470 = early_reset_static_par0_go_out;
wire _guard20471 = _guard20469 & _guard20470;
wire _guard20472 = fsm_out == 1'd0;
wire _guard20473 = cond_wire583_out;
wire _guard20474 = _guard20472 & _guard20473;
wire _guard20475 = fsm_out == 1'd0;
wire _guard20476 = _guard20474 & _guard20475;
wire _guard20477 = fsm_out == 1'd0;
wire _guard20478 = cond_wire585_out;
wire _guard20479 = _guard20477 & _guard20478;
wire _guard20480 = fsm_out == 1'd0;
wire _guard20481 = _guard20479 & _guard20480;
wire _guard20482 = _guard20476 | _guard20481;
wire _guard20483 = early_reset_static_par0_go_out;
wire _guard20484 = _guard20482 & _guard20483;
wire _guard20485 = fsm_out == 1'd0;
wire _guard20486 = cond_wire583_out;
wire _guard20487 = _guard20485 & _guard20486;
wire _guard20488 = fsm_out == 1'd0;
wire _guard20489 = _guard20487 & _guard20488;
wire _guard20490 = fsm_out == 1'd0;
wire _guard20491 = cond_wire585_out;
wire _guard20492 = _guard20490 & _guard20491;
wire _guard20493 = fsm_out == 1'd0;
wire _guard20494 = _guard20492 & _guard20493;
wire _guard20495 = _guard20489 | _guard20494;
wire _guard20496 = early_reset_static_par0_go_out;
wire _guard20497 = _guard20495 & _guard20496;
wire _guard20498 = fsm_out == 1'd0;
wire _guard20499 = cond_wire583_out;
wire _guard20500 = _guard20498 & _guard20499;
wire _guard20501 = fsm_out == 1'd0;
wire _guard20502 = _guard20500 & _guard20501;
wire _guard20503 = fsm_out == 1'd0;
wire _guard20504 = cond_wire585_out;
wire _guard20505 = _guard20503 & _guard20504;
wire _guard20506 = fsm_out == 1'd0;
wire _guard20507 = _guard20505 & _guard20506;
wire _guard20508 = _guard20502 | _guard20507;
wire _guard20509 = early_reset_static_par0_go_out;
wire _guard20510 = _guard20508 & _guard20509;
wire _guard20511 = cond_wire599_out;
wire _guard20512 = early_reset_static_par0_go_out;
wire _guard20513 = _guard20511 & _guard20512;
wire _guard20514 = cond_wire599_out;
wire _guard20515 = early_reset_static_par0_go_out;
wire _guard20516 = _guard20514 & _guard20515;
wire _guard20517 = cond_wire580_out;
wire _guard20518 = early_reset_static_par0_go_out;
wire _guard20519 = _guard20517 & _guard20518;
wire _guard20520 = cond_wire580_out;
wire _guard20521 = early_reset_static_par0_go_out;
wire _guard20522 = _guard20520 & _guard20521;
wire _guard20523 = cond_wire645_out;
wire _guard20524 = early_reset_static_par0_go_out;
wire _guard20525 = _guard20523 & _guard20524;
wire _guard20526 = cond_wire645_out;
wire _guard20527 = early_reset_static_par0_go_out;
wire _guard20528 = _guard20526 & _guard20527;
wire _guard20529 = cond_wire658_out;
wire _guard20530 = early_reset_static_par0_go_out;
wire _guard20531 = _guard20529 & _guard20530;
wire _guard20532 = cond_wire656_out;
wire _guard20533 = early_reset_static_par0_go_out;
wire _guard20534 = _guard20532 & _guard20533;
wire _guard20535 = fsm_out == 1'd0;
wire _guard20536 = cond_wire656_out;
wire _guard20537 = _guard20535 & _guard20536;
wire _guard20538 = fsm_out == 1'd0;
wire _guard20539 = _guard20537 & _guard20538;
wire _guard20540 = fsm_out == 1'd0;
wire _guard20541 = cond_wire658_out;
wire _guard20542 = _guard20540 & _guard20541;
wire _guard20543 = fsm_out == 1'd0;
wire _guard20544 = _guard20542 & _guard20543;
wire _guard20545 = _guard20539 | _guard20544;
wire _guard20546 = early_reset_static_par0_go_out;
wire _guard20547 = _guard20545 & _guard20546;
wire _guard20548 = fsm_out == 1'd0;
wire _guard20549 = cond_wire656_out;
wire _guard20550 = _guard20548 & _guard20549;
wire _guard20551 = fsm_out == 1'd0;
wire _guard20552 = _guard20550 & _guard20551;
wire _guard20553 = fsm_out == 1'd0;
wire _guard20554 = cond_wire658_out;
wire _guard20555 = _guard20553 & _guard20554;
wire _guard20556 = fsm_out == 1'd0;
wire _guard20557 = _guard20555 & _guard20556;
wire _guard20558 = _guard20552 | _guard20557;
wire _guard20559 = early_reset_static_par0_go_out;
wire _guard20560 = _guard20558 & _guard20559;
wire _guard20561 = fsm_out == 1'd0;
wire _guard20562 = cond_wire656_out;
wire _guard20563 = _guard20561 & _guard20562;
wire _guard20564 = fsm_out == 1'd0;
wire _guard20565 = _guard20563 & _guard20564;
wire _guard20566 = fsm_out == 1'd0;
wire _guard20567 = cond_wire658_out;
wire _guard20568 = _guard20566 & _guard20567;
wire _guard20569 = fsm_out == 1'd0;
wire _guard20570 = _guard20568 & _guard20569;
wire _guard20571 = _guard20565 | _guard20570;
wire _guard20572 = early_reset_static_par0_go_out;
wire _guard20573 = _guard20571 & _guard20572;
wire _guard20574 = cond_wire670_out;
wire _guard20575 = early_reset_static_par0_go_out;
wire _guard20576 = _guard20574 & _guard20575;
wire _guard20577 = cond_wire670_out;
wire _guard20578 = early_reset_static_par0_go_out;
wire _guard20579 = _guard20577 & _guard20578;
wire _guard20580 = cond_wire683_out;
wire _guard20581 = early_reset_static_par0_go_out;
wire _guard20582 = _guard20580 & _guard20581;
wire _guard20583 = cond_wire681_out;
wire _guard20584 = early_reset_static_par0_go_out;
wire _guard20585 = _guard20583 & _guard20584;
wire _guard20586 = fsm_out == 1'd0;
wire _guard20587 = cond_wire681_out;
wire _guard20588 = _guard20586 & _guard20587;
wire _guard20589 = fsm_out == 1'd0;
wire _guard20590 = _guard20588 & _guard20589;
wire _guard20591 = fsm_out == 1'd0;
wire _guard20592 = cond_wire683_out;
wire _guard20593 = _guard20591 & _guard20592;
wire _guard20594 = fsm_out == 1'd0;
wire _guard20595 = _guard20593 & _guard20594;
wire _guard20596 = _guard20590 | _guard20595;
wire _guard20597 = early_reset_static_par0_go_out;
wire _guard20598 = _guard20596 & _guard20597;
wire _guard20599 = fsm_out == 1'd0;
wire _guard20600 = cond_wire681_out;
wire _guard20601 = _guard20599 & _guard20600;
wire _guard20602 = fsm_out == 1'd0;
wire _guard20603 = _guard20601 & _guard20602;
wire _guard20604 = fsm_out == 1'd0;
wire _guard20605 = cond_wire683_out;
wire _guard20606 = _guard20604 & _guard20605;
wire _guard20607 = fsm_out == 1'd0;
wire _guard20608 = _guard20606 & _guard20607;
wire _guard20609 = _guard20603 | _guard20608;
wire _guard20610 = early_reset_static_par0_go_out;
wire _guard20611 = _guard20609 & _guard20610;
wire _guard20612 = fsm_out == 1'd0;
wire _guard20613 = cond_wire681_out;
wire _guard20614 = _guard20612 & _guard20613;
wire _guard20615 = fsm_out == 1'd0;
wire _guard20616 = _guard20614 & _guard20615;
wire _guard20617 = fsm_out == 1'd0;
wire _guard20618 = cond_wire683_out;
wire _guard20619 = _guard20617 & _guard20618;
wire _guard20620 = fsm_out == 1'd0;
wire _guard20621 = _guard20619 & _guard20620;
wire _guard20622 = _guard20616 | _guard20621;
wire _guard20623 = early_reset_static_par0_go_out;
wire _guard20624 = _guard20622 & _guard20623;
wire _guard20625 = cond_wire617_out;
wire _guard20626 = early_reset_static_par0_go_out;
wire _guard20627 = _guard20625 & _guard20626;
wire _guard20628 = cond_wire617_out;
wire _guard20629 = early_reset_static_par0_go_out;
wire _guard20630 = _guard20628 & _guard20629;
wire _guard20631 = cond_wire727_out;
wire _guard20632 = early_reset_static_par0_go_out;
wire _guard20633 = _guard20631 & _guard20632;
wire _guard20634 = cond_wire725_out;
wire _guard20635 = early_reset_static_par0_go_out;
wire _guard20636 = _guard20634 & _guard20635;
wire _guard20637 = fsm_out == 1'd0;
wire _guard20638 = cond_wire725_out;
wire _guard20639 = _guard20637 & _guard20638;
wire _guard20640 = fsm_out == 1'd0;
wire _guard20641 = _guard20639 & _guard20640;
wire _guard20642 = fsm_out == 1'd0;
wire _guard20643 = cond_wire727_out;
wire _guard20644 = _guard20642 & _guard20643;
wire _guard20645 = fsm_out == 1'd0;
wire _guard20646 = _guard20644 & _guard20645;
wire _guard20647 = _guard20641 | _guard20646;
wire _guard20648 = early_reset_static_par0_go_out;
wire _guard20649 = _guard20647 & _guard20648;
wire _guard20650 = fsm_out == 1'd0;
wire _guard20651 = cond_wire725_out;
wire _guard20652 = _guard20650 & _guard20651;
wire _guard20653 = fsm_out == 1'd0;
wire _guard20654 = _guard20652 & _guard20653;
wire _guard20655 = fsm_out == 1'd0;
wire _guard20656 = cond_wire727_out;
wire _guard20657 = _guard20655 & _guard20656;
wire _guard20658 = fsm_out == 1'd0;
wire _guard20659 = _guard20657 & _guard20658;
wire _guard20660 = _guard20654 | _guard20659;
wire _guard20661 = early_reset_static_par0_go_out;
wire _guard20662 = _guard20660 & _guard20661;
wire _guard20663 = fsm_out == 1'd0;
wire _guard20664 = cond_wire725_out;
wire _guard20665 = _guard20663 & _guard20664;
wire _guard20666 = fsm_out == 1'd0;
wire _guard20667 = _guard20665 & _guard20666;
wire _guard20668 = fsm_out == 1'd0;
wire _guard20669 = cond_wire727_out;
wire _guard20670 = _guard20668 & _guard20669;
wire _guard20671 = fsm_out == 1'd0;
wire _guard20672 = _guard20670 & _guard20671;
wire _guard20673 = _guard20667 | _guard20672;
wire _guard20674 = early_reset_static_par0_go_out;
wire _guard20675 = _guard20673 & _guard20674;
wire _guard20676 = cond_wire661_out;
wire _guard20677 = early_reset_static_par0_go_out;
wire _guard20678 = _guard20676 & _guard20677;
wire _guard20679 = cond_wire661_out;
wire _guard20680 = early_reset_static_par0_go_out;
wire _guard20681 = _guard20679 & _guard20680;
wire _guard20682 = cond_wire682_out;
wire _guard20683 = early_reset_static_par0_go_out;
wire _guard20684 = _guard20682 & _guard20683;
wire _guard20685 = cond_wire682_out;
wire _guard20686 = early_reset_static_par0_go_out;
wire _guard20687 = _guard20685 & _guard20686;
wire _guard20688 = cond_wire751_out;
wire _guard20689 = early_reset_static_par0_go_out;
wire _guard20690 = _guard20688 & _guard20689;
wire _guard20691 = cond_wire751_out;
wire _guard20692 = early_reset_static_par0_go_out;
wire _guard20693 = _guard20691 & _guard20692;
wire _guard20694 = cond_wire702_out;
wire _guard20695 = early_reset_static_par0_go_out;
wire _guard20696 = _guard20694 & _guard20695;
wire _guard20697 = cond_wire702_out;
wire _guard20698 = early_reset_static_par0_go_out;
wire _guard20699 = _guard20697 & _guard20698;
wire _guard20700 = cond_wire706_out;
wire _guard20701 = early_reset_static_par0_go_out;
wire _guard20702 = _guard20700 & _guard20701;
wire _guard20703 = cond_wire706_out;
wire _guard20704 = early_reset_static_par0_go_out;
wire _guard20705 = _guard20703 & _guard20704;
wire _guard20706 = cond_wire784_out;
wire _guard20707 = early_reset_static_par0_go_out;
wire _guard20708 = _guard20706 & _guard20707;
wire _guard20709 = cond_wire782_out;
wire _guard20710 = early_reset_static_par0_go_out;
wire _guard20711 = _guard20709 & _guard20710;
wire _guard20712 = fsm_out == 1'd0;
wire _guard20713 = cond_wire782_out;
wire _guard20714 = _guard20712 & _guard20713;
wire _guard20715 = fsm_out == 1'd0;
wire _guard20716 = _guard20714 & _guard20715;
wire _guard20717 = fsm_out == 1'd0;
wire _guard20718 = cond_wire784_out;
wire _guard20719 = _guard20717 & _guard20718;
wire _guard20720 = fsm_out == 1'd0;
wire _guard20721 = _guard20719 & _guard20720;
wire _guard20722 = _guard20716 | _guard20721;
wire _guard20723 = early_reset_static_par0_go_out;
wire _guard20724 = _guard20722 & _guard20723;
wire _guard20725 = fsm_out == 1'd0;
wire _guard20726 = cond_wire782_out;
wire _guard20727 = _guard20725 & _guard20726;
wire _guard20728 = fsm_out == 1'd0;
wire _guard20729 = _guard20727 & _guard20728;
wire _guard20730 = fsm_out == 1'd0;
wire _guard20731 = cond_wire784_out;
wire _guard20732 = _guard20730 & _guard20731;
wire _guard20733 = fsm_out == 1'd0;
wire _guard20734 = _guard20732 & _guard20733;
wire _guard20735 = _guard20729 | _guard20734;
wire _guard20736 = early_reset_static_par0_go_out;
wire _guard20737 = _guard20735 & _guard20736;
wire _guard20738 = fsm_out == 1'd0;
wire _guard20739 = cond_wire782_out;
wire _guard20740 = _guard20738 & _guard20739;
wire _guard20741 = fsm_out == 1'd0;
wire _guard20742 = _guard20740 & _guard20741;
wire _guard20743 = fsm_out == 1'd0;
wire _guard20744 = cond_wire784_out;
wire _guard20745 = _guard20743 & _guard20744;
wire _guard20746 = fsm_out == 1'd0;
wire _guard20747 = _guard20745 & _guard20746;
wire _guard20748 = _guard20742 | _guard20747;
wire _guard20749 = early_reset_static_par0_go_out;
wire _guard20750 = _guard20748 & _guard20749;
wire _guard20751 = cond_wire788_out;
wire _guard20752 = early_reset_static_par0_go_out;
wire _guard20753 = _guard20751 & _guard20752;
wire _guard20754 = cond_wire786_out;
wire _guard20755 = early_reset_static_par0_go_out;
wire _guard20756 = _guard20754 & _guard20755;
wire _guard20757 = fsm_out == 1'd0;
wire _guard20758 = cond_wire786_out;
wire _guard20759 = _guard20757 & _guard20758;
wire _guard20760 = fsm_out == 1'd0;
wire _guard20761 = _guard20759 & _guard20760;
wire _guard20762 = fsm_out == 1'd0;
wire _guard20763 = cond_wire788_out;
wire _guard20764 = _guard20762 & _guard20763;
wire _guard20765 = fsm_out == 1'd0;
wire _guard20766 = _guard20764 & _guard20765;
wire _guard20767 = _guard20761 | _guard20766;
wire _guard20768 = early_reset_static_par0_go_out;
wire _guard20769 = _guard20767 & _guard20768;
wire _guard20770 = fsm_out == 1'd0;
wire _guard20771 = cond_wire786_out;
wire _guard20772 = _guard20770 & _guard20771;
wire _guard20773 = fsm_out == 1'd0;
wire _guard20774 = _guard20772 & _guard20773;
wire _guard20775 = fsm_out == 1'd0;
wire _guard20776 = cond_wire788_out;
wire _guard20777 = _guard20775 & _guard20776;
wire _guard20778 = fsm_out == 1'd0;
wire _guard20779 = _guard20777 & _guard20778;
wire _guard20780 = _guard20774 | _guard20779;
wire _guard20781 = early_reset_static_par0_go_out;
wire _guard20782 = _guard20780 & _guard20781;
wire _guard20783 = fsm_out == 1'd0;
wire _guard20784 = cond_wire786_out;
wire _guard20785 = _guard20783 & _guard20784;
wire _guard20786 = fsm_out == 1'd0;
wire _guard20787 = _guard20785 & _guard20786;
wire _guard20788 = fsm_out == 1'd0;
wire _guard20789 = cond_wire788_out;
wire _guard20790 = _guard20788 & _guard20789;
wire _guard20791 = fsm_out == 1'd0;
wire _guard20792 = _guard20790 & _guard20791;
wire _guard20793 = _guard20787 | _guard20792;
wire _guard20794 = early_reset_static_par0_go_out;
wire _guard20795 = _guard20793 & _guard20794;
wire _guard20796 = cond_wire800_out;
wire _guard20797 = early_reset_static_par0_go_out;
wire _guard20798 = _guard20796 & _guard20797;
wire _guard20799 = cond_wire800_out;
wire _guard20800 = early_reset_static_par0_go_out;
wire _guard20801 = _guard20799 & _guard20800;
wire _guard20802 = cond_wire817_out;
wire _guard20803 = early_reset_static_par0_go_out;
wire _guard20804 = _guard20802 & _guard20803;
wire _guard20805 = cond_wire815_out;
wire _guard20806 = early_reset_static_par0_go_out;
wire _guard20807 = _guard20805 & _guard20806;
wire _guard20808 = fsm_out == 1'd0;
wire _guard20809 = cond_wire815_out;
wire _guard20810 = _guard20808 & _guard20809;
wire _guard20811 = fsm_out == 1'd0;
wire _guard20812 = _guard20810 & _guard20811;
wire _guard20813 = fsm_out == 1'd0;
wire _guard20814 = cond_wire817_out;
wire _guard20815 = _guard20813 & _guard20814;
wire _guard20816 = fsm_out == 1'd0;
wire _guard20817 = _guard20815 & _guard20816;
wire _guard20818 = _guard20812 | _guard20817;
wire _guard20819 = early_reset_static_par0_go_out;
wire _guard20820 = _guard20818 & _guard20819;
wire _guard20821 = fsm_out == 1'd0;
wire _guard20822 = cond_wire815_out;
wire _guard20823 = _guard20821 & _guard20822;
wire _guard20824 = fsm_out == 1'd0;
wire _guard20825 = _guard20823 & _guard20824;
wire _guard20826 = fsm_out == 1'd0;
wire _guard20827 = cond_wire817_out;
wire _guard20828 = _guard20826 & _guard20827;
wire _guard20829 = fsm_out == 1'd0;
wire _guard20830 = _guard20828 & _guard20829;
wire _guard20831 = _guard20825 | _guard20830;
wire _guard20832 = early_reset_static_par0_go_out;
wire _guard20833 = _guard20831 & _guard20832;
wire _guard20834 = fsm_out == 1'd0;
wire _guard20835 = cond_wire815_out;
wire _guard20836 = _guard20834 & _guard20835;
wire _guard20837 = fsm_out == 1'd0;
wire _guard20838 = _guard20836 & _guard20837;
wire _guard20839 = fsm_out == 1'd0;
wire _guard20840 = cond_wire817_out;
wire _guard20841 = _guard20839 & _guard20840;
wire _guard20842 = fsm_out == 1'd0;
wire _guard20843 = _guard20841 & _guard20842;
wire _guard20844 = _guard20838 | _guard20843;
wire _guard20845 = early_reset_static_par0_go_out;
wire _guard20846 = _guard20844 & _guard20845;
wire _guard20847 = cond_wire816_out;
wire _guard20848 = early_reset_static_par0_go_out;
wire _guard20849 = _guard20847 & _guard20848;
wire _guard20850 = cond_wire816_out;
wire _guard20851 = early_reset_static_par0_go_out;
wire _guard20852 = _guard20850 & _guard20851;
wire _guard20853 = cond_wire820_out;
wire _guard20854 = early_reset_static_par0_go_out;
wire _guard20855 = _guard20853 & _guard20854;
wire _guard20856 = cond_wire820_out;
wire _guard20857 = early_reset_static_par0_go_out;
wire _guard20858 = _guard20856 & _guard20857;
wire _guard20859 = cond_wire849_out;
wire _guard20860 = early_reset_static_par0_go_out;
wire _guard20861 = _guard20859 & _guard20860;
wire _guard20862 = cond_wire847_out;
wire _guard20863 = early_reset_static_par0_go_out;
wire _guard20864 = _guard20862 & _guard20863;
wire _guard20865 = fsm_out == 1'd0;
wire _guard20866 = cond_wire847_out;
wire _guard20867 = _guard20865 & _guard20866;
wire _guard20868 = fsm_out == 1'd0;
wire _guard20869 = _guard20867 & _guard20868;
wire _guard20870 = fsm_out == 1'd0;
wire _guard20871 = cond_wire849_out;
wire _guard20872 = _guard20870 & _guard20871;
wire _guard20873 = fsm_out == 1'd0;
wire _guard20874 = _guard20872 & _guard20873;
wire _guard20875 = _guard20869 | _guard20874;
wire _guard20876 = early_reset_static_par0_go_out;
wire _guard20877 = _guard20875 & _guard20876;
wire _guard20878 = fsm_out == 1'd0;
wire _guard20879 = cond_wire847_out;
wire _guard20880 = _guard20878 & _guard20879;
wire _guard20881 = fsm_out == 1'd0;
wire _guard20882 = _guard20880 & _guard20881;
wire _guard20883 = fsm_out == 1'd0;
wire _guard20884 = cond_wire849_out;
wire _guard20885 = _guard20883 & _guard20884;
wire _guard20886 = fsm_out == 1'd0;
wire _guard20887 = _guard20885 & _guard20886;
wire _guard20888 = _guard20882 | _guard20887;
wire _guard20889 = early_reset_static_par0_go_out;
wire _guard20890 = _guard20888 & _guard20889;
wire _guard20891 = fsm_out == 1'd0;
wire _guard20892 = cond_wire847_out;
wire _guard20893 = _guard20891 & _guard20892;
wire _guard20894 = fsm_out == 1'd0;
wire _guard20895 = _guard20893 & _guard20894;
wire _guard20896 = fsm_out == 1'd0;
wire _guard20897 = cond_wire849_out;
wire _guard20898 = _guard20896 & _guard20897;
wire _guard20899 = fsm_out == 1'd0;
wire _guard20900 = _guard20898 & _guard20899;
wire _guard20901 = _guard20895 | _guard20900;
wire _guard20902 = early_reset_static_par0_go_out;
wire _guard20903 = _guard20901 & _guard20902;
wire _guard20904 = cond_wire857_out;
wire _guard20905 = early_reset_static_par0_go_out;
wire _guard20906 = _guard20904 & _guard20905;
wire _guard20907 = cond_wire855_out;
wire _guard20908 = early_reset_static_par0_go_out;
wire _guard20909 = _guard20907 & _guard20908;
wire _guard20910 = fsm_out == 1'd0;
wire _guard20911 = cond_wire855_out;
wire _guard20912 = _guard20910 & _guard20911;
wire _guard20913 = fsm_out == 1'd0;
wire _guard20914 = _guard20912 & _guard20913;
wire _guard20915 = fsm_out == 1'd0;
wire _guard20916 = cond_wire857_out;
wire _guard20917 = _guard20915 & _guard20916;
wire _guard20918 = fsm_out == 1'd0;
wire _guard20919 = _guard20917 & _guard20918;
wire _guard20920 = _guard20914 | _guard20919;
wire _guard20921 = early_reset_static_par0_go_out;
wire _guard20922 = _guard20920 & _guard20921;
wire _guard20923 = fsm_out == 1'd0;
wire _guard20924 = cond_wire855_out;
wire _guard20925 = _guard20923 & _guard20924;
wire _guard20926 = fsm_out == 1'd0;
wire _guard20927 = _guard20925 & _guard20926;
wire _guard20928 = fsm_out == 1'd0;
wire _guard20929 = cond_wire857_out;
wire _guard20930 = _guard20928 & _guard20929;
wire _guard20931 = fsm_out == 1'd0;
wire _guard20932 = _guard20930 & _guard20931;
wire _guard20933 = _guard20927 | _guard20932;
wire _guard20934 = early_reset_static_par0_go_out;
wire _guard20935 = _guard20933 & _guard20934;
wire _guard20936 = fsm_out == 1'd0;
wire _guard20937 = cond_wire855_out;
wire _guard20938 = _guard20936 & _guard20937;
wire _guard20939 = fsm_out == 1'd0;
wire _guard20940 = _guard20938 & _guard20939;
wire _guard20941 = fsm_out == 1'd0;
wire _guard20942 = cond_wire857_out;
wire _guard20943 = _guard20941 & _guard20942;
wire _guard20944 = fsm_out == 1'd0;
wire _guard20945 = _guard20943 & _guard20944;
wire _guard20946 = _guard20940 | _guard20945;
wire _guard20947 = early_reset_static_par0_go_out;
wire _guard20948 = _guard20946 & _guard20947;
wire _guard20949 = cond_wire791_out;
wire _guard20950 = early_reset_static_par0_go_out;
wire _guard20951 = _guard20949 & _guard20950;
wire _guard20952 = cond_wire791_out;
wire _guard20953 = early_reset_static_par0_go_out;
wire _guard20954 = _guard20952 & _guard20953;
wire _guard20955 = cond_wire873_out;
wire _guard20956 = early_reset_static_par0_go_out;
wire _guard20957 = _guard20955 & _guard20956;
wire _guard20958 = cond_wire873_out;
wire _guard20959 = early_reset_static_par0_go_out;
wire _guard20960 = _guard20958 & _guard20959;
wire _guard20961 = cond_wire898_out;
wire _guard20962 = early_reset_static_par0_go_out;
wire _guard20963 = _guard20961 & _guard20962;
wire _guard20964 = cond_wire896_out;
wire _guard20965 = early_reset_static_par0_go_out;
wire _guard20966 = _guard20964 & _guard20965;
wire _guard20967 = fsm_out == 1'd0;
wire _guard20968 = cond_wire896_out;
wire _guard20969 = _guard20967 & _guard20968;
wire _guard20970 = fsm_out == 1'd0;
wire _guard20971 = _guard20969 & _guard20970;
wire _guard20972 = fsm_out == 1'd0;
wire _guard20973 = cond_wire898_out;
wire _guard20974 = _guard20972 & _guard20973;
wire _guard20975 = fsm_out == 1'd0;
wire _guard20976 = _guard20974 & _guard20975;
wire _guard20977 = _guard20971 | _guard20976;
wire _guard20978 = early_reset_static_par0_go_out;
wire _guard20979 = _guard20977 & _guard20978;
wire _guard20980 = fsm_out == 1'd0;
wire _guard20981 = cond_wire896_out;
wire _guard20982 = _guard20980 & _guard20981;
wire _guard20983 = fsm_out == 1'd0;
wire _guard20984 = _guard20982 & _guard20983;
wire _guard20985 = fsm_out == 1'd0;
wire _guard20986 = cond_wire898_out;
wire _guard20987 = _guard20985 & _guard20986;
wire _guard20988 = fsm_out == 1'd0;
wire _guard20989 = _guard20987 & _guard20988;
wire _guard20990 = _guard20984 | _guard20989;
wire _guard20991 = early_reset_static_par0_go_out;
wire _guard20992 = _guard20990 & _guard20991;
wire _guard20993 = fsm_out == 1'd0;
wire _guard20994 = cond_wire896_out;
wire _guard20995 = _guard20993 & _guard20994;
wire _guard20996 = fsm_out == 1'd0;
wire _guard20997 = _guard20995 & _guard20996;
wire _guard20998 = fsm_out == 1'd0;
wire _guard20999 = cond_wire898_out;
wire _guard21000 = _guard20998 & _guard20999;
wire _guard21001 = fsm_out == 1'd0;
wire _guard21002 = _guard21000 & _guard21001;
wire _guard21003 = _guard20997 | _guard21002;
wire _guard21004 = early_reset_static_par0_go_out;
wire _guard21005 = _guard21003 & _guard21004;
wire _guard21006 = cond_wire939_out;
wire _guard21007 = early_reset_static_par0_go_out;
wire _guard21008 = _guard21006 & _guard21007;
wire _guard21009 = cond_wire937_out;
wire _guard21010 = early_reset_static_par0_go_out;
wire _guard21011 = _guard21009 & _guard21010;
wire _guard21012 = fsm_out == 1'd0;
wire _guard21013 = cond_wire937_out;
wire _guard21014 = _guard21012 & _guard21013;
wire _guard21015 = fsm_out == 1'd0;
wire _guard21016 = _guard21014 & _guard21015;
wire _guard21017 = fsm_out == 1'd0;
wire _guard21018 = cond_wire939_out;
wire _guard21019 = _guard21017 & _guard21018;
wire _guard21020 = fsm_out == 1'd0;
wire _guard21021 = _guard21019 & _guard21020;
wire _guard21022 = _guard21016 | _guard21021;
wire _guard21023 = early_reset_static_par0_go_out;
wire _guard21024 = _guard21022 & _guard21023;
wire _guard21025 = fsm_out == 1'd0;
wire _guard21026 = cond_wire937_out;
wire _guard21027 = _guard21025 & _guard21026;
wire _guard21028 = fsm_out == 1'd0;
wire _guard21029 = _guard21027 & _guard21028;
wire _guard21030 = fsm_out == 1'd0;
wire _guard21031 = cond_wire939_out;
wire _guard21032 = _guard21030 & _guard21031;
wire _guard21033 = fsm_out == 1'd0;
wire _guard21034 = _guard21032 & _guard21033;
wire _guard21035 = _guard21029 | _guard21034;
wire _guard21036 = early_reset_static_par0_go_out;
wire _guard21037 = _guard21035 & _guard21036;
wire _guard21038 = fsm_out == 1'd0;
wire _guard21039 = cond_wire937_out;
wire _guard21040 = _guard21038 & _guard21039;
wire _guard21041 = fsm_out == 1'd0;
wire _guard21042 = _guard21040 & _guard21041;
wire _guard21043 = fsm_out == 1'd0;
wire _guard21044 = cond_wire939_out;
wire _guard21045 = _guard21043 & _guard21044;
wire _guard21046 = fsm_out == 1'd0;
wire _guard21047 = _guard21045 & _guard21046;
wire _guard21048 = _guard21042 | _guard21047;
wire _guard21049 = early_reset_static_par0_go_out;
wire _guard21050 = _guard21048 & _guard21049;
wire _guard21051 = cond_wire885_out;
wire _guard21052 = early_reset_static_par0_go_out;
wire _guard21053 = _guard21051 & _guard21052;
wire _guard21054 = cond_wire885_out;
wire _guard21055 = early_reset_static_par0_go_out;
wire _guard21056 = _guard21054 & _guard21055;
wire _guard21057 = cond_wire967_out;
wire _guard21058 = early_reset_static_par0_go_out;
wire _guard21059 = _guard21057 & _guard21058;
wire _guard21060 = cond_wire965_out;
wire _guard21061 = early_reset_static_par0_go_out;
wire _guard21062 = _guard21060 & _guard21061;
wire _guard21063 = fsm_out == 1'd0;
wire _guard21064 = cond_wire965_out;
wire _guard21065 = _guard21063 & _guard21064;
wire _guard21066 = fsm_out == 1'd0;
wire _guard21067 = _guard21065 & _guard21066;
wire _guard21068 = fsm_out == 1'd0;
wire _guard21069 = cond_wire967_out;
wire _guard21070 = _guard21068 & _guard21069;
wire _guard21071 = fsm_out == 1'd0;
wire _guard21072 = _guard21070 & _guard21071;
wire _guard21073 = _guard21067 | _guard21072;
wire _guard21074 = early_reset_static_par0_go_out;
wire _guard21075 = _guard21073 & _guard21074;
wire _guard21076 = fsm_out == 1'd0;
wire _guard21077 = cond_wire965_out;
wire _guard21078 = _guard21076 & _guard21077;
wire _guard21079 = fsm_out == 1'd0;
wire _guard21080 = _guard21078 & _guard21079;
wire _guard21081 = fsm_out == 1'd0;
wire _guard21082 = cond_wire967_out;
wire _guard21083 = _guard21081 & _guard21082;
wire _guard21084 = fsm_out == 1'd0;
wire _guard21085 = _guard21083 & _guard21084;
wire _guard21086 = _guard21080 | _guard21085;
wire _guard21087 = early_reset_static_par0_go_out;
wire _guard21088 = _guard21086 & _guard21087;
wire _guard21089 = fsm_out == 1'd0;
wire _guard21090 = cond_wire965_out;
wire _guard21091 = _guard21089 & _guard21090;
wire _guard21092 = fsm_out == 1'd0;
wire _guard21093 = _guard21091 & _guard21092;
wire _guard21094 = fsm_out == 1'd0;
wire _guard21095 = cond_wire967_out;
wire _guard21096 = _guard21094 & _guard21095;
wire _guard21097 = fsm_out == 1'd0;
wire _guard21098 = _guard21096 & _guard21097;
wire _guard21099 = _guard21093 | _guard21098;
wire _guard21100 = early_reset_static_par0_go_out;
wire _guard21101 = _guard21099 & _guard21100;
wire _guard21102 = cond_wire978_out;
wire _guard21103 = early_reset_static_par0_go_out;
wire _guard21104 = _guard21102 & _guard21103;
wire _guard21105 = cond_wire978_out;
wire _guard21106 = early_reset_static_par0_go_out;
wire _guard21107 = _guard21105 & _guard21106;
wire _guard21108 = cond_wire991_out;
wire _guard21109 = early_reset_static_par0_go_out;
wire _guard21110 = _guard21108 & _guard21109;
wire _guard21111 = cond_wire991_out;
wire _guard21112 = early_reset_static_par0_go_out;
wire _guard21113 = _guard21111 & _guard21112;
wire _guard21114 = cond_wire934_out;
wire _guard21115 = early_reset_static_par0_go_out;
wire _guard21116 = _guard21114 & _guard21115;
wire _guard21117 = cond_wire934_out;
wire _guard21118 = early_reset_static_par0_go_out;
wire _guard21119 = _guard21117 & _guard21118;
wire _guard21120 = cond_wire1004_out;
wire _guard21121 = early_reset_static_par0_go_out;
wire _guard21122 = _guard21120 & _guard21121;
wire _guard21123 = cond_wire1002_out;
wire _guard21124 = early_reset_static_par0_go_out;
wire _guard21125 = _guard21123 & _guard21124;
wire _guard21126 = fsm_out == 1'd0;
wire _guard21127 = cond_wire1002_out;
wire _guard21128 = _guard21126 & _guard21127;
wire _guard21129 = fsm_out == 1'd0;
wire _guard21130 = _guard21128 & _guard21129;
wire _guard21131 = fsm_out == 1'd0;
wire _guard21132 = cond_wire1004_out;
wire _guard21133 = _guard21131 & _guard21132;
wire _guard21134 = fsm_out == 1'd0;
wire _guard21135 = _guard21133 & _guard21134;
wire _guard21136 = _guard21130 | _guard21135;
wire _guard21137 = early_reset_static_par0_go_out;
wire _guard21138 = _guard21136 & _guard21137;
wire _guard21139 = fsm_out == 1'd0;
wire _guard21140 = cond_wire1002_out;
wire _guard21141 = _guard21139 & _guard21140;
wire _guard21142 = fsm_out == 1'd0;
wire _guard21143 = _guard21141 & _guard21142;
wire _guard21144 = fsm_out == 1'd0;
wire _guard21145 = cond_wire1004_out;
wire _guard21146 = _guard21144 & _guard21145;
wire _guard21147 = fsm_out == 1'd0;
wire _guard21148 = _guard21146 & _guard21147;
wire _guard21149 = _guard21143 | _guard21148;
wire _guard21150 = early_reset_static_par0_go_out;
wire _guard21151 = _guard21149 & _guard21150;
wire _guard21152 = fsm_out == 1'd0;
wire _guard21153 = cond_wire1002_out;
wire _guard21154 = _guard21152 & _guard21153;
wire _guard21155 = fsm_out == 1'd0;
wire _guard21156 = _guard21154 & _guard21155;
wire _guard21157 = fsm_out == 1'd0;
wire _guard21158 = cond_wire1004_out;
wire _guard21159 = _guard21157 & _guard21158;
wire _guard21160 = fsm_out == 1'd0;
wire _guard21161 = _guard21159 & _guard21160;
wire _guard21162 = _guard21156 | _guard21161;
wire _guard21163 = early_reset_static_par0_go_out;
wire _guard21164 = _guard21162 & _guard21163;
wire _guard21165 = cond_wire1016_out;
wire _guard21166 = early_reset_static_par0_go_out;
wire _guard21167 = _guard21165 & _guard21166;
wire _guard21168 = cond_wire1014_out;
wire _guard21169 = early_reset_static_par0_go_out;
wire _guard21170 = _guard21168 & _guard21169;
wire _guard21171 = fsm_out == 1'd0;
wire _guard21172 = cond_wire1014_out;
wire _guard21173 = _guard21171 & _guard21172;
wire _guard21174 = fsm_out == 1'd0;
wire _guard21175 = _guard21173 & _guard21174;
wire _guard21176 = fsm_out == 1'd0;
wire _guard21177 = cond_wire1016_out;
wire _guard21178 = _guard21176 & _guard21177;
wire _guard21179 = fsm_out == 1'd0;
wire _guard21180 = _guard21178 & _guard21179;
wire _guard21181 = _guard21175 | _guard21180;
wire _guard21182 = early_reset_static_par0_go_out;
wire _guard21183 = _guard21181 & _guard21182;
wire _guard21184 = fsm_out == 1'd0;
wire _guard21185 = cond_wire1014_out;
wire _guard21186 = _guard21184 & _guard21185;
wire _guard21187 = fsm_out == 1'd0;
wire _guard21188 = _guard21186 & _guard21187;
wire _guard21189 = fsm_out == 1'd0;
wire _guard21190 = cond_wire1016_out;
wire _guard21191 = _guard21189 & _guard21190;
wire _guard21192 = fsm_out == 1'd0;
wire _guard21193 = _guard21191 & _guard21192;
wire _guard21194 = _guard21188 | _guard21193;
wire _guard21195 = early_reset_static_par0_go_out;
wire _guard21196 = _guard21194 & _guard21195;
wire _guard21197 = fsm_out == 1'd0;
wire _guard21198 = cond_wire1014_out;
wire _guard21199 = _guard21197 & _guard21198;
wire _guard21200 = fsm_out == 1'd0;
wire _guard21201 = _guard21199 & _guard21200;
wire _guard21202 = fsm_out == 1'd0;
wire _guard21203 = cond_wire1016_out;
wire _guard21204 = _guard21202 & _guard21203;
wire _guard21205 = fsm_out == 1'd0;
wire _guard21206 = _guard21204 & _guard21205;
wire _guard21207 = _guard21201 | _guard21206;
wire _guard21208 = early_reset_static_par0_go_out;
wire _guard21209 = _guard21207 & _guard21208;
wire _guard21210 = cond_wire1051_out;
wire _guard21211 = early_reset_static_par0_go_out;
wire _guard21212 = _guard21210 & _guard21211;
wire _guard21213 = cond_wire1050_out;
wire _guard21214 = early_reset_static_par0_go_out;
wire _guard21215 = _guard21213 & _guard21214;
wire _guard21216 = fsm_out == 1'd0;
wire _guard21217 = cond_wire1050_out;
wire _guard21218 = _guard21216 & _guard21217;
wire _guard21219 = fsm_out == 1'd0;
wire _guard21220 = _guard21218 & _guard21219;
wire _guard21221 = fsm_out == 1'd0;
wire _guard21222 = cond_wire1051_out;
wire _guard21223 = _guard21221 & _guard21222;
wire _guard21224 = fsm_out == 1'd0;
wire _guard21225 = _guard21223 & _guard21224;
wire _guard21226 = _guard21220 | _guard21225;
wire _guard21227 = early_reset_static_par0_go_out;
wire _guard21228 = _guard21226 & _guard21227;
wire _guard21229 = fsm_out == 1'd0;
wire _guard21230 = cond_wire1050_out;
wire _guard21231 = _guard21229 & _guard21230;
wire _guard21232 = fsm_out == 1'd0;
wire _guard21233 = _guard21231 & _guard21232;
wire _guard21234 = fsm_out == 1'd0;
wire _guard21235 = cond_wire1051_out;
wire _guard21236 = _guard21234 & _guard21235;
wire _guard21237 = fsm_out == 1'd0;
wire _guard21238 = _guard21236 & _guard21237;
wire _guard21239 = _guard21233 | _guard21238;
wire _guard21240 = early_reset_static_par0_go_out;
wire _guard21241 = _guard21239 & _guard21240;
wire _guard21242 = fsm_out == 1'd0;
wire _guard21243 = cond_wire1050_out;
wire _guard21244 = _guard21242 & _guard21243;
wire _guard21245 = fsm_out == 1'd0;
wire _guard21246 = _guard21244 & _guard21245;
wire _guard21247 = fsm_out == 1'd0;
wire _guard21248 = cond_wire1051_out;
wire _guard21249 = _guard21247 & _guard21248;
wire _guard21250 = fsm_out == 1'd0;
wire _guard21251 = _guard21249 & _guard21250;
wire _guard21252 = _guard21246 | _guard21251;
wire _guard21253 = early_reset_static_par0_go_out;
wire _guard21254 = _guard21252 & _guard21253;
wire _guard21255 = cond_wire9_out;
wire _guard21256 = early_reset_static_par0_go_out;
wire _guard21257 = _guard21255 & _guard21256;
wire _guard21258 = cond_wire9_out;
wire _guard21259 = early_reset_static_par0_go_out;
wire _guard21260 = _guard21258 & _guard21259;
wire _guard21261 = cond_wire24_out;
wire _guard21262 = early_reset_static_par0_go_out;
wire _guard21263 = _guard21261 & _guard21262;
wire _guard21264 = cond_wire24_out;
wire _guard21265 = early_reset_static_par0_go_out;
wire _guard21266 = _guard21264 & _guard21265;
wire _guard21267 = cond_wire44_out;
wire _guard21268 = early_reset_static_par0_go_out;
wire _guard21269 = _guard21267 & _guard21268;
wire _guard21270 = cond_wire44_out;
wire _guard21271 = early_reset_static_par0_go_out;
wire _guard21272 = _guard21270 & _guard21271;
wire _guard21273 = fsm0_out == 6'd0;
wire _guard21274 = early_reset_static_seq_go_out;
wire _guard21275 = _guard21273 & _guard21274;
wire _guard21276 = cond_wire64_out;
wire _guard21277 = early_reset_static_par0_go_out;
wire _guard21278 = _guard21276 & _guard21277;
wire _guard21279 = _guard21275 | _guard21278;
wire _guard21280 = fsm0_out == 6'd0;
wire _guard21281 = early_reset_static_seq_go_out;
wire _guard21282 = _guard21280 & _guard21281;
wire _guard21283 = cond_wire64_out;
wire _guard21284 = early_reset_static_par0_go_out;
wire _guard21285 = _guard21283 & _guard21284;
wire _guard21286 = cond_wire534_out;
wire _guard21287 = early_reset_static_par0_go_out;
wire _guard21288 = _guard21286 & _guard21287;
wire _guard21289 = cond_wire534_out;
wire _guard21290 = early_reset_static_par0_go_out;
wire _guard21291 = _guard21289 & _guard21290;
wire _guard21292 = early_reset_static_par0_go_out;
wire _guard21293 = early_reset_static_par0_go_out;
wire _guard21294 = early_reset_static_par0_go_out;
wire _guard21295 = early_reset_static_par0_go_out;
wire _guard21296 = early_reset_static_par0_go_out;
wire _guard21297 = early_reset_static_par0_go_out;
wire _guard21298 = early_reset_static_par0_go_out;
wire _guard21299 = early_reset_static_par0_go_out;
wire _guard21300 = early_reset_static_par0_go_out;
wire _guard21301 = early_reset_static_par0_go_out;
wire _guard21302 = fsm0_out == 6'd0;
wire _guard21303 = early_reset_static_seq_go_out;
wire _guard21304 = _guard21302 & _guard21303;
wire _guard21305 = early_reset_static_par0_go_out;
wire _guard21306 = _guard21304 | _guard21305;
wire _guard21307 = fsm0_out == 6'd0;
wire _guard21308 = early_reset_static_seq_go_out;
wire _guard21309 = _guard21307 & _guard21308;
wire _guard21310 = early_reset_static_par0_go_out;
wire _guard21311 = early_reset_static_par0_go_out;
wire _guard21312 = early_reset_static_par0_go_out;
wire _guard21313 = early_reset_static_par0_go_out;
wire _guard21314 = early_reset_static_par0_go_out;
wire _guard21315 = fsm0_out == 6'd0;
wire _guard21316 = early_reset_static_seq_go_out;
wire _guard21317 = _guard21315 & _guard21316;
wire _guard21318 = early_reset_static_par0_go_out;
wire _guard21319 = _guard21317 | _guard21318;
wire _guard21320 = early_reset_static_par0_go_out;
wire _guard21321 = fsm0_out == 6'd0;
wire _guard21322 = early_reset_static_seq_go_out;
wire _guard21323 = _guard21321 & _guard21322;
wire _guard21324 = fsm0_out == 6'd0;
wire _guard21325 = early_reset_static_seq_go_out;
wire _guard21326 = _guard21324 & _guard21325;
wire _guard21327 = early_reset_static_par0_go_out;
wire _guard21328 = _guard21326 | _guard21327;
wire _guard21329 = early_reset_static_par0_go_out;
wire _guard21330 = fsm0_out == 6'd0;
wire _guard21331 = early_reset_static_seq_go_out;
wire _guard21332 = _guard21330 & _guard21331;
wire _guard21333 = early_reset_static_par0_go_out;
wire _guard21334 = early_reset_static_par0_go_out;
wire _guard21335 = early_reset_static_par0_go_out;
wire _guard21336 = early_reset_static_par0_go_out;
wire _guard21337 = early_reset_static_par0_go_out;
wire _guard21338 = early_reset_static_par0_go_out;
wire _guard21339 = early_reset_static_par0_go_out;
wire _guard21340 = early_reset_static_par0_go_out;
wire _guard21341 = fsm0_out == 6'd0;
wire _guard21342 = early_reset_static_seq_go_out;
wire _guard21343 = _guard21341 & _guard21342;
wire _guard21344 = early_reset_static_par0_go_out;
wire _guard21345 = _guard21343 | _guard21344;
wire _guard21346 = early_reset_static_par0_go_out;
wire _guard21347 = fsm0_out == 6'd0;
wire _guard21348 = early_reset_static_seq_go_out;
wire _guard21349 = _guard21347 & _guard21348;
wire _guard21350 = early_reset_static_par0_go_out;
wire _guard21351 = early_reset_static_par0_go_out;
wire _guard21352 = fsm0_out == 6'd0;
wire _guard21353 = early_reset_static_seq_go_out;
wire _guard21354 = _guard21352 & _guard21353;
wire _guard21355 = early_reset_static_par0_go_out;
wire _guard21356 = _guard21354 | _guard21355;
wire _guard21357 = early_reset_static_par0_go_out;
wire _guard21358 = fsm0_out == 6'd0;
wire _guard21359 = early_reset_static_seq_go_out;
wire _guard21360 = _guard21358 & _guard21359;
wire _guard21361 = early_reset_static_par0_go_out;
wire _guard21362 = early_reset_static_par0_go_out;
wire _guard21363 = fsm0_out == 6'd0;
wire _guard21364 = early_reset_static_seq_go_out;
wire _guard21365 = _guard21363 & _guard21364;
wire _guard21366 = early_reset_static_par0_go_out;
wire _guard21367 = _guard21365 | _guard21366;
wire _guard21368 = early_reset_static_par0_go_out;
wire _guard21369 = fsm0_out == 6'd0;
wire _guard21370 = early_reset_static_seq_go_out;
wire _guard21371 = _guard21369 & _guard21370;
wire _guard21372 = fsm0_out == 6'd0;
wire _guard21373 = early_reset_static_seq_go_out;
wire _guard21374 = _guard21372 & _guard21373;
wire _guard21375 = early_reset_static_par0_go_out;
wire _guard21376 = _guard21374 | _guard21375;
wire _guard21377 = early_reset_static_par0_go_out;
wire _guard21378 = fsm0_out == 6'd0;
wire _guard21379 = early_reset_static_seq_go_out;
wire _guard21380 = _guard21378 & _guard21379;
wire _guard21381 = fsm0_out == 6'd0;
wire _guard21382 = early_reset_static_seq_go_out;
wire _guard21383 = _guard21381 & _guard21382;
wire _guard21384 = early_reset_static_par0_go_out;
wire _guard21385 = _guard21383 | _guard21384;
wire _guard21386 = fsm0_out == 6'd0;
wire _guard21387 = early_reset_static_seq_go_out;
wire _guard21388 = _guard21386 & _guard21387;
wire _guard21389 = early_reset_static_par0_go_out;
wire _guard21390 = early_reset_static_par0_go_out;
wire _guard21391 = early_reset_static_par0_go_out;
wire _guard21392 = early_reset_static_par0_go_out;
wire _guard21393 = ~_guard0;
wire _guard21394 = early_reset_static_par0_go_out;
wire _guard21395 = _guard21393 & _guard21394;
wire _guard21396 = early_reset_static_par0_go_out;
wire _guard21397 = ~_guard0;
wire _guard21398 = early_reset_static_par0_go_out;
wire _guard21399 = _guard21397 & _guard21398;
wire _guard21400 = early_reset_static_par0_go_out;
wire _guard21401 = ~_guard0;
wire _guard21402 = early_reset_static_par0_go_out;
wire _guard21403 = _guard21401 & _guard21402;
wire _guard21404 = ~_guard0;
wire _guard21405 = early_reset_static_par0_go_out;
wire _guard21406 = _guard21404 & _guard21405;
wire _guard21407 = early_reset_static_par0_go_out;
wire _guard21408 = ~_guard0;
wire _guard21409 = early_reset_static_par0_go_out;
wire _guard21410 = _guard21408 & _guard21409;
wire _guard21411 = early_reset_static_par0_go_out;
wire _guard21412 = early_reset_static_par0_go_out;
wire _guard21413 = ~_guard0;
wire _guard21414 = early_reset_static_par0_go_out;
wire _guard21415 = _guard21413 & _guard21414;
wire _guard21416 = early_reset_static_par0_go_out;
wire _guard21417 = ~_guard0;
wire _guard21418 = early_reset_static_par0_go_out;
wire _guard21419 = _guard21417 & _guard21418;
wire _guard21420 = early_reset_static_par0_go_out;
wire _guard21421 = early_reset_static_par0_go_out;
wire _guard21422 = early_reset_static_par0_go_out;
wire _guard21423 = ~_guard0;
wire _guard21424 = early_reset_static_par0_go_out;
wire _guard21425 = _guard21423 & _guard21424;
wire _guard21426 = early_reset_static_par0_go_out;
wire _guard21427 = early_reset_static_par0_go_out;
wire _guard21428 = early_reset_static_par0_go_out;
wire _guard21429 = early_reset_static_par0_go_out;
wire _guard21430 = early_reset_static_par0_go_out;
wire _guard21431 = early_reset_static_par0_go_out;
wire _guard21432 = ~_guard0;
wire _guard21433 = early_reset_static_par0_go_out;
wire _guard21434 = _guard21432 & _guard21433;
wire _guard21435 = early_reset_static_par0_go_out;
wire _guard21436 = ~_guard0;
wire _guard21437 = early_reset_static_par0_go_out;
wire _guard21438 = _guard21436 & _guard21437;
wire _guard21439 = early_reset_static_par0_go_out;
wire _guard21440 = early_reset_static_par0_go_out;
wire _guard21441 = early_reset_static_par0_go_out;
wire _guard21442 = early_reset_static_par0_go_out;
wire _guard21443 = early_reset_static_par0_go_out;
wire _guard21444 = ~_guard0;
wire _guard21445 = early_reset_static_par0_go_out;
wire _guard21446 = _guard21444 & _guard21445;
wire _guard21447 = early_reset_static_par0_go_out;
wire _guard21448 = early_reset_static_par0_go_out;
wire _guard21449 = early_reset_static_par0_go_out;
wire _guard21450 = early_reset_static_par0_go_out;
wire _guard21451 = ~_guard0;
wire _guard21452 = early_reset_static_par0_go_out;
wire _guard21453 = _guard21451 & _guard21452;
wire _guard21454 = early_reset_static_par0_go_out;
wire _guard21455 = early_reset_static_par0_go_out;
wire _guard21456 = early_reset_static_par0_go_out;
wire _guard21457 = ~_guard0;
wire _guard21458 = early_reset_static_par0_go_out;
wire _guard21459 = _guard21457 & _guard21458;
wire _guard21460 = early_reset_static_par0_go_out;
wire _guard21461 = early_reset_static_par0_go_out;
wire _guard21462 = early_reset_static_par0_go_out;
wire _guard21463 = early_reset_static_par0_go_out;
wire _guard21464 = early_reset_static_par0_go_out;
wire _guard21465 = ~_guard0;
wire _guard21466 = early_reset_static_par0_go_out;
wire _guard21467 = _guard21465 & _guard21466;
wire _guard21468 = early_reset_static_par0_go_out;
wire _guard21469 = ~_guard0;
wire _guard21470 = early_reset_static_par0_go_out;
wire _guard21471 = _guard21469 & _guard21470;
wire _guard21472 = early_reset_static_par0_go_out;
wire _guard21473 = early_reset_static_par0_go_out;
wire _guard21474 = ~_guard0;
wire _guard21475 = early_reset_static_par0_go_out;
wire _guard21476 = _guard21474 & _guard21475;
wire _guard21477 = early_reset_static_par0_go_out;
wire _guard21478 = early_reset_static_par0_go_out;
wire _guard21479 = ~_guard0;
wire _guard21480 = early_reset_static_par0_go_out;
wire _guard21481 = _guard21479 & _guard21480;
wire _guard21482 = early_reset_static_par0_go_out;
wire _guard21483 = ~_guard0;
wire _guard21484 = early_reset_static_par0_go_out;
wire _guard21485 = _guard21483 & _guard21484;
wire _guard21486 = early_reset_static_par0_go_out;
wire _guard21487 = early_reset_static_par0_go_out;
wire _guard21488 = early_reset_static_par0_go_out;
wire _guard21489 = early_reset_static_par0_go_out;
wire _guard21490 = early_reset_static_par0_go_out;
wire _guard21491 = early_reset_static_par0_go_out;
wire _guard21492 = ~_guard0;
wire _guard21493 = early_reset_static_par0_go_out;
wire _guard21494 = _guard21492 & _guard21493;
wire _guard21495 = early_reset_static_par0_go_out;
wire _guard21496 = ~_guard0;
wire _guard21497 = early_reset_static_par0_go_out;
wire _guard21498 = _guard21496 & _guard21497;
wire _guard21499 = early_reset_static_par0_go_out;
wire _guard21500 = early_reset_static_par0_go_out;
wire _guard21501 = ~_guard0;
wire _guard21502 = early_reset_static_par0_go_out;
wire _guard21503 = _guard21501 & _guard21502;
wire _guard21504 = early_reset_static_par0_go_out;
wire _guard21505 = ~_guard0;
wire _guard21506 = early_reset_static_par0_go_out;
wire _guard21507 = _guard21505 & _guard21506;
wire _guard21508 = early_reset_static_par0_go_out;
wire _guard21509 = early_reset_static_par0_go_out;
wire _guard21510 = early_reset_static_par0_go_out;
wire _guard21511 = early_reset_static_par0_go_out;
wire _guard21512 = early_reset_static_par0_go_out;
wire _guard21513 = ~_guard0;
wire _guard21514 = early_reset_static_par0_go_out;
wire _guard21515 = _guard21513 & _guard21514;
wire _guard21516 = early_reset_static_par0_go_out;
wire _guard21517 = ~_guard0;
wire _guard21518 = early_reset_static_par0_go_out;
wire _guard21519 = _guard21517 & _guard21518;
wire _guard21520 = early_reset_static_par0_go_out;
wire _guard21521 = ~_guard0;
wire _guard21522 = early_reset_static_par0_go_out;
wire _guard21523 = _guard21521 & _guard21522;
wire _guard21524 = early_reset_static_par0_go_out;
wire _guard21525 = early_reset_static_par0_go_out;
wire _guard21526 = early_reset_static_par0_go_out;
wire _guard21527 = ~_guard0;
wire _guard21528 = early_reset_static_par0_go_out;
wire _guard21529 = _guard21527 & _guard21528;
wire _guard21530 = early_reset_static_par0_go_out;
wire _guard21531 = early_reset_static_par0_go_out;
wire _guard21532 = early_reset_static_par0_go_out;
wire _guard21533 = early_reset_static_par0_go_out;
wire _guard21534 = ~_guard0;
wire _guard21535 = early_reset_static_par0_go_out;
wire _guard21536 = _guard21534 & _guard21535;
wire _guard21537 = early_reset_static_par0_go_out;
wire _guard21538 = early_reset_static_par0_go_out;
wire _guard21539 = ~_guard0;
wire _guard21540 = early_reset_static_par0_go_out;
wire _guard21541 = _guard21539 & _guard21540;
wire _guard21542 = early_reset_static_par0_go_out;
wire _guard21543 = ~_guard0;
wire _guard21544 = early_reset_static_par0_go_out;
wire _guard21545 = _guard21543 & _guard21544;
wire _guard21546 = early_reset_static_par0_go_out;
wire _guard21547 = ~_guard0;
wire _guard21548 = early_reset_static_par0_go_out;
wire _guard21549 = _guard21547 & _guard21548;
wire _guard21550 = early_reset_static_par0_go_out;
wire _guard21551 = early_reset_static_par0_go_out;
wire _guard21552 = ~_guard0;
wire _guard21553 = early_reset_static_par0_go_out;
wire _guard21554 = _guard21552 & _guard21553;
wire _guard21555 = early_reset_static_par0_go_out;
wire _guard21556 = ~_guard0;
wire _guard21557 = early_reset_static_par0_go_out;
wire _guard21558 = _guard21556 & _guard21557;
wire _guard21559 = early_reset_static_par0_go_out;
wire _guard21560 = ~_guard0;
wire _guard21561 = early_reset_static_par0_go_out;
wire _guard21562 = _guard21560 & _guard21561;
wire _guard21563 = early_reset_static_par0_go_out;
wire _guard21564 = early_reset_static_par0_go_out;
wire _guard21565 = ~_guard0;
wire _guard21566 = early_reset_static_par0_go_out;
wire _guard21567 = _guard21565 & _guard21566;
wire _guard21568 = early_reset_static_par0_go_out;
wire _guard21569 = early_reset_static_par0_go_out;
wire _guard21570 = early_reset_static_par0_go_out;
wire _guard21571 = ~_guard0;
wire _guard21572 = early_reset_static_par0_go_out;
wire _guard21573 = _guard21571 & _guard21572;
wire _guard21574 = early_reset_static_par0_go_out;
wire _guard21575 = early_reset_static_par0_go_out;
wire _guard21576 = early_reset_static_par0_go_out;
wire _guard21577 = early_reset_static_par0_go_out;
wire _guard21578 = early_reset_static_par0_go_out;
wire _guard21579 = early_reset_static_par0_go_out;
wire _guard21580 = early_reset_static_par0_go_out;
wire _guard21581 = early_reset_static_par0_go_out;
wire _guard21582 = early_reset_static_par0_go_out;
wire _guard21583 = early_reset_static_par0_go_out;
wire _guard21584 = early_reset_static_par0_go_out;
wire _guard21585 = early_reset_static_par0_go_out;
wire _guard21586 = ~_guard0;
wire _guard21587 = early_reset_static_par0_go_out;
wire _guard21588 = _guard21586 & _guard21587;
wire _guard21589 = early_reset_static_par0_go_out;
wire _guard21590 = early_reset_static_par0_go_out;
wire _guard21591 = early_reset_static_par0_go_out;
wire _guard21592 = early_reset_static_par0_go_out;
wire _guard21593 = ~_guard0;
wire _guard21594 = early_reset_static_par0_go_out;
wire _guard21595 = _guard21593 & _guard21594;
wire _guard21596 = early_reset_static_par0_go_out;
wire _guard21597 = early_reset_static_par0_go_out;
wire _guard21598 = early_reset_static_par0_go_out;
wire _guard21599 = early_reset_static_par0_go_out;
wire _guard21600 = ~_guard0;
wire _guard21601 = early_reset_static_par0_go_out;
wire _guard21602 = _guard21600 & _guard21601;
wire _guard21603 = early_reset_static_par0_go_out;
wire _guard21604 = early_reset_static_par0_go_out;
wire _guard21605 = ~_guard0;
wire _guard21606 = early_reset_static_par0_go_out;
wire _guard21607 = _guard21605 & _guard21606;
wire _guard21608 = early_reset_static_par0_go_out;
wire _guard21609 = early_reset_static_par0_go_out;
wire _guard21610 = early_reset_static_par0_go_out;
wire _guard21611 = ~_guard0;
wire _guard21612 = early_reset_static_par0_go_out;
wire _guard21613 = _guard21611 & _guard21612;
wire _guard21614 = ~_guard0;
wire _guard21615 = early_reset_static_par0_go_out;
wire _guard21616 = _guard21614 & _guard21615;
wire _guard21617 = early_reset_static_par0_go_out;
wire _guard21618 = early_reset_static_par0_go_out;
wire _guard21619 = early_reset_static_par0_go_out;
wire _guard21620 = early_reset_static_par0_go_out;
wire _guard21621 = early_reset_static_par0_go_out;
wire _guard21622 = ~_guard0;
wire _guard21623 = early_reset_static_par0_go_out;
wire _guard21624 = _guard21622 & _guard21623;
wire _guard21625 = early_reset_static_par0_go_out;
wire _guard21626 = early_reset_static_par0_go_out;
wire _guard21627 = ~_guard0;
wire _guard21628 = early_reset_static_par0_go_out;
wire _guard21629 = _guard21627 & _guard21628;
wire _guard21630 = early_reset_static_par0_go_out;
wire _guard21631 = early_reset_static_par0_go_out;
wire _guard21632 = ~_guard0;
wire _guard21633 = early_reset_static_par0_go_out;
wire _guard21634 = _guard21632 & _guard21633;
wire _guard21635 = early_reset_static_par0_go_out;
wire _guard21636 = early_reset_static_par0_go_out;
wire _guard21637 = early_reset_static_par0_go_out;
wire _guard21638 = early_reset_static_par0_go_out;
wire _guard21639 = early_reset_static_par0_go_out;
wire _guard21640 = early_reset_static_par0_go_out;
wire _guard21641 = ~_guard0;
wire _guard21642 = early_reset_static_par0_go_out;
wire _guard21643 = _guard21641 & _guard21642;
wire _guard21644 = early_reset_static_par0_go_out;
wire _guard21645 = early_reset_static_par0_go_out;
wire _guard21646 = early_reset_static_par0_go_out;
wire _guard21647 = early_reset_static_par0_go_out;
wire _guard21648 = ~_guard0;
wire _guard21649 = early_reset_static_par0_go_out;
wire _guard21650 = _guard21648 & _guard21649;
wire _guard21651 = early_reset_static_par0_go_out;
wire _guard21652 = ~_guard0;
wire _guard21653 = early_reset_static_par0_go_out;
wire _guard21654 = _guard21652 & _guard21653;
wire _guard21655 = early_reset_static_par0_go_out;
wire _guard21656 = early_reset_static_par0_go_out;
wire _guard21657 = early_reset_static_par0_go_out;
wire _guard21658 = early_reset_static_par0_go_out;
wire _guard21659 = ~_guard0;
wire _guard21660 = early_reset_static_par0_go_out;
wire _guard21661 = _guard21659 & _guard21660;
wire _guard21662 = ~_guard0;
wire _guard21663 = early_reset_static_par0_go_out;
wire _guard21664 = _guard21662 & _guard21663;
wire _guard21665 = early_reset_static_par0_go_out;
wire _guard21666 = early_reset_static_par0_go_out;
wire _guard21667 = early_reset_static_par0_go_out;
wire _guard21668 = early_reset_static_par0_go_out;
wire _guard21669 = ~_guard0;
wire _guard21670 = early_reset_static_par0_go_out;
wire _guard21671 = _guard21669 & _guard21670;
wire _guard21672 = early_reset_static_par0_go_out;
wire _guard21673 = early_reset_static_par0_go_out;
wire _guard21674 = early_reset_static_par0_go_out;
wire _guard21675 = early_reset_static_par0_go_out;
wire _guard21676 = early_reset_static_par0_go_out;
wire _guard21677 = early_reset_static_par0_go_out;
wire _guard21678 = early_reset_static_par0_go_out;
wire _guard21679 = ~_guard0;
wire _guard21680 = early_reset_static_par0_go_out;
wire _guard21681 = _guard21679 & _guard21680;
wire _guard21682 = early_reset_static_par0_go_out;
wire _guard21683 = early_reset_static_par0_go_out;
wire _guard21684 = early_reset_static_par0_go_out;
wire _guard21685 = early_reset_static_par0_go_out;
wire _guard21686 = ~_guard0;
wire _guard21687 = early_reset_static_par0_go_out;
wire _guard21688 = _guard21686 & _guard21687;
wire _guard21689 = early_reset_static_par0_go_out;
wire _guard21690 = ~_guard0;
wire _guard21691 = early_reset_static_par0_go_out;
wire _guard21692 = _guard21690 & _guard21691;
wire _guard21693 = early_reset_static_par0_go_out;
wire _guard21694 = early_reset_static_par0_go_out;
wire _guard21695 = early_reset_static_par0_go_out;
wire _guard21696 = early_reset_static_par0_go_out;
wire _guard21697 = ~_guard0;
wire _guard21698 = early_reset_static_par0_go_out;
wire _guard21699 = _guard21697 & _guard21698;
wire _guard21700 = early_reset_static_par0_go_out;
wire _guard21701 = ~_guard0;
wire _guard21702 = early_reset_static_par0_go_out;
wire _guard21703 = _guard21701 & _guard21702;
wire _guard21704 = early_reset_static_par0_go_out;
wire _guard21705 = ~_guard0;
wire _guard21706 = early_reset_static_par0_go_out;
wire _guard21707 = _guard21705 & _guard21706;
wire _guard21708 = early_reset_static_par0_go_out;
wire _guard21709 = early_reset_static_par0_go_out;
wire _guard21710 = ~_guard0;
wire _guard21711 = early_reset_static_par0_go_out;
wire _guard21712 = _guard21710 & _guard21711;
wire _guard21713 = early_reset_static_par0_go_out;
wire _guard21714 = early_reset_static_par0_go_out;
wire _guard21715 = early_reset_static_par0_go_out;
wire _guard21716 = early_reset_static_par0_go_out;
wire _guard21717 = early_reset_static_par0_go_out;
wire _guard21718 = early_reset_static_par0_go_out;
wire _guard21719 = early_reset_static_par0_go_out;
wire _guard21720 = ~_guard0;
wire _guard21721 = early_reset_static_par0_go_out;
wire _guard21722 = _guard21720 & _guard21721;
wire _guard21723 = early_reset_static_par0_go_out;
wire _guard21724 = ~_guard0;
wire _guard21725 = early_reset_static_par0_go_out;
wire _guard21726 = _guard21724 & _guard21725;
wire _guard21727 = early_reset_static_par0_go_out;
wire _guard21728 = ~_guard0;
wire _guard21729 = early_reset_static_par0_go_out;
wire _guard21730 = _guard21728 & _guard21729;
wire _guard21731 = early_reset_static_par0_go_out;
wire _guard21732 = ~_guard0;
wire _guard21733 = early_reset_static_par0_go_out;
wire _guard21734 = _guard21732 & _guard21733;
wire _guard21735 = early_reset_static_par0_go_out;
wire _guard21736 = ~_guard0;
wire _guard21737 = early_reset_static_par0_go_out;
wire _guard21738 = _guard21736 & _guard21737;
wire _guard21739 = early_reset_static_par0_go_out;
wire _guard21740 = ~_guard0;
wire _guard21741 = early_reset_static_par0_go_out;
wire _guard21742 = _guard21740 & _guard21741;
wire _guard21743 = early_reset_static_par0_go_out;
wire _guard21744 = ~_guard0;
wire _guard21745 = early_reset_static_par0_go_out;
wire _guard21746 = _guard21744 & _guard21745;
wire _guard21747 = early_reset_static_par0_go_out;
wire _guard21748 = early_reset_static_par0_go_out;
wire _guard21749 = ~_guard0;
wire _guard21750 = early_reset_static_par0_go_out;
wire _guard21751 = _guard21749 & _guard21750;
wire _guard21752 = early_reset_static_par0_go_out;
wire _guard21753 = ~_guard0;
wire _guard21754 = early_reset_static_par0_go_out;
wire _guard21755 = _guard21753 & _guard21754;
wire _guard21756 = early_reset_static_par0_go_out;
wire _guard21757 = ~_guard0;
wire _guard21758 = early_reset_static_par0_go_out;
wire _guard21759 = _guard21757 & _guard21758;
wire _guard21760 = early_reset_static_par0_go_out;
wire _guard21761 = early_reset_static_par0_go_out;
wire _guard21762 = ~_guard0;
wire _guard21763 = early_reset_static_par0_go_out;
wire _guard21764 = _guard21762 & _guard21763;
wire _guard21765 = early_reset_static_par0_go_out;
wire _guard21766 = ~_guard0;
wire _guard21767 = early_reset_static_par0_go_out;
wire _guard21768 = _guard21766 & _guard21767;
wire _guard21769 = early_reset_static_par0_go_out;
wire _guard21770 = early_reset_static_par0_go_out;
wire _guard21771 = early_reset_static_par0_go_out;
wire _guard21772 = ~_guard0;
wire _guard21773 = early_reset_static_par0_go_out;
wire _guard21774 = _guard21772 & _guard21773;
wire _guard21775 = early_reset_static_par0_go_out;
wire _guard21776 = early_reset_static_par0_go_out;
wire _guard21777 = early_reset_static_par0_go_out;
wire _guard21778 = early_reset_static_par0_go_out;
wire _guard21779 = ~_guard0;
wire _guard21780 = early_reset_static_par0_go_out;
wire _guard21781 = _guard21779 & _guard21780;
wire _guard21782 = early_reset_static_par0_go_out;
wire _guard21783 = early_reset_static_par0_go_out;
wire _guard21784 = early_reset_static_par0_go_out;
wire _guard21785 = early_reset_static_par0_go_out;
wire _guard21786 = cond_wire14_out;
wire _guard21787 = early_reset_static_par0_go_out;
wire _guard21788 = _guard21786 & _guard21787;
wire _guard21789 = cond_wire14_out;
wire _guard21790 = early_reset_static_par0_go_out;
wire _guard21791 = _guard21789 & _guard21790;
wire _guard21792 = cond_wire32_out;
wire _guard21793 = early_reset_static_par0_go_out;
wire _guard21794 = _guard21792 & _guard21793;
wire _guard21795 = cond_wire30_out;
wire _guard21796 = early_reset_static_par0_go_out;
wire _guard21797 = _guard21795 & _guard21796;
wire _guard21798 = fsm_out == 1'd0;
wire _guard21799 = cond_wire30_out;
wire _guard21800 = _guard21798 & _guard21799;
wire _guard21801 = fsm_out == 1'd0;
wire _guard21802 = _guard21800 & _guard21801;
wire _guard21803 = fsm_out == 1'd0;
wire _guard21804 = cond_wire32_out;
wire _guard21805 = _guard21803 & _guard21804;
wire _guard21806 = fsm_out == 1'd0;
wire _guard21807 = _guard21805 & _guard21806;
wire _guard21808 = _guard21802 | _guard21807;
wire _guard21809 = early_reset_static_par0_go_out;
wire _guard21810 = _guard21808 & _guard21809;
wire _guard21811 = fsm_out == 1'd0;
wire _guard21812 = cond_wire30_out;
wire _guard21813 = _guard21811 & _guard21812;
wire _guard21814 = fsm_out == 1'd0;
wire _guard21815 = _guard21813 & _guard21814;
wire _guard21816 = fsm_out == 1'd0;
wire _guard21817 = cond_wire32_out;
wire _guard21818 = _guard21816 & _guard21817;
wire _guard21819 = fsm_out == 1'd0;
wire _guard21820 = _guard21818 & _guard21819;
wire _guard21821 = _guard21815 | _guard21820;
wire _guard21822 = early_reset_static_par0_go_out;
wire _guard21823 = _guard21821 & _guard21822;
wire _guard21824 = fsm_out == 1'd0;
wire _guard21825 = cond_wire30_out;
wire _guard21826 = _guard21824 & _guard21825;
wire _guard21827 = fsm_out == 1'd0;
wire _guard21828 = _guard21826 & _guard21827;
wire _guard21829 = fsm_out == 1'd0;
wire _guard21830 = cond_wire32_out;
wire _guard21831 = _guard21829 & _guard21830;
wire _guard21832 = fsm_out == 1'd0;
wire _guard21833 = _guard21831 & _guard21832;
wire _guard21834 = _guard21828 | _guard21833;
wire _guard21835 = early_reset_static_par0_go_out;
wire _guard21836 = _guard21834 & _guard21835;
wire _guard21837 = cond_wire36_out;
wire _guard21838 = early_reset_static_par0_go_out;
wire _guard21839 = _guard21837 & _guard21838;
wire _guard21840 = cond_wire36_out;
wire _guard21841 = early_reset_static_par0_go_out;
wire _guard21842 = _guard21840 & _guard21841;
wire _guard21843 = cond_wire61_out;
wire _guard21844 = early_reset_static_par0_go_out;
wire _guard21845 = _guard21843 & _guard21844;
wire _guard21846 = cond_wire61_out;
wire _guard21847 = early_reset_static_par0_go_out;
wire _guard21848 = _guard21846 & _guard21847;
wire _guard21849 = cond_wire137_out;
wire _guard21850 = early_reset_static_par0_go_out;
wire _guard21851 = _guard21849 & _guard21850;
wire _guard21852 = cond_wire137_out;
wire _guard21853 = early_reset_static_par0_go_out;
wire _guard21854 = _guard21852 & _guard21853;
wire _guard21855 = cond_wire85_out;
wire _guard21856 = early_reset_static_par0_go_out;
wire _guard21857 = _guard21855 & _guard21856;
wire _guard21858 = cond_wire85_out;
wire _guard21859 = early_reset_static_par0_go_out;
wire _guard21860 = _guard21858 & _guard21859;
wire _guard21861 = cond_wire121_out;
wire _guard21862 = early_reset_static_par0_go_out;
wire _guard21863 = _guard21861 & _guard21862;
wire _guard21864 = cond_wire121_out;
wire _guard21865 = early_reset_static_par0_go_out;
wire _guard21866 = _guard21864 & _guard21865;
wire _guard21867 = cond_wire219_out;
wire _guard21868 = early_reset_static_par0_go_out;
wire _guard21869 = _guard21867 & _guard21868;
wire _guard21870 = cond_wire219_out;
wire _guard21871 = early_reset_static_par0_go_out;
wire _guard21872 = _guard21870 & _guard21871;
wire _guard21873 = cond_wire174_out;
wire _guard21874 = early_reset_static_par0_go_out;
wire _guard21875 = _guard21873 & _guard21874;
wire _guard21876 = cond_wire174_out;
wire _guard21877 = early_reset_static_par0_go_out;
wire _guard21878 = _guard21876 & _guard21877;
wire _guard21879 = cond_wire198_out;
wire _guard21880 = early_reset_static_par0_go_out;
wire _guard21881 = _guard21879 & _guard21880;
wire _guard21882 = cond_wire198_out;
wire _guard21883 = early_reset_static_par0_go_out;
wire _guard21884 = _guard21882 & _guard21883;
wire _guard21885 = cond_wire276_out;
wire _guard21886 = early_reset_static_par0_go_out;
wire _guard21887 = _guard21885 & _guard21886;
wire _guard21888 = cond_wire276_out;
wire _guard21889 = early_reset_static_par0_go_out;
wire _guard21890 = _guard21888 & _guard21889;
wire _guard21891 = cond_wire289_out;
wire _guard21892 = early_reset_static_par0_go_out;
wire _guard21893 = _guard21891 & _guard21892;
wire _guard21894 = cond_wire287_out;
wire _guard21895 = early_reset_static_par0_go_out;
wire _guard21896 = _guard21894 & _guard21895;
wire _guard21897 = fsm_out == 1'd0;
wire _guard21898 = cond_wire287_out;
wire _guard21899 = _guard21897 & _guard21898;
wire _guard21900 = fsm_out == 1'd0;
wire _guard21901 = _guard21899 & _guard21900;
wire _guard21902 = fsm_out == 1'd0;
wire _guard21903 = cond_wire289_out;
wire _guard21904 = _guard21902 & _guard21903;
wire _guard21905 = fsm_out == 1'd0;
wire _guard21906 = _guard21904 & _guard21905;
wire _guard21907 = _guard21901 | _guard21906;
wire _guard21908 = early_reset_static_par0_go_out;
wire _guard21909 = _guard21907 & _guard21908;
wire _guard21910 = fsm_out == 1'd0;
wire _guard21911 = cond_wire287_out;
wire _guard21912 = _guard21910 & _guard21911;
wire _guard21913 = fsm_out == 1'd0;
wire _guard21914 = _guard21912 & _guard21913;
wire _guard21915 = fsm_out == 1'd0;
wire _guard21916 = cond_wire289_out;
wire _guard21917 = _guard21915 & _guard21916;
wire _guard21918 = fsm_out == 1'd0;
wire _guard21919 = _guard21917 & _guard21918;
wire _guard21920 = _guard21914 | _guard21919;
wire _guard21921 = early_reset_static_par0_go_out;
wire _guard21922 = _guard21920 & _guard21921;
wire _guard21923 = fsm_out == 1'd0;
wire _guard21924 = cond_wire287_out;
wire _guard21925 = _guard21923 & _guard21924;
wire _guard21926 = fsm_out == 1'd0;
wire _guard21927 = _guard21925 & _guard21926;
wire _guard21928 = fsm_out == 1'd0;
wire _guard21929 = cond_wire289_out;
wire _guard21930 = _guard21928 & _guard21929;
wire _guard21931 = fsm_out == 1'd0;
wire _guard21932 = _guard21930 & _guard21931;
wire _guard21933 = _guard21927 | _guard21932;
wire _guard21934 = early_reset_static_par0_go_out;
wire _guard21935 = _guard21933 & _guard21934;
wire _guard21936 = cond_wire243_out;
wire _guard21937 = early_reset_static_par0_go_out;
wire _guard21938 = _guard21936 & _guard21937;
wire _guard21939 = cond_wire243_out;
wire _guard21940 = early_reset_static_par0_go_out;
wire _guard21941 = _guard21939 & _guard21940;
wire _guard21942 = cond_wire317_out;
wire _guard21943 = early_reset_static_par0_go_out;
wire _guard21944 = _guard21942 & _guard21943;
wire _guard21945 = cond_wire315_out;
wire _guard21946 = early_reset_static_par0_go_out;
wire _guard21947 = _guard21945 & _guard21946;
wire _guard21948 = fsm_out == 1'd0;
wire _guard21949 = cond_wire315_out;
wire _guard21950 = _guard21948 & _guard21949;
wire _guard21951 = fsm_out == 1'd0;
wire _guard21952 = _guard21950 & _guard21951;
wire _guard21953 = fsm_out == 1'd0;
wire _guard21954 = cond_wire317_out;
wire _guard21955 = _guard21953 & _guard21954;
wire _guard21956 = fsm_out == 1'd0;
wire _guard21957 = _guard21955 & _guard21956;
wire _guard21958 = _guard21952 | _guard21957;
wire _guard21959 = early_reset_static_par0_go_out;
wire _guard21960 = _guard21958 & _guard21959;
wire _guard21961 = fsm_out == 1'd0;
wire _guard21962 = cond_wire315_out;
wire _guard21963 = _guard21961 & _guard21962;
wire _guard21964 = fsm_out == 1'd0;
wire _guard21965 = _guard21963 & _guard21964;
wire _guard21966 = fsm_out == 1'd0;
wire _guard21967 = cond_wire317_out;
wire _guard21968 = _guard21966 & _guard21967;
wire _guard21969 = fsm_out == 1'd0;
wire _guard21970 = _guard21968 & _guard21969;
wire _guard21971 = _guard21965 | _guard21970;
wire _guard21972 = early_reset_static_par0_go_out;
wire _guard21973 = _guard21971 & _guard21972;
wire _guard21974 = fsm_out == 1'd0;
wire _guard21975 = cond_wire315_out;
wire _guard21976 = _guard21974 & _guard21975;
wire _guard21977 = fsm_out == 1'd0;
wire _guard21978 = _guard21976 & _guard21977;
wire _guard21979 = fsm_out == 1'd0;
wire _guard21980 = cond_wire317_out;
wire _guard21981 = _guard21979 & _guard21980;
wire _guard21982 = fsm_out == 1'd0;
wire _guard21983 = _guard21981 & _guard21982;
wire _guard21984 = _guard21978 | _guard21983;
wire _guard21985 = early_reset_static_par0_go_out;
wire _guard21986 = _guard21984 & _guard21985;
wire _guard21987 = cond_wire267_out;
wire _guard21988 = early_reset_static_par0_go_out;
wire _guard21989 = _guard21987 & _guard21988;
wire _guard21990 = cond_wire267_out;
wire _guard21991 = early_reset_static_par0_go_out;
wire _guard21992 = _guard21990 & _guard21991;
wire _guard21993 = cond_wire339_out;
wire _guard21994 = early_reset_static_par0_go_out;
wire _guard21995 = _guard21993 & _guard21994;
wire _guard21996 = cond_wire339_out;
wire _guard21997 = early_reset_static_par0_go_out;
wire _guard21998 = _guard21996 & _guard21997;
wire _guard21999 = cond_wire386_out;
wire _guard22000 = early_reset_static_par0_go_out;
wire _guard22001 = _guard21999 & _guard22000;
wire _guard22002 = cond_wire384_out;
wire _guard22003 = early_reset_static_par0_go_out;
wire _guard22004 = _guard22002 & _guard22003;
wire _guard22005 = fsm_out == 1'd0;
wire _guard22006 = cond_wire384_out;
wire _guard22007 = _guard22005 & _guard22006;
wire _guard22008 = fsm_out == 1'd0;
wire _guard22009 = _guard22007 & _guard22008;
wire _guard22010 = fsm_out == 1'd0;
wire _guard22011 = cond_wire386_out;
wire _guard22012 = _guard22010 & _guard22011;
wire _guard22013 = fsm_out == 1'd0;
wire _guard22014 = _guard22012 & _guard22013;
wire _guard22015 = _guard22009 | _guard22014;
wire _guard22016 = early_reset_static_par0_go_out;
wire _guard22017 = _guard22015 & _guard22016;
wire _guard22018 = fsm_out == 1'd0;
wire _guard22019 = cond_wire384_out;
wire _guard22020 = _guard22018 & _guard22019;
wire _guard22021 = fsm_out == 1'd0;
wire _guard22022 = _guard22020 & _guard22021;
wire _guard22023 = fsm_out == 1'd0;
wire _guard22024 = cond_wire386_out;
wire _guard22025 = _guard22023 & _guard22024;
wire _guard22026 = fsm_out == 1'd0;
wire _guard22027 = _guard22025 & _guard22026;
wire _guard22028 = _guard22022 | _guard22027;
wire _guard22029 = early_reset_static_par0_go_out;
wire _guard22030 = _guard22028 & _guard22029;
wire _guard22031 = fsm_out == 1'd0;
wire _guard22032 = cond_wire384_out;
wire _guard22033 = _guard22031 & _guard22032;
wire _guard22034 = fsm_out == 1'd0;
wire _guard22035 = _guard22033 & _guard22034;
wire _guard22036 = fsm_out == 1'd0;
wire _guard22037 = cond_wire386_out;
wire _guard22038 = _guard22036 & _guard22037;
wire _guard22039 = fsm_out == 1'd0;
wire _guard22040 = _guard22038 & _guard22039;
wire _guard22041 = _guard22035 | _guard22040;
wire _guard22042 = early_reset_static_par0_go_out;
wire _guard22043 = _guard22041 & _guard22042;
wire _guard22044 = cond_wire324_out;
wire _guard22045 = early_reset_static_par0_go_out;
wire _guard22046 = _guard22044 & _guard22045;
wire _guard22047 = cond_wire324_out;
wire _guard22048 = early_reset_static_par0_go_out;
wire _guard22049 = _guard22047 & _guard22048;
wire _guard22050 = cond_wire385_out;
wire _guard22051 = early_reset_static_par0_go_out;
wire _guard22052 = _guard22050 & _guard22051;
wire _guard22053 = cond_wire385_out;
wire _guard22054 = early_reset_static_par0_go_out;
wire _guard22055 = _guard22053 & _guard22054;
wire _guard22056 = cond_wire402_out;
wire _guard22057 = early_reset_static_par0_go_out;
wire _guard22058 = _guard22056 & _guard22057;
wire _guard22059 = cond_wire400_out;
wire _guard22060 = early_reset_static_par0_go_out;
wire _guard22061 = _guard22059 & _guard22060;
wire _guard22062 = fsm_out == 1'd0;
wire _guard22063 = cond_wire400_out;
wire _guard22064 = _guard22062 & _guard22063;
wire _guard22065 = fsm_out == 1'd0;
wire _guard22066 = _guard22064 & _guard22065;
wire _guard22067 = fsm_out == 1'd0;
wire _guard22068 = cond_wire402_out;
wire _guard22069 = _guard22067 & _guard22068;
wire _guard22070 = fsm_out == 1'd0;
wire _guard22071 = _guard22069 & _guard22070;
wire _guard22072 = _guard22066 | _guard22071;
wire _guard22073 = early_reset_static_par0_go_out;
wire _guard22074 = _guard22072 & _guard22073;
wire _guard22075 = fsm_out == 1'd0;
wire _guard22076 = cond_wire400_out;
wire _guard22077 = _guard22075 & _guard22076;
wire _guard22078 = fsm_out == 1'd0;
wire _guard22079 = _guard22077 & _guard22078;
wire _guard22080 = fsm_out == 1'd0;
wire _guard22081 = cond_wire402_out;
wire _guard22082 = _guard22080 & _guard22081;
wire _guard22083 = fsm_out == 1'd0;
wire _guard22084 = _guard22082 & _guard22083;
wire _guard22085 = _guard22079 | _guard22084;
wire _guard22086 = early_reset_static_par0_go_out;
wire _guard22087 = _guard22085 & _guard22086;
wire _guard22088 = fsm_out == 1'd0;
wire _guard22089 = cond_wire400_out;
wire _guard22090 = _guard22088 & _guard22089;
wire _guard22091 = fsm_out == 1'd0;
wire _guard22092 = _guard22090 & _guard22091;
wire _guard22093 = fsm_out == 1'd0;
wire _guard22094 = cond_wire402_out;
wire _guard22095 = _guard22093 & _guard22094;
wire _guard22096 = fsm_out == 1'd0;
wire _guard22097 = _guard22095 & _guard22096;
wire _guard22098 = _guard22092 | _guard22097;
wire _guard22099 = early_reset_static_par0_go_out;
wire _guard22100 = _guard22098 & _guard22099;
wire _guard22101 = cond_wire431_out;
wire _guard22102 = early_reset_static_par0_go_out;
wire _guard22103 = _guard22101 & _guard22102;
wire _guard22104 = cond_wire429_out;
wire _guard22105 = early_reset_static_par0_go_out;
wire _guard22106 = _guard22104 & _guard22105;
wire _guard22107 = fsm_out == 1'd0;
wire _guard22108 = cond_wire429_out;
wire _guard22109 = _guard22107 & _guard22108;
wire _guard22110 = fsm_out == 1'd0;
wire _guard22111 = _guard22109 & _guard22110;
wire _guard22112 = fsm_out == 1'd0;
wire _guard22113 = cond_wire431_out;
wire _guard22114 = _guard22112 & _guard22113;
wire _guard22115 = fsm_out == 1'd0;
wire _guard22116 = _guard22114 & _guard22115;
wire _guard22117 = _guard22111 | _guard22116;
wire _guard22118 = early_reset_static_par0_go_out;
wire _guard22119 = _guard22117 & _guard22118;
wire _guard22120 = fsm_out == 1'd0;
wire _guard22121 = cond_wire429_out;
wire _guard22122 = _guard22120 & _guard22121;
wire _guard22123 = fsm_out == 1'd0;
wire _guard22124 = _guard22122 & _guard22123;
wire _guard22125 = fsm_out == 1'd0;
wire _guard22126 = cond_wire431_out;
wire _guard22127 = _guard22125 & _guard22126;
wire _guard22128 = fsm_out == 1'd0;
wire _guard22129 = _guard22127 & _guard22128;
wire _guard22130 = _guard22124 | _guard22129;
wire _guard22131 = early_reset_static_par0_go_out;
wire _guard22132 = _guard22130 & _guard22131;
wire _guard22133 = fsm_out == 1'd0;
wire _guard22134 = cond_wire429_out;
wire _guard22135 = _guard22133 & _guard22134;
wire _guard22136 = fsm_out == 1'd0;
wire _guard22137 = _guard22135 & _guard22136;
wire _guard22138 = fsm_out == 1'd0;
wire _guard22139 = cond_wire431_out;
wire _guard22140 = _guard22138 & _guard22139;
wire _guard22141 = fsm_out == 1'd0;
wire _guard22142 = _guard22140 & _guard22141;
wire _guard22143 = _guard22137 | _guard22142;
wire _guard22144 = early_reset_static_par0_go_out;
wire _guard22145 = _guard22143 & _guard22144;
wire _guard22146 = cond_wire377_out;
wire _guard22147 = early_reset_static_par0_go_out;
wire _guard22148 = _guard22146 & _guard22147;
wire _guard22149 = cond_wire377_out;
wire _guard22150 = early_reset_static_par0_go_out;
wire _guard22151 = _guard22149 & _guard22150;
wire _guard22152 = cond_wire480_out;
wire _guard22153 = early_reset_static_par0_go_out;
wire _guard22154 = _guard22152 & _guard22153;
wire _guard22155 = cond_wire478_out;
wire _guard22156 = early_reset_static_par0_go_out;
wire _guard22157 = _guard22155 & _guard22156;
wire _guard22158 = fsm_out == 1'd0;
wire _guard22159 = cond_wire478_out;
wire _guard22160 = _guard22158 & _guard22159;
wire _guard22161 = fsm_out == 1'd0;
wire _guard22162 = _guard22160 & _guard22161;
wire _guard22163 = fsm_out == 1'd0;
wire _guard22164 = cond_wire480_out;
wire _guard22165 = _guard22163 & _guard22164;
wire _guard22166 = fsm_out == 1'd0;
wire _guard22167 = _guard22165 & _guard22166;
wire _guard22168 = _guard22162 | _guard22167;
wire _guard22169 = early_reset_static_par0_go_out;
wire _guard22170 = _guard22168 & _guard22169;
wire _guard22171 = fsm_out == 1'd0;
wire _guard22172 = cond_wire478_out;
wire _guard22173 = _guard22171 & _guard22172;
wire _guard22174 = fsm_out == 1'd0;
wire _guard22175 = _guard22173 & _guard22174;
wire _guard22176 = fsm_out == 1'd0;
wire _guard22177 = cond_wire480_out;
wire _guard22178 = _guard22176 & _guard22177;
wire _guard22179 = fsm_out == 1'd0;
wire _guard22180 = _guard22178 & _guard22179;
wire _guard22181 = _guard22175 | _guard22180;
wire _guard22182 = early_reset_static_par0_go_out;
wire _guard22183 = _guard22181 & _guard22182;
wire _guard22184 = fsm_out == 1'd0;
wire _guard22185 = cond_wire478_out;
wire _guard22186 = _guard22184 & _guard22185;
wire _guard22187 = fsm_out == 1'd0;
wire _guard22188 = _guard22186 & _guard22187;
wire _guard22189 = fsm_out == 1'd0;
wire _guard22190 = cond_wire480_out;
wire _guard22191 = _guard22189 & _guard22190;
wire _guard22192 = fsm_out == 1'd0;
wire _guard22193 = _guard22191 & _guard22192;
wire _guard22194 = _guard22188 | _guard22193;
wire _guard22195 = early_reset_static_par0_go_out;
wire _guard22196 = _guard22194 & _guard22195;
wire _guard22197 = cond_wire500_out;
wire _guard22198 = early_reset_static_par0_go_out;
wire _guard22199 = _guard22197 & _guard22198;
wire _guard22200 = cond_wire498_out;
wire _guard22201 = early_reset_static_par0_go_out;
wire _guard22202 = _guard22200 & _guard22201;
wire _guard22203 = fsm_out == 1'd0;
wire _guard22204 = cond_wire498_out;
wire _guard22205 = _guard22203 & _guard22204;
wire _guard22206 = fsm_out == 1'd0;
wire _guard22207 = _guard22205 & _guard22206;
wire _guard22208 = fsm_out == 1'd0;
wire _guard22209 = cond_wire500_out;
wire _guard22210 = _guard22208 & _guard22209;
wire _guard22211 = fsm_out == 1'd0;
wire _guard22212 = _guard22210 & _guard22211;
wire _guard22213 = _guard22207 | _guard22212;
wire _guard22214 = early_reset_static_par0_go_out;
wire _guard22215 = _guard22213 & _guard22214;
wire _guard22216 = fsm_out == 1'd0;
wire _guard22217 = cond_wire498_out;
wire _guard22218 = _guard22216 & _guard22217;
wire _guard22219 = fsm_out == 1'd0;
wire _guard22220 = _guard22218 & _guard22219;
wire _guard22221 = fsm_out == 1'd0;
wire _guard22222 = cond_wire500_out;
wire _guard22223 = _guard22221 & _guard22222;
wire _guard22224 = fsm_out == 1'd0;
wire _guard22225 = _guard22223 & _guard22224;
wire _guard22226 = _guard22220 | _guard22225;
wire _guard22227 = early_reset_static_par0_go_out;
wire _guard22228 = _guard22226 & _guard22227;
wire _guard22229 = fsm_out == 1'd0;
wire _guard22230 = cond_wire498_out;
wire _guard22231 = _guard22229 & _guard22230;
wire _guard22232 = fsm_out == 1'd0;
wire _guard22233 = _guard22231 & _guard22232;
wire _guard22234 = fsm_out == 1'd0;
wire _guard22235 = cond_wire500_out;
wire _guard22236 = _guard22234 & _guard22235;
wire _guard22237 = fsm_out == 1'd0;
wire _guard22238 = _guard22236 & _guard22237;
wire _guard22239 = _guard22233 | _guard22238;
wire _guard22240 = early_reset_static_par0_go_out;
wire _guard22241 = _guard22239 & _guard22240;
wire _guard22242 = cond_wire442_out;
wire _guard22243 = early_reset_static_par0_go_out;
wire _guard22244 = _guard22242 & _guard22243;
wire _guard22245 = cond_wire442_out;
wire _guard22246 = early_reset_static_par0_go_out;
wire _guard22247 = _guard22245 & _guard22246;
wire _guard22248 = cond_wire462_out;
wire _guard22249 = early_reset_static_par0_go_out;
wire _guard22250 = _guard22248 & _guard22249;
wire _guard22251 = cond_wire462_out;
wire _guard22252 = early_reset_static_par0_go_out;
wire _guard22253 = _guard22251 & _guard22252;
wire _guard22254 = cond_wire466_out;
wire _guard22255 = early_reset_static_par0_go_out;
wire _guard22256 = _guard22254 & _guard22255;
wire _guard22257 = cond_wire466_out;
wire _guard22258 = early_reset_static_par0_go_out;
wire _guard22259 = _guard22257 & _guard22258;
wire _guard22260 = cond_wire536_out;
wire _guard22261 = early_reset_static_par0_go_out;
wire _guard22262 = _guard22260 & _guard22261;
wire _guard22263 = cond_wire536_out;
wire _guard22264 = early_reset_static_par0_go_out;
wire _guard22265 = _guard22263 & _guard22264;
wire _guard22266 = cond_wire577_out;
wire _guard22267 = early_reset_static_par0_go_out;
wire _guard22268 = _guard22266 & _guard22267;
wire _guard22269 = cond_wire575_out;
wire _guard22270 = early_reset_static_par0_go_out;
wire _guard22271 = _guard22269 & _guard22270;
wire _guard22272 = fsm_out == 1'd0;
wire _guard22273 = cond_wire575_out;
wire _guard22274 = _guard22272 & _guard22273;
wire _guard22275 = fsm_out == 1'd0;
wire _guard22276 = _guard22274 & _guard22275;
wire _guard22277 = fsm_out == 1'd0;
wire _guard22278 = cond_wire577_out;
wire _guard22279 = _guard22277 & _guard22278;
wire _guard22280 = fsm_out == 1'd0;
wire _guard22281 = _guard22279 & _guard22280;
wire _guard22282 = _guard22276 | _guard22281;
wire _guard22283 = early_reset_static_par0_go_out;
wire _guard22284 = _guard22282 & _guard22283;
wire _guard22285 = fsm_out == 1'd0;
wire _guard22286 = cond_wire575_out;
wire _guard22287 = _guard22285 & _guard22286;
wire _guard22288 = fsm_out == 1'd0;
wire _guard22289 = _guard22287 & _guard22288;
wire _guard22290 = fsm_out == 1'd0;
wire _guard22291 = cond_wire577_out;
wire _guard22292 = _guard22290 & _guard22291;
wire _guard22293 = fsm_out == 1'd0;
wire _guard22294 = _guard22292 & _guard22293;
wire _guard22295 = _guard22289 | _guard22294;
wire _guard22296 = early_reset_static_par0_go_out;
wire _guard22297 = _guard22295 & _guard22296;
wire _guard22298 = fsm_out == 1'd0;
wire _guard22299 = cond_wire575_out;
wire _guard22300 = _guard22298 & _guard22299;
wire _guard22301 = fsm_out == 1'd0;
wire _guard22302 = _guard22300 & _guard22301;
wire _guard22303 = fsm_out == 1'd0;
wire _guard22304 = cond_wire577_out;
wire _guard22305 = _guard22303 & _guard22304;
wire _guard22306 = fsm_out == 1'd0;
wire _guard22307 = _guard22305 & _guard22306;
wire _guard22308 = _guard22302 | _guard22307;
wire _guard22309 = early_reset_static_par0_go_out;
wire _guard22310 = _guard22308 & _guard22309;
wire _guard22311 = cond_wire584_out;
wire _guard22312 = early_reset_static_par0_go_out;
wire _guard22313 = _guard22311 & _guard22312;
wire _guard22314 = cond_wire584_out;
wire _guard22315 = early_reset_static_par0_go_out;
wire _guard22316 = _guard22314 & _guard22315;
wire _guard22317 = cond_wire593_out;
wire _guard22318 = early_reset_static_par0_go_out;
wire _guard22319 = _guard22317 & _guard22318;
wire _guard22320 = cond_wire591_out;
wire _guard22321 = early_reset_static_par0_go_out;
wire _guard22322 = _guard22320 & _guard22321;
wire _guard22323 = fsm_out == 1'd0;
wire _guard22324 = cond_wire591_out;
wire _guard22325 = _guard22323 & _guard22324;
wire _guard22326 = fsm_out == 1'd0;
wire _guard22327 = _guard22325 & _guard22326;
wire _guard22328 = fsm_out == 1'd0;
wire _guard22329 = cond_wire593_out;
wire _guard22330 = _guard22328 & _guard22329;
wire _guard22331 = fsm_out == 1'd0;
wire _guard22332 = _guard22330 & _guard22331;
wire _guard22333 = _guard22327 | _guard22332;
wire _guard22334 = early_reset_static_par0_go_out;
wire _guard22335 = _guard22333 & _guard22334;
wire _guard22336 = fsm_out == 1'd0;
wire _guard22337 = cond_wire591_out;
wire _guard22338 = _guard22336 & _guard22337;
wire _guard22339 = fsm_out == 1'd0;
wire _guard22340 = _guard22338 & _guard22339;
wire _guard22341 = fsm_out == 1'd0;
wire _guard22342 = cond_wire593_out;
wire _guard22343 = _guard22341 & _guard22342;
wire _guard22344 = fsm_out == 1'd0;
wire _guard22345 = _guard22343 & _guard22344;
wire _guard22346 = _guard22340 | _guard22345;
wire _guard22347 = early_reset_static_par0_go_out;
wire _guard22348 = _guard22346 & _guard22347;
wire _guard22349 = fsm_out == 1'd0;
wire _guard22350 = cond_wire591_out;
wire _guard22351 = _guard22349 & _guard22350;
wire _guard22352 = fsm_out == 1'd0;
wire _guard22353 = _guard22351 & _guard22352;
wire _guard22354 = fsm_out == 1'd0;
wire _guard22355 = cond_wire593_out;
wire _guard22356 = _guard22354 & _guard22355;
wire _guard22357 = fsm_out == 1'd0;
wire _guard22358 = _guard22356 & _guard22357;
wire _guard22359 = _guard22353 | _guard22358;
wire _guard22360 = early_reset_static_par0_go_out;
wire _guard22361 = _guard22359 & _guard22360;
wire _guard22362 = cond_wire544_out;
wire _guard22363 = early_reset_static_par0_go_out;
wire _guard22364 = _guard22362 & _guard22363;
wire _guard22365 = cond_wire544_out;
wire _guard22366 = early_reset_static_par0_go_out;
wire _guard22367 = _guard22365 & _guard22366;
wire _guard22368 = cond_wire641_out;
wire _guard22369 = early_reset_static_par0_go_out;
wire _guard22370 = _guard22368 & _guard22369;
wire _guard22371 = cond_wire641_out;
wire _guard22372 = early_reset_static_par0_go_out;
wire _guard22373 = _guard22371 & _guard22372;
wire _guard22374 = cond_wire666_out;
wire _guard22375 = early_reset_static_par0_go_out;
wire _guard22376 = _guard22374 & _guard22375;
wire _guard22377 = cond_wire666_out;
wire _guard22378 = early_reset_static_par0_go_out;
wire _guard22379 = _guard22377 & _guard22378;
wire _guard22380 = cond_wire711_out;
wire _guard22381 = early_reset_static_par0_go_out;
wire _guard22382 = _guard22380 & _guard22381;
wire _guard22383 = cond_wire709_out;
wire _guard22384 = early_reset_static_par0_go_out;
wire _guard22385 = _guard22383 & _guard22384;
wire _guard22386 = fsm_out == 1'd0;
wire _guard22387 = cond_wire709_out;
wire _guard22388 = _guard22386 & _guard22387;
wire _guard22389 = fsm_out == 1'd0;
wire _guard22390 = _guard22388 & _guard22389;
wire _guard22391 = fsm_out == 1'd0;
wire _guard22392 = cond_wire711_out;
wire _guard22393 = _guard22391 & _guard22392;
wire _guard22394 = fsm_out == 1'd0;
wire _guard22395 = _guard22393 & _guard22394;
wire _guard22396 = _guard22390 | _guard22395;
wire _guard22397 = early_reset_static_par0_go_out;
wire _guard22398 = _guard22396 & _guard22397;
wire _guard22399 = fsm_out == 1'd0;
wire _guard22400 = cond_wire709_out;
wire _guard22401 = _guard22399 & _guard22400;
wire _guard22402 = fsm_out == 1'd0;
wire _guard22403 = _guard22401 & _guard22402;
wire _guard22404 = fsm_out == 1'd0;
wire _guard22405 = cond_wire711_out;
wire _guard22406 = _guard22404 & _guard22405;
wire _guard22407 = fsm_out == 1'd0;
wire _guard22408 = _guard22406 & _guard22407;
wire _guard22409 = _guard22403 | _guard22408;
wire _guard22410 = early_reset_static_par0_go_out;
wire _guard22411 = _guard22409 & _guard22410;
wire _guard22412 = fsm_out == 1'd0;
wire _guard22413 = cond_wire709_out;
wire _guard22414 = _guard22412 & _guard22413;
wire _guard22415 = fsm_out == 1'd0;
wire _guard22416 = _guard22414 & _guard22415;
wire _guard22417 = fsm_out == 1'd0;
wire _guard22418 = cond_wire711_out;
wire _guard22419 = _guard22417 & _guard22418;
wire _guard22420 = fsm_out == 1'd0;
wire _guard22421 = _guard22419 & _guard22420;
wire _guard22422 = _guard22416 | _guard22421;
wire _guard22423 = early_reset_static_par0_go_out;
wire _guard22424 = _guard22422 & _guard22423;
wire _guard22425 = cond_wire645_out;
wire _guard22426 = early_reset_static_par0_go_out;
wire _guard22427 = _guard22425 & _guard22426;
wire _guard22428 = cond_wire645_out;
wire _guard22429 = early_reset_static_par0_go_out;
wire _guard22430 = _guard22428 & _guard22429;
wire _guard22431 = cond_wire710_out;
wire _guard22432 = early_reset_static_par0_go_out;
wire _guard22433 = _guard22431 & _guard22432;
wire _guard22434 = cond_wire710_out;
wire _guard22435 = early_reset_static_par0_go_out;
wire _guard22436 = _guard22434 & _guard22435;
wire _guard22437 = cond_wire666_out;
wire _guard22438 = early_reset_static_par0_go_out;
wire _guard22439 = _guard22437 & _guard22438;
wire _guard22440 = cond_wire666_out;
wire _guard22441 = early_reset_static_par0_go_out;
wire _guard22442 = _guard22440 & _guard22441;
wire _guard22443 = cond_wire731_out;
wire _guard22444 = early_reset_static_par0_go_out;
wire _guard22445 = _guard22443 & _guard22444;
wire _guard22446 = cond_wire731_out;
wire _guard22447 = early_reset_static_par0_go_out;
wire _guard22448 = _guard22446 & _guard22447;
wire _guard22449 = cond_wire772_out;
wire _guard22450 = early_reset_static_par0_go_out;
wire _guard22451 = _guard22449 & _guard22450;
wire _guard22452 = cond_wire770_out;
wire _guard22453 = early_reset_static_par0_go_out;
wire _guard22454 = _guard22452 & _guard22453;
wire _guard22455 = fsm_out == 1'd0;
wire _guard22456 = cond_wire770_out;
wire _guard22457 = _guard22455 & _guard22456;
wire _guard22458 = fsm_out == 1'd0;
wire _guard22459 = _guard22457 & _guard22458;
wire _guard22460 = fsm_out == 1'd0;
wire _guard22461 = cond_wire772_out;
wire _guard22462 = _guard22460 & _guard22461;
wire _guard22463 = fsm_out == 1'd0;
wire _guard22464 = _guard22462 & _guard22463;
wire _guard22465 = _guard22459 | _guard22464;
wire _guard22466 = early_reset_static_par0_go_out;
wire _guard22467 = _guard22465 & _guard22466;
wire _guard22468 = fsm_out == 1'd0;
wire _guard22469 = cond_wire770_out;
wire _guard22470 = _guard22468 & _guard22469;
wire _guard22471 = fsm_out == 1'd0;
wire _guard22472 = _guard22470 & _guard22471;
wire _guard22473 = fsm_out == 1'd0;
wire _guard22474 = cond_wire772_out;
wire _guard22475 = _guard22473 & _guard22474;
wire _guard22476 = fsm_out == 1'd0;
wire _guard22477 = _guard22475 & _guard22476;
wire _guard22478 = _guard22472 | _guard22477;
wire _guard22479 = early_reset_static_par0_go_out;
wire _guard22480 = _guard22478 & _guard22479;
wire _guard22481 = fsm_out == 1'd0;
wire _guard22482 = cond_wire770_out;
wire _guard22483 = _guard22481 & _guard22482;
wire _guard22484 = fsm_out == 1'd0;
wire _guard22485 = _guard22483 & _guard22484;
wire _guard22486 = fsm_out == 1'd0;
wire _guard22487 = cond_wire772_out;
wire _guard22488 = _guard22486 & _guard22487;
wire _guard22489 = fsm_out == 1'd0;
wire _guard22490 = _guard22488 & _guard22489;
wire _guard22491 = _guard22485 | _guard22490;
wire _guard22492 = early_reset_static_par0_go_out;
wire _guard22493 = _guard22491 & _guard22492;
wire _guard22494 = cond_wire852_out;
wire _guard22495 = early_reset_static_par0_go_out;
wire _guard22496 = _guard22494 & _guard22495;
wire _guard22497 = cond_wire852_out;
wire _guard22498 = early_reset_static_par0_go_out;
wire _guard22499 = _guard22497 & _guard22498;
wire _guard22500 = cond_wire924_out;
wire _guard22501 = early_reset_static_par0_go_out;
wire _guard22502 = _guard22500 & _guard22501;
wire _guard22503 = cond_wire924_out;
wire _guard22504 = early_reset_static_par0_go_out;
wire _guard22505 = _guard22503 & _guard22504;
wire _guard22506 = cond_wire869_out;
wire _guard22507 = early_reset_static_par0_go_out;
wire _guard22508 = _guard22506 & _guard22507;
wire _guard22509 = cond_wire869_out;
wire _guard22510 = early_reset_static_par0_go_out;
wire _guard22511 = _guard22509 & _guard22510;
wire _guard22512 = cond_wire873_out;
wire _guard22513 = early_reset_static_par0_go_out;
wire _guard22514 = _guard22512 & _guard22513;
wire _guard22515 = cond_wire873_out;
wire _guard22516 = early_reset_static_par0_go_out;
wire _guard22517 = _guard22515 & _guard22516;
wire _guard22518 = cond_wire1003_out;
wire _guard22519 = early_reset_static_par0_go_out;
wire _guard22520 = _guard22518 & _guard22519;
wire _guard22521 = cond_wire1003_out;
wire _guard22522 = early_reset_static_par0_go_out;
wire _guard22523 = _guard22521 & _guard22522;
wire _guard22524 = cond_wire1020_out;
wire _guard22525 = early_reset_static_par0_go_out;
wire _guard22526 = _guard22524 & _guard22525;
wire _guard22527 = cond_wire1018_out;
wire _guard22528 = early_reset_static_par0_go_out;
wire _guard22529 = _guard22527 & _guard22528;
wire _guard22530 = fsm_out == 1'd0;
wire _guard22531 = cond_wire1018_out;
wire _guard22532 = _guard22530 & _guard22531;
wire _guard22533 = fsm_out == 1'd0;
wire _guard22534 = _guard22532 & _guard22533;
wire _guard22535 = fsm_out == 1'd0;
wire _guard22536 = cond_wire1020_out;
wire _guard22537 = _guard22535 & _guard22536;
wire _guard22538 = fsm_out == 1'd0;
wire _guard22539 = _guard22537 & _guard22538;
wire _guard22540 = _guard22534 | _guard22539;
wire _guard22541 = early_reset_static_par0_go_out;
wire _guard22542 = _guard22540 & _guard22541;
wire _guard22543 = fsm_out == 1'd0;
wire _guard22544 = cond_wire1018_out;
wire _guard22545 = _guard22543 & _guard22544;
wire _guard22546 = fsm_out == 1'd0;
wire _guard22547 = _guard22545 & _guard22546;
wire _guard22548 = fsm_out == 1'd0;
wire _guard22549 = cond_wire1020_out;
wire _guard22550 = _guard22548 & _guard22549;
wire _guard22551 = fsm_out == 1'd0;
wire _guard22552 = _guard22550 & _guard22551;
wire _guard22553 = _guard22547 | _guard22552;
wire _guard22554 = early_reset_static_par0_go_out;
wire _guard22555 = _guard22553 & _guard22554;
wire _guard22556 = fsm_out == 1'd0;
wire _guard22557 = cond_wire1018_out;
wire _guard22558 = _guard22556 & _guard22557;
wire _guard22559 = fsm_out == 1'd0;
wire _guard22560 = _guard22558 & _guard22559;
wire _guard22561 = fsm_out == 1'd0;
wire _guard22562 = cond_wire1020_out;
wire _guard22563 = _guard22561 & _guard22562;
wire _guard22564 = fsm_out == 1'd0;
wire _guard22565 = _guard22563 & _guard22564;
wire _guard22566 = _guard22560 | _guard22565;
wire _guard22567 = early_reset_static_par0_go_out;
wire _guard22568 = _guard22566 & _guard22567;
wire _guard22569 = fsm0_out == 6'd0;
wire _guard22570 = early_reset_static_seq_go_out;
wire _guard22571 = _guard22569 & _guard22570;
wire _guard22572 = cond_wire9_out;
wire _guard22573 = early_reset_static_par0_go_out;
wire _guard22574 = _guard22572 & _guard22573;
wire _guard22575 = _guard22571 | _guard22574;
wire _guard22576 = fsm0_out == 6'd0;
wire _guard22577 = early_reset_static_seq_go_out;
wire _guard22578 = _guard22576 & _guard22577;
wire _guard22579 = cond_wire9_out;
wire _guard22580 = early_reset_static_par0_go_out;
wire _guard22581 = _guard22579 & _guard22580;
wire _guard22582 = cond_wire54_out;
wire _guard22583 = early_reset_static_par0_go_out;
wire _guard22584 = _guard22582 & _guard22583;
wire _guard22585 = cond_wire54_out;
wire _guard22586 = early_reset_static_par0_go_out;
wire _guard22587 = _guard22585 & _guard22586;
wire _guard22588 = fsm0_out == 6'd0;
wire _guard22589 = early_reset_static_seq_go_out;
wire _guard22590 = _guard22588 & _guard22589;
wire _guard22591 = cond_wire144_out;
wire _guard22592 = early_reset_static_par0_go_out;
wire _guard22593 = _guard22591 & _guard22592;
wire _guard22594 = _guard22590 | _guard22593;
wire _guard22595 = fsm0_out == 6'd0;
wire _guard22596 = early_reset_static_seq_go_out;
wire _guard22597 = _guard22595 & _guard22596;
wire _guard22598 = cond_wire144_out;
wire _guard22599 = early_reset_static_par0_go_out;
wire _guard22600 = _guard22598 & _guard22599;
wire _guard22601 = fsm0_out == 6'd0;
wire _guard22602 = early_reset_static_seq_go_out;
wire _guard22603 = _guard22601 & _guard22602;
wire _guard22604 = cond_wire404_out;
wire _guard22605 = early_reset_static_par0_go_out;
wire _guard22606 = _guard22604 & _guard22605;
wire _guard22607 = _guard22603 | _guard22606;
wire _guard22608 = fsm0_out == 6'd0;
wire _guard22609 = early_reset_static_seq_go_out;
wire _guard22610 = _guard22608 & _guard22609;
wire _guard22611 = cond_wire404_out;
wire _guard22612 = early_reset_static_par0_go_out;
wire _guard22613 = _guard22611 & _guard22612;
wire _guard22614 = cond_wire924_out;
wire _guard22615 = early_reset_static_par0_go_out;
wire _guard22616 = _guard22614 & _guard22615;
wire _guard22617 = cond_wire924_out;
wire _guard22618 = early_reset_static_par0_go_out;
wire _guard22619 = _guard22617 & _guard22618;
wire _guard22620 = early_reset_static_par0_go_out;
wire _guard22621 = early_reset_static_par0_go_out;
wire _guard22622 = early_reset_static_par0_go_out;
wire _guard22623 = early_reset_static_par0_go_out;
wire _guard22624 = fsm0_out == 6'd0;
wire _guard22625 = early_reset_static_seq_go_out;
wire _guard22626 = _guard22624 & _guard22625;
wire _guard22627 = early_reset_static_par0_go_out;
wire _guard22628 = _guard22626 | _guard22627;
wire _guard22629 = fsm0_out == 6'd0;
wire _guard22630 = early_reset_static_seq_go_out;
wire _guard22631 = _guard22629 & _guard22630;
wire _guard22632 = early_reset_static_par0_go_out;
wire _guard22633 = early_reset_static_par0_go_out;
wire _guard22634 = early_reset_static_par0_go_out;
wire _guard22635 = fsm0_out == 6'd0;
wire _guard22636 = early_reset_static_seq_go_out;
wire _guard22637 = _guard22635 & _guard22636;
wire _guard22638 = early_reset_static_par0_go_out;
wire _guard22639 = _guard22637 | _guard22638;
wire _guard22640 = fsm0_out == 6'd0;
wire _guard22641 = early_reset_static_seq_go_out;
wire _guard22642 = _guard22640 & _guard22641;
wire _guard22643 = early_reset_static_par0_go_out;
wire _guard22644 = early_reset_static_par0_go_out;
wire _guard22645 = early_reset_static_par0_go_out;
wire _guard22646 = early_reset_static_par0_go_out;
wire _guard22647 = early_reset_static_par0_go_out;
wire _guard22648 = early_reset_static_par0_go_out;
wire _guard22649 = early_reset_static_par0_go_out;
wire _guard22650 = fsm0_out == 6'd0;
wire _guard22651 = early_reset_static_seq_go_out;
wire _guard22652 = _guard22650 & _guard22651;
wire _guard22653 = early_reset_static_par0_go_out;
wire _guard22654 = _guard22652 | _guard22653;
wire _guard22655 = early_reset_static_par0_go_out;
wire _guard22656 = fsm0_out == 6'd0;
wire _guard22657 = early_reset_static_seq_go_out;
wire _guard22658 = _guard22656 & _guard22657;
wire _guard22659 = early_reset_static_par0_go_out;
wire _guard22660 = early_reset_static_par0_go_out;
wire _guard22661 = early_reset_static_par0_go_out;
wire _guard22662 = early_reset_static_par0_go_out;
wire _guard22663 = fsm0_out == 6'd0;
wire _guard22664 = early_reset_static_seq_go_out;
wire _guard22665 = _guard22663 & _guard22664;
wire _guard22666 = early_reset_static_par0_go_out;
wire _guard22667 = _guard22665 | _guard22666;
wire _guard22668 = early_reset_static_par0_go_out;
wire _guard22669 = fsm0_out == 6'd0;
wire _guard22670 = early_reset_static_seq_go_out;
wire _guard22671 = _guard22669 & _guard22670;
wire _guard22672 = early_reset_static_par0_go_out;
wire _guard22673 = early_reset_static_par0_go_out;
wire _guard22674 = early_reset_static_par0_go_out;
wire _guard22675 = early_reset_static_par0_go_out;
wire _guard22676 = fsm0_out == 6'd0;
wire _guard22677 = early_reset_static_seq_go_out;
wire _guard22678 = _guard22676 & _guard22677;
wire _guard22679 = early_reset_static_par0_go_out;
wire _guard22680 = _guard22678 | _guard22679;
wire _guard22681 = fsm0_out == 6'd0;
wire _guard22682 = early_reset_static_seq_go_out;
wire _guard22683 = _guard22681 & _guard22682;
wire _guard22684 = early_reset_static_par0_go_out;
wire _guard22685 = fsm0_out == 6'd0;
wire _guard22686 = early_reset_static_seq_go_out;
wire _guard22687 = _guard22685 & _guard22686;
wire _guard22688 = early_reset_static_par0_go_out;
wire _guard22689 = _guard22687 | _guard22688;
wire _guard22690 = fsm0_out == 6'd0;
wire _guard22691 = early_reset_static_seq_go_out;
wire _guard22692 = _guard22690 & _guard22691;
wire _guard22693 = early_reset_static_par0_go_out;
wire _guard22694 = early_reset_static_par0_go_out;
wire _guard22695 = early_reset_static_par0_go_out;
wire _guard22696 = early_reset_static_par0_go_out;
wire _guard22697 = early_reset_static_par0_go_out;
wire _guard22698 = early_reset_static_par0_go_out;
wire _guard22699 = early_reset_static_par0_go_out;
wire _guard22700 = fsm0_out == 6'd0;
wire _guard22701 = early_reset_static_seq_go_out;
wire _guard22702 = _guard22700 & _guard22701;
wire _guard22703 = early_reset_static_par0_go_out;
wire _guard22704 = _guard22702 | _guard22703;
wire _guard22705 = early_reset_static_par0_go_out;
wire _guard22706 = fsm0_out == 6'd0;
wire _guard22707 = early_reset_static_seq_go_out;
wire _guard22708 = _guard22706 & _guard22707;
wire _guard22709 = early_reset_static_par0_go_out;
wire _guard22710 = early_reset_static_par0_go_out;
wire _guard22711 = early_reset_static_par0_go_out;
wire _guard22712 = early_reset_static_par0_go_out;
wire _guard22713 = ~_guard0;
wire _guard22714 = early_reset_static_par0_go_out;
wire _guard22715 = _guard22713 & _guard22714;
wire _guard22716 = early_reset_static_par0_go_out;
wire _guard22717 = early_reset_static_par0_go_out;
wire _guard22718 = early_reset_static_par0_go_out;
wire _guard22719 = early_reset_static_par0_go_out;
wire _guard22720 = early_reset_static_par0_go_out;
wire _guard22721 = early_reset_static_par0_go_out;
wire _guard22722 = ~_guard0;
wire _guard22723 = early_reset_static_par0_go_out;
wire _guard22724 = _guard22722 & _guard22723;
wire _guard22725 = early_reset_static_par0_go_out;
wire _guard22726 = early_reset_static_par0_go_out;
wire _guard22727 = early_reset_static_par0_go_out;
wire _guard22728 = early_reset_static_par0_go_out;
wire _guard22729 = ~_guard0;
wire _guard22730 = early_reset_static_par0_go_out;
wire _guard22731 = _guard22729 & _guard22730;
wire _guard22732 = early_reset_static_par0_go_out;
wire _guard22733 = early_reset_static_par0_go_out;
wire _guard22734 = ~_guard0;
wire _guard22735 = early_reset_static_par0_go_out;
wire _guard22736 = _guard22734 & _guard22735;
wire _guard22737 = early_reset_static_par0_go_out;
wire _guard22738 = ~_guard0;
wire _guard22739 = early_reset_static_par0_go_out;
wire _guard22740 = _guard22738 & _guard22739;
wire _guard22741 = early_reset_static_par0_go_out;
wire _guard22742 = ~_guard0;
wire _guard22743 = early_reset_static_par0_go_out;
wire _guard22744 = _guard22742 & _guard22743;
wire _guard22745 = early_reset_static_par0_go_out;
wire _guard22746 = early_reset_static_par0_go_out;
wire _guard22747 = early_reset_static_par0_go_out;
wire _guard22748 = early_reset_static_par0_go_out;
wire _guard22749 = early_reset_static_par0_go_out;
wire _guard22750 = ~_guard0;
wire _guard22751 = early_reset_static_par0_go_out;
wire _guard22752 = _guard22750 & _guard22751;
wire _guard22753 = early_reset_static_par0_go_out;
wire _guard22754 = early_reset_static_par0_go_out;
wire _guard22755 = early_reset_static_par0_go_out;
wire _guard22756 = early_reset_static_par0_go_out;
wire _guard22757 = early_reset_static_par0_go_out;
wire _guard22758 = early_reset_static_par0_go_out;
wire _guard22759 = early_reset_static_par0_go_out;
wire _guard22760 = early_reset_static_par0_go_out;
wire _guard22761 = early_reset_static_par0_go_out;
wire _guard22762 = early_reset_static_par0_go_out;
wire _guard22763 = early_reset_static_par0_go_out;
wire _guard22764 = early_reset_static_par0_go_out;
wire _guard22765 = early_reset_static_par0_go_out;
wire _guard22766 = ~_guard0;
wire _guard22767 = early_reset_static_par0_go_out;
wire _guard22768 = _guard22766 & _guard22767;
wire _guard22769 = early_reset_static_par0_go_out;
wire _guard22770 = early_reset_static_par0_go_out;
wire _guard22771 = early_reset_static_par0_go_out;
wire _guard22772 = early_reset_static_par0_go_out;
wire _guard22773 = ~_guard0;
wire _guard22774 = early_reset_static_par0_go_out;
wire _guard22775 = _guard22773 & _guard22774;
wire _guard22776 = early_reset_static_par0_go_out;
wire _guard22777 = early_reset_static_par0_go_out;
wire _guard22778 = early_reset_static_par0_go_out;
wire _guard22779 = early_reset_static_par0_go_out;
wire _guard22780 = early_reset_static_par0_go_out;
wire _guard22781 = early_reset_static_par0_go_out;
wire _guard22782 = early_reset_static_par0_go_out;
wire _guard22783 = early_reset_static_par0_go_out;
wire _guard22784 = ~_guard0;
wire _guard22785 = early_reset_static_par0_go_out;
wire _guard22786 = _guard22784 & _guard22785;
wire _guard22787 = ~_guard0;
wire _guard22788 = early_reset_static_par0_go_out;
wire _guard22789 = _guard22787 & _guard22788;
wire _guard22790 = early_reset_static_par0_go_out;
wire _guard22791 = early_reset_static_par0_go_out;
wire _guard22792 = early_reset_static_par0_go_out;
wire _guard22793 = early_reset_static_par0_go_out;
wire _guard22794 = ~_guard0;
wire _guard22795 = early_reset_static_par0_go_out;
wire _guard22796 = _guard22794 & _guard22795;
wire _guard22797 = early_reset_static_par0_go_out;
wire _guard22798 = early_reset_static_par0_go_out;
wire _guard22799 = ~_guard0;
wire _guard22800 = early_reset_static_par0_go_out;
wire _guard22801 = _guard22799 & _guard22800;
wire _guard22802 = early_reset_static_par0_go_out;
wire _guard22803 = early_reset_static_par0_go_out;
wire _guard22804 = ~_guard0;
wire _guard22805 = early_reset_static_par0_go_out;
wire _guard22806 = _guard22804 & _guard22805;
wire _guard22807 = early_reset_static_par0_go_out;
wire _guard22808 = ~_guard0;
wire _guard22809 = early_reset_static_par0_go_out;
wire _guard22810 = _guard22808 & _guard22809;
wire _guard22811 = early_reset_static_par0_go_out;
wire _guard22812 = early_reset_static_par0_go_out;
wire _guard22813 = early_reset_static_par0_go_out;
wire _guard22814 = ~_guard0;
wire _guard22815 = early_reset_static_par0_go_out;
wire _guard22816 = _guard22814 & _guard22815;
wire _guard22817 = early_reset_static_par0_go_out;
wire _guard22818 = early_reset_static_par0_go_out;
wire _guard22819 = early_reset_static_par0_go_out;
wire _guard22820 = early_reset_static_par0_go_out;
wire _guard22821 = ~_guard0;
wire _guard22822 = early_reset_static_par0_go_out;
wire _guard22823 = _guard22821 & _guard22822;
wire _guard22824 = early_reset_static_par0_go_out;
wire _guard22825 = early_reset_static_par0_go_out;
wire _guard22826 = ~_guard0;
wire _guard22827 = early_reset_static_par0_go_out;
wire _guard22828 = _guard22826 & _guard22827;
wire _guard22829 = early_reset_static_par0_go_out;
wire _guard22830 = early_reset_static_par0_go_out;
wire _guard22831 = early_reset_static_par0_go_out;
wire _guard22832 = early_reset_static_par0_go_out;
wire _guard22833 = early_reset_static_par0_go_out;
wire _guard22834 = early_reset_static_par0_go_out;
wire _guard22835 = early_reset_static_par0_go_out;
wire _guard22836 = early_reset_static_par0_go_out;
wire _guard22837 = early_reset_static_par0_go_out;
wire _guard22838 = early_reset_static_par0_go_out;
wire _guard22839 = early_reset_static_par0_go_out;
wire _guard22840 = early_reset_static_par0_go_out;
wire _guard22841 = early_reset_static_par0_go_out;
wire _guard22842 = early_reset_static_par0_go_out;
wire _guard22843 = ~_guard0;
wire _guard22844 = early_reset_static_par0_go_out;
wire _guard22845 = _guard22843 & _guard22844;
wire _guard22846 = early_reset_static_par0_go_out;
wire _guard22847 = early_reset_static_par0_go_out;
wire _guard22848 = early_reset_static_par0_go_out;
wire _guard22849 = early_reset_static_par0_go_out;
wire _guard22850 = early_reset_static_par0_go_out;
wire _guard22851 = early_reset_static_par0_go_out;
wire _guard22852 = early_reset_static_par0_go_out;
wire _guard22853 = early_reset_static_par0_go_out;
wire _guard22854 = early_reset_static_par0_go_out;
wire _guard22855 = early_reset_static_par0_go_out;
wire _guard22856 = ~_guard0;
wire _guard22857 = early_reset_static_par0_go_out;
wire _guard22858 = _guard22856 & _guard22857;
wire _guard22859 = ~_guard0;
wire _guard22860 = early_reset_static_par0_go_out;
wire _guard22861 = _guard22859 & _guard22860;
wire _guard22862 = early_reset_static_par0_go_out;
wire _guard22863 = early_reset_static_par0_go_out;
wire _guard22864 = early_reset_static_par0_go_out;
wire _guard22865 = early_reset_static_par0_go_out;
wire _guard22866 = early_reset_static_par0_go_out;
wire _guard22867 = early_reset_static_par0_go_out;
wire _guard22868 = early_reset_static_par0_go_out;
wire _guard22869 = ~_guard0;
wire _guard22870 = early_reset_static_par0_go_out;
wire _guard22871 = _guard22869 & _guard22870;
wire _guard22872 = early_reset_static_par0_go_out;
wire _guard22873 = early_reset_static_par0_go_out;
wire _guard22874 = early_reset_static_par0_go_out;
wire _guard22875 = ~_guard0;
wire _guard22876 = early_reset_static_par0_go_out;
wire _guard22877 = _guard22875 & _guard22876;
wire _guard22878 = early_reset_static_par0_go_out;
wire _guard22879 = early_reset_static_par0_go_out;
wire _guard22880 = ~_guard0;
wire _guard22881 = early_reset_static_par0_go_out;
wire _guard22882 = _guard22880 & _guard22881;
wire _guard22883 = ~_guard0;
wire _guard22884 = early_reset_static_par0_go_out;
wire _guard22885 = _guard22883 & _guard22884;
wire _guard22886 = early_reset_static_par0_go_out;
wire _guard22887 = early_reset_static_par0_go_out;
wire _guard22888 = early_reset_static_par0_go_out;
wire _guard22889 = early_reset_static_par0_go_out;
wire _guard22890 = early_reset_static_par0_go_out;
wire _guard22891 = early_reset_static_par0_go_out;
wire _guard22892 = ~_guard0;
wire _guard22893 = early_reset_static_par0_go_out;
wire _guard22894 = _guard22892 & _guard22893;
wire _guard22895 = early_reset_static_par0_go_out;
wire _guard22896 = early_reset_static_par0_go_out;
wire _guard22897 = early_reset_static_par0_go_out;
wire _guard22898 = early_reset_static_par0_go_out;
wire _guard22899 = early_reset_static_par0_go_out;
wire _guard22900 = ~_guard0;
wire _guard22901 = early_reset_static_par0_go_out;
wire _guard22902 = _guard22900 & _guard22901;
wire _guard22903 = early_reset_static_par0_go_out;
wire _guard22904 = early_reset_static_par0_go_out;
wire _guard22905 = early_reset_static_par0_go_out;
wire _guard22906 = early_reset_static_par0_go_out;
wire _guard22907 = early_reset_static_par0_go_out;
wire _guard22908 = early_reset_static_par0_go_out;
wire _guard22909 = ~_guard0;
wire _guard22910 = early_reset_static_par0_go_out;
wire _guard22911 = _guard22909 & _guard22910;
wire _guard22912 = early_reset_static_par0_go_out;
wire _guard22913 = ~_guard0;
wire _guard22914 = early_reset_static_par0_go_out;
wire _guard22915 = _guard22913 & _guard22914;
wire _guard22916 = early_reset_static_par0_go_out;
wire _guard22917 = early_reset_static_par0_go_out;
wire _guard22918 = early_reset_static_par0_go_out;
wire _guard22919 = early_reset_static_par0_go_out;
wire _guard22920 = ~_guard0;
wire _guard22921 = early_reset_static_par0_go_out;
wire _guard22922 = _guard22920 & _guard22921;
wire _guard22923 = early_reset_static_par0_go_out;
wire _guard22924 = early_reset_static_par0_go_out;
wire _guard22925 = ~_guard0;
wire _guard22926 = early_reset_static_par0_go_out;
wire _guard22927 = _guard22925 & _guard22926;
wire _guard22928 = early_reset_static_par0_go_out;
wire _guard22929 = early_reset_static_par0_go_out;
wire _guard22930 = early_reset_static_par0_go_out;
wire _guard22931 = early_reset_static_par0_go_out;
wire _guard22932 = ~_guard0;
wire _guard22933 = early_reset_static_par0_go_out;
wire _guard22934 = _guard22932 & _guard22933;
wire _guard22935 = ~_guard0;
wire _guard22936 = early_reset_static_par0_go_out;
wire _guard22937 = _guard22935 & _guard22936;
wire _guard22938 = early_reset_static_par0_go_out;
wire _guard22939 = early_reset_static_par0_go_out;
wire _guard22940 = early_reset_static_par0_go_out;
wire _guard22941 = early_reset_static_par0_go_out;
wire _guard22942 = ~_guard0;
wire _guard22943 = early_reset_static_par0_go_out;
wire _guard22944 = _guard22942 & _guard22943;
wire _guard22945 = early_reset_static_par0_go_out;
wire _guard22946 = early_reset_static_par0_go_out;
wire _guard22947 = ~_guard0;
wire _guard22948 = early_reset_static_par0_go_out;
wire _guard22949 = _guard22947 & _guard22948;
wire _guard22950 = early_reset_static_par0_go_out;
wire _guard22951 = ~_guard0;
wire _guard22952 = early_reset_static_par0_go_out;
wire _guard22953 = _guard22951 & _guard22952;
wire _guard22954 = early_reset_static_par0_go_out;
wire _guard22955 = early_reset_static_par0_go_out;
wire _guard22956 = ~_guard0;
wire _guard22957 = early_reset_static_par0_go_out;
wire _guard22958 = _guard22956 & _guard22957;
wire _guard22959 = early_reset_static_par0_go_out;
wire _guard22960 = early_reset_static_par0_go_out;
wire _guard22961 = early_reset_static_par0_go_out;
wire _guard22962 = ~_guard0;
wire _guard22963 = early_reset_static_par0_go_out;
wire _guard22964 = _guard22962 & _guard22963;
wire _guard22965 = early_reset_static_par0_go_out;
wire _guard22966 = early_reset_static_par0_go_out;
wire _guard22967 = early_reset_static_par0_go_out;
wire _guard22968 = ~_guard0;
wire _guard22969 = early_reset_static_par0_go_out;
wire _guard22970 = _guard22968 & _guard22969;
wire _guard22971 = early_reset_static_par0_go_out;
wire _guard22972 = early_reset_static_par0_go_out;
wire _guard22973 = early_reset_static_par0_go_out;
wire _guard22974 = early_reset_static_par0_go_out;
wire _guard22975 = early_reset_static_par0_go_out;
wire _guard22976 = early_reset_static_par0_go_out;
wire _guard22977 = ~_guard0;
wire _guard22978 = early_reset_static_par0_go_out;
wire _guard22979 = _guard22977 & _guard22978;
wire _guard22980 = early_reset_static_par0_go_out;
wire _guard22981 = early_reset_static_par0_go_out;
wire _guard22982 = early_reset_static_par0_go_out;
wire _guard22983 = early_reset_static_par0_go_out;
wire _guard22984 = early_reset_static_par0_go_out;
wire _guard22985 = early_reset_static_par0_go_out;
wire _guard22986 = early_reset_static_par0_go_out;
wire _guard22987 = early_reset_static_par0_go_out;
wire _guard22988 = early_reset_static_par0_go_out;
wire _guard22989 = early_reset_static_par0_go_out;
wire _guard22990 = ~_guard0;
wire _guard22991 = early_reset_static_par0_go_out;
wire _guard22992 = _guard22990 & _guard22991;
wire _guard22993 = ~_guard0;
wire _guard22994 = early_reset_static_par0_go_out;
wire _guard22995 = _guard22993 & _guard22994;
wire _guard22996 = early_reset_static_par0_go_out;
wire _guard22997 = ~_guard0;
wire _guard22998 = early_reset_static_par0_go_out;
wire _guard22999 = _guard22997 & _guard22998;
wire _guard23000 = early_reset_static_par0_go_out;
wire _guard23001 = early_reset_static_par0_go_out;
wire _guard23002 = early_reset_static_par0_go_out;
wire _guard23003 = early_reset_static_par0_go_out;
wire _guard23004 = ~_guard0;
wire _guard23005 = early_reset_static_par0_go_out;
wire _guard23006 = _guard23004 & _guard23005;
wire _guard23007 = ~_guard0;
wire _guard23008 = early_reset_static_par0_go_out;
wire _guard23009 = _guard23007 & _guard23008;
wire _guard23010 = early_reset_static_par0_go_out;
wire _guard23011 = early_reset_static_par0_go_out;
wire _guard23012 = early_reset_static_par0_go_out;
wire _guard23013 = early_reset_static_par0_go_out;
wire _guard23014 = early_reset_static_par0_go_out;
wire _guard23015 = early_reset_static_par0_go_out;
wire _guard23016 = early_reset_static_par0_go_out;
wire _guard23017 = early_reset_static_par0_go_out;
wire _guard23018 = ~_guard0;
wire _guard23019 = early_reset_static_par0_go_out;
wire _guard23020 = _guard23018 & _guard23019;
wire _guard23021 = ~_guard0;
wire _guard23022 = early_reset_static_par0_go_out;
wire _guard23023 = _guard23021 & _guard23022;
wire _guard23024 = early_reset_static_par0_go_out;
wire _guard23025 = early_reset_static_par0_go_out;
wire _guard23026 = early_reset_static_par0_go_out;
wire _guard23027 = early_reset_static_par0_go_out;
wire _guard23028 = early_reset_static_par0_go_out;
wire _guard23029 = early_reset_static_par0_go_out;
wire _guard23030 = early_reset_static_par0_go_out;
wire _guard23031 = ~_guard0;
wire _guard23032 = early_reset_static_par0_go_out;
wire _guard23033 = _guard23031 & _guard23032;
wire _guard23034 = early_reset_static_par0_go_out;
wire _guard23035 = early_reset_static_par0_go_out;
wire _guard23036 = ~_guard0;
wire _guard23037 = early_reset_static_par0_go_out;
wire _guard23038 = _guard23036 & _guard23037;
wire _guard23039 = ~_guard0;
wire _guard23040 = early_reset_static_par0_go_out;
wire _guard23041 = _guard23039 & _guard23040;
wire _guard23042 = early_reset_static_par0_go_out;
wire _guard23043 = ~_guard0;
wire _guard23044 = early_reset_static_par0_go_out;
wire _guard23045 = _guard23043 & _guard23044;
wire _guard23046 = early_reset_static_par0_go_out;
wire _guard23047 = ~_guard0;
wire _guard23048 = early_reset_static_par0_go_out;
wire _guard23049 = _guard23047 & _guard23048;
wire _guard23050 = early_reset_static_par0_go_out;
wire _guard23051 = early_reset_static_par0_go_out;
wire _guard23052 = early_reset_static_par0_go_out;
wire _guard23053 = early_reset_static_par0_go_out;
wire _guard23054 = early_reset_static_par0_go_out;
wire _guard23055 = early_reset_static_par0_go_out;
wire _guard23056 = ~_guard0;
wire _guard23057 = early_reset_static_par0_go_out;
wire _guard23058 = _guard23056 & _guard23057;
wire _guard23059 = early_reset_static_par0_go_out;
wire _guard23060 = early_reset_static_par0_go_out;
wire _guard23061 = ~_guard0;
wire _guard23062 = early_reset_static_par0_go_out;
wire _guard23063 = _guard23061 & _guard23062;
wire _guard23064 = early_reset_static_par0_go_out;
wire _guard23065 = ~_guard0;
wire _guard23066 = early_reset_static_par0_go_out;
wire _guard23067 = _guard23065 & _guard23066;
wire _guard23068 = early_reset_static_par0_go_out;
wire _guard23069 = early_reset_static_par0_go_out;
wire _guard23070 = ~_guard0;
wire _guard23071 = early_reset_static_par0_go_out;
wire _guard23072 = _guard23070 & _guard23071;
wire _guard23073 = early_reset_static_par0_go_out;
wire _guard23074 = early_reset_static_par0_go_out;
wire _guard23075 = ~_guard0;
wire _guard23076 = early_reset_static_par0_go_out;
wire _guard23077 = _guard23075 & _guard23076;
wire _guard23078 = early_reset_static_par0_go_out;
wire _guard23079 = early_reset_static_par0_go_out;
wire _guard23080 = ~_guard0;
wire _guard23081 = early_reset_static_par0_go_out;
wire _guard23082 = _guard23080 & _guard23081;
wire _guard23083 = early_reset_static_par0_go_out;
wire _guard23084 = early_reset_static_par0_go_out;
wire _guard23085 = early_reset_static_par0_go_out;
wire _guard23086 = early_reset_static_par0_go_out;
wire _guard23087 = early_reset_static_par0_go_out;
wire _guard23088 = early_reset_static_par0_go_out;
wire _guard23089 = early_reset_static_par0_go_out;
wire _guard23090 = early_reset_static_par0_go_out;
wire _guard23091 = early_reset_static_par0_go_out;
wire _guard23092 = ~_guard0;
wire _guard23093 = early_reset_static_par0_go_out;
wire _guard23094 = _guard23092 & _guard23093;
wire _guard23095 = ~_guard0;
wire _guard23096 = early_reset_static_par0_go_out;
wire _guard23097 = _guard23095 & _guard23096;
wire _guard23098 = early_reset_static_par0_go_out;
wire _guard23099 = ~_guard0;
wire _guard23100 = early_reset_static_par0_go_out;
wire _guard23101 = _guard23099 & _guard23100;
wire _guard23102 = early_reset_static_par0_go_out;
wire _guard23103 = ~_guard0;
wire _guard23104 = early_reset_static_par0_go_out;
wire _guard23105 = _guard23103 & _guard23104;
wire _guard23106 = early_reset_static_par0_go_out;
wire _guard23107 = early_reset_static_par0_go_out;
wire _guard23108 = early_reset_static_par0_go_out;
wire _guard23109 = ~_guard0;
wire _guard23110 = early_reset_static_par0_go_out;
wire _guard23111 = _guard23109 & _guard23110;
wire _guard23112 = early_reset_static_par0_go_out;
wire _guard23113 = early_reset_static_par0_go_out;
wire _guard23114 = early_reset_static_par0_go_out;
wire _guard23115 = early_reset_static_par0_go_out;
wire _guard23116 = early_reset_static_par0_go_out;
wire _guard23117 = early_reset_static_par0_go_out;
wire _guard23118 = early_reset_static_par0_go_out;
wire _guard23119 = ~_guard0;
wire _guard23120 = early_reset_static_par0_go_out;
wire _guard23121 = _guard23119 & _guard23120;
wire _guard23122 = early_reset_static_par0_go_out;
wire _guard23123 = early_reset_static_par0_go_out;
wire _guard23124 = early_reset_static_par0_go_out;
wire _guard23125 = ~_guard0;
wire _guard23126 = early_reset_static_par0_go_out;
wire _guard23127 = _guard23125 & _guard23126;
wire _guard23128 = early_reset_static_par0_go_out;
wire _guard23129 = early_reset_static_par0_go_out;
wire _guard23130 = ~_guard0;
wire _guard23131 = early_reset_static_par0_go_out;
wire _guard23132 = _guard23130 & _guard23131;
wire _guard23133 = early_reset_static_par0_go_out;
wire _guard23134 = ~_guard0;
wire _guard23135 = early_reset_static_par0_go_out;
wire _guard23136 = _guard23134 & _guard23135;
wire _guard23137 = early_reset_static_par0_go_out;
wire _guard23138 = early_reset_static_par0_go_out;
wire _guard23139 = early_reset_static_par0_go_out;
wire _guard23140 = ~_guard0;
wire _guard23141 = early_reset_static_par0_go_out;
wire _guard23142 = _guard23140 & _guard23141;
wire _guard23143 = early_reset_static_par0_go_out;
wire _guard23144 = early_reset_static_par0_go_out;
wire _guard23145 = early_reset_static_par0_go_out;
wire _guard23146 = early_reset_static_par0_go_out;
wire _guard23147 = early_reset_static_par0_go_out;
wire _guard23148 = early_reset_static_par0_go_out;
wire _guard23149 = early_reset_static_par0_go_out;
wire _guard23150 = ~_guard0;
wire _guard23151 = early_reset_static_par0_go_out;
wire _guard23152 = _guard23150 & _guard23151;
wire _guard23153 = cond_wire_out;
wire _guard23154 = early_reset_static_par0_go_out;
wire _guard23155 = _guard23153 & _guard23154;
wire _guard23156 = cond_wire_out;
wire _guard23157 = early_reset_static_par0_go_out;
wire _guard23158 = _guard23156 & _guard23157;
wire _guard23159 = cond_wire24_out;
wire _guard23160 = early_reset_static_par0_go_out;
wire _guard23161 = _guard23159 & _guard23160;
wire _guard23162 = cond_wire24_out;
wire _guard23163 = early_reset_static_par0_go_out;
wire _guard23164 = _guard23162 & _guard23163;
wire _guard23165 = cond_wire39_out;
wire _guard23166 = early_reset_static_par0_go_out;
wire _guard23167 = _guard23165 & _guard23166;
wire _guard23168 = cond_wire39_out;
wire _guard23169 = early_reset_static_par0_go_out;
wire _guard23170 = _guard23168 & _guard23169;
wire _guard23171 = cond_wire86_out;
wire _guard23172 = early_reset_static_par0_go_out;
wire _guard23173 = _guard23171 & _guard23172;
wire _guard23174 = cond_wire84_out;
wire _guard23175 = early_reset_static_par0_go_out;
wire _guard23176 = _guard23174 & _guard23175;
wire _guard23177 = fsm_out == 1'd0;
wire _guard23178 = cond_wire84_out;
wire _guard23179 = _guard23177 & _guard23178;
wire _guard23180 = fsm_out == 1'd0;
wire _guard23181 = _guard23179 & _guard23180;
wire _guard23182 = fsm_out == 1'd0;
wire _guard23183 = cond_wire86_out;
wire _guard23184 = _guard23182 & _guard23183;
wire _guard23185 = fsm_out == 1'd0;
wire _guard23186 = _guard23184 & _guard23185;
wire _guard23187 = _guard23181 | _guard23186;
wire _guard23188 = early_reset_static_par0_go_out;
wire _guard23189 = _guard23187 & _guard23188;
wire _guard23190 = fsm_out == 1'd0;
wire _guard23191 = cond_wire84_out;
wire _guard23192 = _guard23190 & _guard23191;
wire _guard23193 = fsm_out == 1'd0;
wire _guard23194 = _guard23192 & _guard23193;
wire _guard23195 = fsm_out == 1'd0;
wire _guard23196 = cond_wire86_out;
wire _guard23197 = _guard23195 & _guard23196;
wire _guard23198 = fsm_out == 1'd0;
wire _guard23199 = _guard23197 & _guard23198;
wire _guard23200 = _guard23194 | _guard23199;
wire _guard23201 = early_reset_static_par0_go_out;
wire _guard23202 = _guard23200 & _guard23201;
wire _guard23203 = fsm_out == 1'd0;
wire _guard23204 = cond_wire84_out;
wire _guard23205 = _guard23203 & _guard23204;
wire _guard23206 = fsm_out == 1'd0;
wire _guard23207 = _guard23205 & _guard23206;
wire _guard23208 = fsm_out == 1'd0;
wire _guard23209 = cond_wire86_out;
wire _guard23210 = _guard23208 & _guard23209;
wire _guard23211 = fsm_out == 1'd0;
wire _guard23212 = _guard23210 & _guard23211;
wire _guard23213 = _guard23207 | _guard23212;
wire _guard23214 = early_reset_static_par0_go_out;
wire _guard23215 = _guard23213 & _guard23214;
wire _guard23216 = cond_wire46_out;
wire _guard23217 = early_reset_static_par0_go_out;
wire _guard23218 = _guard23216 & _guard23217;
wire _guard23219 = cond_wire46_out;
wire _guard23220 = early_reset_static_par0_go_out;
wire _guard23221 = _guard23219 & _guard23220;
wire _guard23222 = cond_wire134_out;
wire _guard23223 = early_reset_static_par0_go_out;
wire _guard23224 = _guard23222 & _guard23223;
wire _guard23225 = cond_wire132_out;
wire _guard23226 = early_reset_static_par0_go_out;
wire _guard23227 = _guard23225 & _guard23226;
wire _guard23228 = fsm_out == 1'd0;
wire _guard23229 = cond_wire132_out;
wire _guard23230 = _guard23228 & _guard23229;
wire _guard23231 = fsm_out == 1'd0;
wire _guard23232 = _guard23230 & _guard23231;
wire _guard23233 = fsm_out == 1'd0;
wire _guard23234 = cond_wire134_out;
wire _guard23235 = _guard23233 & _guard23234;
wire _guard23236 = fsm_out == 1'd0;
wire _guard23237 = _guard23235 & _guard23236;
wire _guard23238 = _guard23232 | _guard23237;
wire _guard23239 = early_reset_static_par0_go_out;
wire _guard23240 = _guard23238 & _guard23239;
wire _guard23241 = fsm_out == 1'd0;
wire _guard23242 = cond_wire132_out;
wire _guard23243 = _guard23241 & _guard23242;
wire _guard23244 = fsm_out == 1'd0;
wire _guard23245 = _guard23243 & _guard23244;
wire _guard23246 = fsm_out == 1'd0;
wire _guard23247 = cond_wire134_out;
wire _guard23248 = _guard23246 & _guard23247;
wire _guard23249 = fsm_out == 1'd0;
wire _guard23250 = _guard23248 & _guard23249;
wire _guard23251 = _guard23245 | _guard23250;
wire _guard23252 = early_reset_static_par0_go_out;
wire _guard23253 = _guard23251 & _guard23252;
wire _guard23254 = fsm_out == 1'd0;
wire _guard23255 = cond_wire132_out;
wire _guard23256 = _guard23254 & _guard23255;
wire _guard23257 = fsm_out == 1'd0;
wire _guard23258 = _guard23256 & _guard23257;
wire _guard23259 = fsm_out == 1'd0;
wire _guard23260 = cond_wire134_out;
wire _guard23261 = _guard23259 & _guard23260;
wire _guard23262 = fsm_out == 1'd0;
wire _guard23263 = _guard23261 & _guard23262;
wire _guard23264 = _guard23258 | _guard23263;
wire _guard23265 = early_reset_static_par0_go_out;
wire _guard23266 = _guard23264 & _guard23265;
wire _guard23267 = cond_wire109_out;
wire _guard23268 = early_reset_static_par0_go_out;
wire _guard23269 = _guard23267 & _guard23268;
wire _guard23270 = cond_wire109_out;
wire _guard23271 = early_reset_static_par0_go_out;
wire _guard23272 = _guard23270 & _guard23271;
wire _guard23273 = cond_wire186_out;
wire _guard23274 = early_reset_static_par0_go_out;
wire _guard23275 = _guard23273 & _guard23274;
wire _guard23276 = cond_wire186_out;
wire _guard23277 = early_reset_static_par0_go_out;
wire _guard23278 = _guard23276 & _guard23277;
wire _guard23279 = cond_wire137_out;
wire _guard23280 = early_reset_static_par0_go_out;
wire _guard23281 = _guard23279 & _guard23280;
wire _guard23282 = cond_wire137_out;
wire _guard23283 = early_reset_static_par0_go_out;
wire _guard23284 = _guard23282 & _guard23283;
wire _guard23285 = cond_wire198_out;
wire _guard23286 = early_reset_static_par0_go_out;
wire _guard23287 = _guard23285 & _guard23286;
wire _guard23288 = cond_wire198_out;
wire _guard23289 = early_reset_static_par0_go_out;
wire _guard23290 = _guard23288 & _guard23289;
wire _guard23291 = cond_wire316_out;
wire _guard23292 = early_reset_static_par0_go_out;
wire _guard23293 = _guard23291 & _guard23292;
wire _guard23294 = cond_wire316_out;
wire _guard23295 = early_reset_static_par0_go_out;
wire _guard23296 = _guard23294 & _guard23295;
wire _guard23297 = cond_wire345_out;
wire _guard23298 = early_reset_static_par0_go_out;
wire _guard23299 = _guard23297 & _guard23298;
wire _guard23300 = cond_wire345_out;
wire _guard23301 = early_reset_static_par0_go_out;
wire _guard23302 = _guard23300 & _guard23301;
wire _guard23303 = cond_wire304_out;
wire _guard23304 = early_reset_static_par0_go_out;
wire _guard23305 = _guard23303 & _guard23304;
wire _guard23306 = cond_wire304_out;
wire _guard23307 = early_reset_static_par0_go_out;
wire _guard23308 = _guard23306 & _guard23307;
wire _guard23309 = cond_wire365_out;
wire _guard23310 = early_reset_static_par0_go_out;
wire _guard23311 = _guard23309 & _guard23310;
wire _guard23312 = cond_wire365_out;
wire _guard23313 = early_reset_static_par0_go_out;
wire _guard23314 = _guard23312 & _guard23313;
wire _guard23315 = cond_wire404_out;
wire _guard23316 = early_reset_static_par0_go_out;
wire _guard23317 = _guard23315 & _guard23316;
wire _guard23318 = cond_wire404_out;
wire _guard23319 = early_reset_static_par0_go_out;
wire _guard23320 = _guard23318 & _guard23319;
wire _guard23321 = cond_wire439_out;
wire _guard23322 = early_reset_static_par0_go_out;
wire _guard23323 = _guard23321 & _guard23322;
wire _guard23324 = cond_wire437_out;
wire _guard23325 = early_reset_static_par0_go_out;
wire _guard23326 = _guard23324 & _guard23325;
wire _guard23327 = fsm_out == 1'd0;
wire _guard23328 = cond_wire437_out;
wire _guard23329 = _guard23327 & _guard23328;
wire _guard23330 = fsm_out == 1'd0;
wire _guard23331 = _guard23329 & _guard23330;
wire _guard23332 = fsm_out == 1'd0;
wire _guard23333 = cond_wire439_out;
wire _guard23334 = _guard23332 & _guard23333;
wire _guard23335 = fsm_out == 1'd0;
wire _guard23336 = _guard23334 & _guard23335;
wire _guard23337 = _guard23331 | _guard23336;
wire _guard23338 = early_reset_static_par0_go_out;
wire _guard23339 = _guard23337 & _guard23338;
wire _guard23340 = fsm_out == 1'd0;
wire _guard23341 = cond_wire437_out;
wire _guard23342 = _guard23340 & _guard23341;
wire _guard23343 = fsm_out == 1'd0;
wire _guard23344 = _guard23342 & _guard23343;
wire _guard23345 = fsm_out == 1'd0;
wire _guard23346 = cond_wire439_out;
wire _guard23347 = _guard23345 & _guard23346;
wire _guard23348 = fsm_out == 1'd0;
wire _guard23349 = _guard23347 & _guard23348;
wire _guard23350 = _guard23344 | _guard23349;
wire _guard23351 = early_reset_static_par0_go_out;
wire _guard23352 = _guard23350 & _guard23351;
wire _guard23353 = fsm_out == 1'd0;
wire _guard23354 = cond_wire437_out;
wire _guard23355 = _guard23353 & _guard23354;
wire _guard23356 = fsm_out == 1'd0;
wire _guard23357 = _guard23355 & _guard23356;
wire _guard23358 = fsm_out == 1'd0;
wire _guard23359 = cond_wire439_out;
wire _guard23360 = _guard23358 & _guard23359;
wire _guard23361 = fsm_out == 1'd0;
wire _guard23362 = _guard23360 & _guard23361;
wire _guard23363 = _guard23357 | _guard23362;
wire _guard23364 = early_reset_static_par0_go_out;
wire _guard23365 = _guard23363 & _guard23364;
wire _guard23366 = cond_wire410_out;
wire _guard23367 = early_reset_static_par0_go_out;
wire _guard23368 = _guard23366 & _guard23367;
wire _guard23369 = cond_wire410_out;
wire _guard23370 = early_reset_static_par0_go_out;
wire _guard23371 = _guard23369 & _guard23370;
wire _guard23372 = cond_wire504_out;
wire _guard23373 = early_reset_static_par0_go_out;
wire _guard23374 = _guard23372 & _guard23373;
wire _guard23375 = cond_wire502_out;
wire _guard23376 = early_reset_static_par0_go_out;
wire _guard23377 = _guard23375 & _guard23376;
wire _guard23378 = fsm_out == 1'd0;
wire _guard23379 = cond_wire502_out;
wire _guard23380 = _guard23378 & _guard23379;
wire _guard23381 = fsm_out == 1'd0;
wire _guard23382 = _guard23380 & _guard23381;
wire _guard23383 = fsm_out == 1'd0;
wire _guard23384 = cond_wire504_out;
wire _guard23385 = _guard23383 & _guard23384;
wire _guard23386 = fsm_out == 1'd0;
wire _guard23387 = _guard23385 & _guard23386;
wire _guard23388 = _guard23382 | _guard23387;
wire _guard23389 = early_reset_static_par0_go_out;
wire _guard23390 = _guard23388 & _guard23389;
wire _guard23391 = fsm_out == 1'd0;
wire _guard23392 = cond_wire502_out;
wire _guard23393 = _guard23391 & _guard23392;
wire _guard23394 = fsm_out == 1'd0;
wire _guard23395 = _guard23393 & _guard23394;
wire _guard23396 = fsm_out == 1'd0;
wire _guard23397 = cond_wire504_out;
wire _guard23398 = _guard23396 & _guard23397;
wire _guard23399 = fsm_out == 1'd0;
wire _guard23400 = _guard23398 & _guard23399;
wire _guard23401 = _guard23395 | _guard23400;
wire _guard23402 = early_reset_static_par0_go_out;
wire _guard23403 = _guard23401 & _guard23402;
wire _guard23404 = fsm_out == 1'd0;
wire _guard23405 = cond_wire502_out;
wire _guard23406 = _guard23404 & _guard23405;
wire _guard23407 = fsm_out == 1'd0;
wire _guard23408 = _guard23406 & _guard23407;
wire _guard23409 = fsm_out == 1'd0;
wire _guard23410 = cond_wire504_out;
wire _guard23411 = _guard23409 & _guard23410;
wire _guard23412 = fsm_out == 1'd0;
wire _guard23413 = _guard23411 & _guard23412;
wire _guard23414 = _guard23408 | _guard23413;
wire _guard23415 = early_reset_static_par0_go_out;
wire _guard23416 = _guard23414 & _guard23415;
wire _guard23417 = cond_wire516_out;
wire _guard23418 = early_reset_static_par0_go_out;
wire _guard23419 = _guard23417 & _guard23418;
wire _guard23420 = cond_wire514_out;
wire _guard23421 = early_reset_static_par0_go_out;
wire _guard23422 = _guard23420 & _guard23421;
wire _guard23423 = fsm_out == 1'd0;
wire _guard23424 = cond_wire514_out;
wire _guard23425 = _guard23423 & _guard23424;
wire _guard23426 = fsm_out == 1'd0;
wire _guard23427 = _guard23425 & _guard23426;
wire _guard23428 = fsm_out == 1'd0;
wire _guard23429 = cond_wire516_out;
wire _guard23430 = _guard23428 & _guard23429;
wire _guard23431 = fsm_out == 1'd0;
wire _guard23432 = _guard23430 & _guard23431;
wire _guard23433 = _guard23427 | _guard23432;
wire _guard23434 = early_reset_static_par0_go_out;
wire _guard23435 = _guard23433 & _guard23434;
wire _guard23436 = fsm_out == 1'd0;
wire _guard23437 = cond_wire514_out;
wire _guard23438 = _guard23436 & _guard23437;
wire _guard23439 = fsm_out == 1'd0;
wire _guard23440 = _guard23438 & _guard23439;
wire _guard23441 = fsm_out == 1'd0;
wire _guard23442 = cond_wire516_out;
wire _guard23443 = _guard23441 & _guard23442;
wire _guard23444 = fsm_out == 1'd0;
wire _guard23445 = _guard23443 & _guard23444;
wire _guard23446 = _guard23440 | _guard23445;
wire _guard23447 = early_reset_static_par0_go_out;
wire _guard23448 = _guard23446 & _guard23447;
wire _guard23449 = fsm_out == 1'd0;
wire _guard23450 = cond_wire514_out;
wire _guard23451 = _guard23449 & _guard23450;
wire _guard23452 = fsm_out == 1'd0;
wire _guard23453 = _guard23451 & _guard23452;
wire _guard23454 = fsm_out == 1'd0;
wire _guard23455 = cond_wire516_out;
wire _guard23456 = _guard23454 & _guard23455;
wire _guard23457 = fsm_out == 1'd0;
wire _guard23458 = _guard23456 & _guard23457;
wire _guard23459 = _guard23453 | _guard23458;
wire _guard23460 = early_reset_static_par0_go_out;
wire _guard23461 = _guard23459 & _guard23460;
wire _guard23462 = cond_wire524_out;
wire _guard23463 = early_reset_static_par0_go_out;
wire _guard23464 = _guard23462 & _guard23463;
wire _guard23465 = cond_wire522_out;
wire _guard23466 = early_reset_static_par0_go_out;
wire _guard23467 = _guard23465 & _guard23466;
wire _guard23468 = fsm_out == 1'd0;
wire _guard23469 = cond_wire522_out;
wire _guard23470 = _guard23468 & _guard23469;
wire _guard23471 = fsm_out == 1'd0;
wire _guard23472 = _guard23470 & _guard23471;
wire _guard23473 = fsm_out == 1'd0;
wire _guard23474 = cond_wire524_out;
wire _guard23475 = _guard23473 & _guard23474;
wire _guard23476 = fsm_out == 1'd0;
wire _guard23477 = _guard23475 & _guard23476;
wire _guard23478 = _guard23472 | _guard23477;
wire _guard23479 = early_reset_static_par0_go_out;
wire _guard23480 = _guard23478 & _guard23479;
wire _guard23481 = fsm_out == 1'd0;
wire _guard23482 = cond_wire522_out;
wire _guard23483 = _guard23481 & _guard23482;
wire _guard23484 = fsm_out == 1'd0;
wire _guard23485 = _guard23483 & _guard23484;
wire _guard23486 = fsm_out == 1'd0;
wire _guard23487 = cond_wire524_out;
wire _guard23488 = _guard23486 & _guard23487;
wire _guard23489 = fsm_out == 1'd0;
wire _guard23490 = _guard23488 & _guard23489;
wire _guard23491 = _guard23485 | _guard23490;
wire _guard23492 = early_reset_static_par0_go_out;
wire _guard23493 = _guard23491 & _guard23492;
wire _guard23494 = fsm_out == 1'd0;
wire _guard23495 = cond_wire522_out;
wire _guard23496 = _guard23494 & _guard23495;
wire _guard23497 = fsm_out == 1'd0;
wire _guard23498 = _guard23496 & _guard23497;
wire _guard23499 = fsm_out == 1'd0;
wire _guard23500 = cond_wire524_out;
wire _guard23501 = _guard23499 & _guard23500;
wire _guard23502 = fsm_out == 1'd0;
wire _guard23503 = _guard23501 & _guard23502;
wire _guard23504 = _guard23498 | _guard23503;
wire _guard23505 = early_reset_static_par0_go_out;
wire _guard23506 = _guard23504 & _guard23505;
wire _guard23507 = cond_wire458_out;
wire _guard23508 = early_reset_static_par0_go_out;
wire _guard23509 = _guard23507 & _guard23508;
wire _guard23510 = cond_wire458_out;
wire _guard23511 = early_reset_static_par0_go_out;
wire _guard23512 = _guard23510 & _guard23511;
wire _guard23513 = cond_wire527_out;
wire _guard23514 = early_reset_static_par0_go_out;
wire _guard23515 = _guard23513 & _guard23514;
wire _guard23516 = cond_wire527_out;
wire _guard23517 = early_reset_static_par0_go_out;
wire _guard23518 = _guard23516 & _guard23517;
wire _guard23519 = cond_wire491_out;
wire _guard23520 = early_reset_static_par0_go_out;
wire _guard23521 = _guard23519 & _guard23520;
wire _guard23522 = cond_wire491_out;
wire _guard23523 = early_reset_static_par0_go_out;
wire _guard23524 = _guard23522 & _guard23523;
wire _guard23525 = cond_wire507_out;
wire _guard23526 = early_reset_static_par0_go_out;
wire _guard23527 = _guard23525 & _guard23526;
wire _guard23528 = cond_wire507_out;
wire _guard23529 = early_reset_static_par0_go_out;
wire _guard23530 = _guard23528 & _guard23529;
wire _guard23531 = cond_wire610_out;
wire _guard23532 = early_reset_static_par0_go_out;
wire _guard23533 = _guard23531 & _guard23532;
wire _guard23534 = cond_wire608_out;
wire _guard23535 = early_reset_static_par0_go_out;
wire _guard23536 = _guard23534 & _guard23535;
wire _guard23537 = fsm_out == 1'd0;
wire _guard23538 = cond_wire608_out;
wire _guard23539 = _guard23537 & _guard23538;
wire _guard23540 = fsm_out == 1'd0;
wire _guard23541 = _guard23539 & _guard23540;
wire _guard23542 = fsm_out == 1'd0;
wire _guard23543 = cond_wire610_out;
wire _guard23544 = _guard23542 & _guard23543;
wire _guard23545 = fsm_out == 1'd0;
wire _guard23546 = _guard23544 & _guard23545;
wire _guard23547 = _guard23541 | _guard23546;
wire _guard23548 = early_reset_static_par0_go_out;
wire _guard23549 = _guard23547 & _guard23548;
wire _guard23550 = fsm_out == 1'd0;
wire _guard23551 = cond_wire608_out;
wire _guard23552 = _guard23550 & _guard23551;
wire _guard23553 = fsm_out == 1'd0;
wire _guard23554 = _guard23552 & _guard23553;
wire _guard23555 = fsm_out == 1'd0;
wire _guard23556 = cond_wire610_out;
wire _guard23557 = _guard23555 & _guard23556;
wire _guard23558 = fsm_out == 1'd0;
wire _guard23559 = _guard23557 & _guard23558;
wire _guard23560 = _guard23554 | _guard23559;
wire _guard23561 = early_reset_static_par0_go_out;
wire _guard23562 = _guard23560 & _guard23561;
wire _guard23563 = fsm_out == 1'd0;
wire _guard23564 = cond_wire608_out;
wire _guard23565 = _guard23563 & _guard23564;
wire _guard23566 = fsm_out == 1'd0;
wire _guard23567 = _guard23565 & _guard23566;
wire _guard23568 = fsm_out == 1'd0;
wire _guard23569 = cond_wire610_out;
wire _guard23570 = _guard23568 & _guard23569;
wire _guard23571 = fsm_out == 1'd0;
wire _guard23572 = _guard23570 & _guard23571;
wire _guard23573 = _guard23567 | _guard23572;
wire _guard23574 = early_reset_static_par0_go_out;
wire _guard23575 = _guard23573 & _guard23574;
wire _guard23576 = cond_wire609_out;
wire _guard23577 = early_reset_static_par0_go_out;
wire _guard23578 = _guard23576 & _guard23577;
wire _guard23579 = cond_wire609_out;
wire _guard23580 = early_reset_static_par0_go_out;
wire _guard23581 = _guard23579 & _guard23580;
wire _guard23582 = cond_wire564_out;
wire _guard23583 = early_reset_static_par0_go_out;
wire _guard23584 = _guard23582 & _guard23583;
wire _guard23585 = cond_wire564_out;
wire _guard23586 = early_reset_static_par0_go_out;
wire _guard23587 = _guard23585 & _guard23586;
wire _guard23588 = cond_wire576_out;
wire _guard23589 = early_reset_static_par0_go_out;
wire _guard23590 = _guard23588 & _guard23589;
wire _guard23591 = cond_wire576_out;
wire _guard23592 = early_reset_static_par0_go_out;
wire _guard23593 = _guard23591 & _guard23592;
wire _guard23594 = cond_wire588_out;
wire _guard23595 = early_reset_static_par0_go_out;
wire _guard23596 = _guard23594 & _guard23595;
wire _guard23597 = cond_wire588_out;
wire _guard23598 = early_reset_static_par0_go_out;
wire _guard23599 = _guard23597 & _guard23598;
wire _guard23600 = cond_wire671_out;
wire _guard23601 = early_reset_static_par0_go_out;
wire _guard23602 = _guard23600 & _guard23601;
wire _guard23603 = cond_wire669_out;
wire _guard23604 = early_reset_static_par0_go_out;
wire _guard23605 = _guard23603 & _guard23604;
wire _guard23606 = fsm_out == 1'd0;
wire _guard23607 = cond_wire669_out;
wire _guard23608 = _guard23606 & _guard23607;
wire _guard23609 = fsm_out == 1'd0;
wire _guard23610 = _guard23608 & _guard23609;
wire _guard23611 = fsm_out == 1'd0;
wire _guard23612 = cond_wire671_out;
wire _guard23613 = _guard23611 & _guard23612;
wire _guard23614 = fsm_out == 1'd0;
wire _guard23615 = _guard23613 & _guard23614;
wire _guard23616 = _guard23610 | _guard23615;
wire _guard23617 = early_reset_static_par0_go_out;
wire _guard23618 = _guard23616 & _guard23617;
wire _guard23619 = fsm_out == 1'd0;
wire _guard23620 = cond_wire669_out;
wire _guard23621 = _guard23619 & _guard23620;
wire _guard23622 = fsm_out == 1'd0;
wire _guard23623 = _guard23621 & _guard23622;
wire _guard23624 = fsm_out == 1'd0;
wire _guard23625 = cond_wire671_out;
wire _guard23626 = _guard23624 & _guard23625;
wire _guard23627 = fsm_out == 1'd0;
wire _guard23628 = _guard23626 & _guard23627;
wire _guard23629 = _guard23623 | _guard23628;
wire _guard23630 = early_reset_static_par0_go_out;
wire _guard23631 = _guard23629 & _guard23630;
wire _guard23632 = fsm_out == 1'd0;
wire _guard23633 = cond_wire669_out;
wire _guard23634 = _guard23632 & _guard23633;
wire _guard23635 = fsm_out == 1'd0;
wire _guard23636 = _guard23634 & _guard23635;
wire _guard23637 = fsm_out == 1'd0;
wire _guard23638 = cond_wire671_out;
wire _guard23639 = _guard23637 & _guard23638;
wire _guard23640 = fsm_out == 1'd0;
wire _guard23641 = _guard23639 & _guard23640;
wire _guard23642 = _guard23636 | _guard23641;
wire _guard23643 = early_reset_static_par0_go_out;
wire _guard23644 = _guard23642 & _guard23643;
wire _guard23645 = cond_wire613_out;
wire _guard23646 = early_reset_static_par0_go_out;
wire _guard23647 = _guard23645 & _guard23646;
wire _guard23648 = cond_wire613_out;
wire _guard23649 = early_reset_static_par0_go_out;
wire _guard23650 = _guard23648 & _guard23649;
wire _guard23651 = cond_wire691_out;
wire _guard23652 = early_reset_static_par0_go_out;
wire _guard23653 = _guard23651 & _guard23652;
wire _guard23654 = cond_wire689_out;
wire _guard23655 = early_reset_static_par0_go_out;
wire _guard23656 = _guard23654 & _guard23655;
wire _guard23657 = fsm_out == 1'd0;
wire _guard23658 = cond_wire689_out;
wire _guard23659 = _guard23657 & _guard23658;
wire _guard23660 = fsm_out == 1'd0;
wire _guard23661 = _guard23659 & _guard23660;
wire _guard23662 = fsm_out == 1'd0;
wire _guard23663 = cond_wire691_out;
wire _guard23664 = _guard23662 & _guard23663;
wire _guard23665 = fsm_out == 1'd0;
wire _guard23666 = _guard23664 & _guard23665;
wire _guard23667 = _guard23661 | _guard23666;
wire _guard23668 = early_reset_static_par0_go_out;
wire _guard23669 = _guard23667 & _guard23668;
wire _guard23670 = fsm_out == 1'd0;
wire _guard23671 = cond_wire689_out;
wire _guard23672 = _guard23670 & _guard23671;
wire _guard23673 = fsm_out == 1'd0;
wire _guard23674 = _guard23672 & _guard23673;
wire _guard23675 = fsm_out == 1'd0;
wire _guard23676 = cond_wire691_out;
wire _guard23677 = _guard23675 & _guard23676;
wire _guard23678 = fsm_out == 1'd0;
wire _guard23679 = _guard23677 & _guard23678;
wire _guard23680 = _guard23674 | _guard23679;
wire _guard23681 = early_reset_static_par0_go_out;
wire _guard23682 = _guard23680 & _guard23681;
wire _guard23683 = fsm_out == 1'd0;
wire _guard23684 = cond_wire689_out;
wire _guard23685 = _guard23683 & _guard23684;
wire _guard23686 = fsm_out == 1'd0;
wire _guard23687 = _guard23685 & _guard23686;
wire _guard23688 = fsm_out == 1'd0;
wire _guard23689 = cond_wire691_out;
wire _guard23690 = _guard23688 & _guard23689;
wire _guard23691 = fsm_out == 1'd0;
wire _guard23692 = _guard23690 & _guard23691;
wire _guard23693 = _guard23687 | _guard23692;
wire _guard23694 = early_reset_static_par0_go_out;
wire _guard23695 = _guard23693 & _guard23694;
wire _guard23696 = cond_wire649_out;
wire _guard23697 = early_reset_static_par0_go_out;
wire _guard23698 = _guard23696 & _guard23697;
wire _guard23699 = cond_wire649_out;
wire _guard23700 = early_reset_static_par0_go_out;
wire _guard23701 = _guard23699 & _guard23700;
wire _guard23702 = cond_wire755_out;
wire _guard23703 = early_reset_static_par0_go_out;
wire _guard23704 = _guard23702 & _guard23703;
wire _guard23705 = cond_wire755_out;
wire _guard23706 = early_reset_static_par0_go_out;
wire _guard23707 = _guard23705 & _guard23706;
wire _guard23708 = cond_wire714_out;
wire _guard23709 = early_reset_static_par0_go_out;
wire _guard23710 = _guard23708 & _guard23709;
wire _guard23711 = cond_wire714_out;
wire _guard23712 = early_reset_static_par0_go_out;
wire _guard23713 = _guard23711 & _guard23712;
wire _guard23714 = cond_wire779_out;
wire _guard23715 = early_reset_static_par0_go_out;
wire _guard23716 = _guard23714 & _guard23715;
wire _guard23717 = cond_wire779_out;
wire _guard23718 = early_reset_static_par0_go_out;
wire _guard23719 = _guard23717 & _guard23718;
wire _guard23720 = cond_wire797_out;
wire _guard23721 = early_reset_static_par0_go_out;
wire _guard23722 = _guard23720 & _guard23721;
wire _guard23723 = cond_wire795_out;
wire _guard23724 = early_reset_static_par0_go_out;
wire _guard23725 = _guard23723 & _guard23724;
wire _guard23726 = fsm_out == 1'd0;
wire _guard23727 = cond_wire795_out;
wire _guard23728 = _guard23726 & _guard23727;
wire _guard23729 = fsm_out == 1'd0;
wire _guard23730 = _guard23728 & _guard23729;
wire _guard23731 = fsm_out == 1'd0;
wire _guard23732 = cond_wire797_out;
wire _guard23733 = _guard23731 & _guard23732;
wire _guard23734 = fsm_out == 1'd0;
wire _guard23735 = _guard23733 & _guard23734;
wire _guard23736 = _guard23730 | _guard23735;
wire _guard23737 = early_reset_static_par0_go_out;
wire _guard23738 = _guard23736 & _guard23737;
wire _guard23739 = fsm_out == 1'd0;
wire _guard23740 = cond_wire795_out;
wire _guard23741 = _guard23739 & _guard23740;
wire _guard23742 = fsm_out == 1'd0;
wire _guard23743 = _guard23741 & _guard23742;
wire _guard23744 = fsm_out == 1'd0;
wire _guard23745 = cond_wire797_out;
wire _guard23746 = _guard23744 & _guard23745;
wire _guard23747 = fsm_out == 1'd0;
wire _guard23748 = _guard23746 & _guard23747;
wire _guard23749 = _guard23743 | _guard23748;
wire _guard23750 = early_reset_static_par0_go_out;
wire _guard23751 = _guard23749 & _guard23750;
wire _guard23752 = fsm_out == 1'd0;
wire _guard23753 = cond_wire795_out;
wire _guard23754 = _guard23752 & _guard23753;
wire _guard23755 = fsm_out == 1'd0;
wire _guard23756 = _guard23754 & _guard23755;
wire _guard23757 = fsm_out == 1'd0;
wire _guard23758 = cond_wire797_out;
wire _guard23759 = _guard23757 & _guard23758;
wire _guard23760 = fsm_out == 1'd0;
wire _guard23761 = _guard23759 & _guard23760;
wire _guard23762 = _guard23756 | _guard23761;
wire _guard23763 = early_reset_static_par0_go_out;
wire _guard23764 = _guard23762 & _guard23763;
wire _guard23765 = cond_wire747_out;
wire _guard23766 = early_reset_static_par0_go_out;
wire _guard23767 = _guard23765 & _guard23766;
wire _guard23768 = cond_wire747_out;
wire _guard23769 = early_reset_static_par0_go_out;
wire _guard23770 = _guard23768 & _guard23769;
wire _guard23771 = cond_wire840_out;
wire _guard23772 = early_reset_static_par0_go_out;
wire _guard23773 = _guard23771 & _guard23772;
wire _guard23774 = cond_wire840_out;
wire _guard23775 = early_reset_static_par0_go_out;
wire _guard23776 = _guard23774 & _guard23775;
wire _guard23777 = cond_wire877_out;
wire _guard23778 = early_reset_static_par0_go_out;
wire _guard23779 = _guard23777 & _guard23778;
wire _guard23780 = cond_wire877_out;
wire _guard23781 = early_reset_static_par0_go_out;
wire _guard23782 = _guard23780 & _guard23781;
wire _guard23783 = cond_wire922_out;
wire _guard23784 = early_reset_static_par0_go_out;
wire _guard23785 = _guard23783 & _guard23784;
wire _guard23786 = cond_wire920_out;
wire _guard23787 = early_reset_static_par0_go_out;
wire _guard23788 = _guard23786 & _guard23787;
wire _guard23789 = fsm_out == 1'd0;
wire _guard23790 = cond_wire920_out;
wire _guard23791 = _guard23789 & _guard23790;
wire _guard23792 = fsm_out == 1'd0;
wire _guard23793 = _guard23791 & _guard23792;
wire _guard23794 = fsm_out == 1'd0;
wire _guard23795 = cond_wire922_out;
wire _guard23796 = _guard23794 & _guard23795;
wire _guard23797 = fsm_out == 1'd0;
wire _guard23798 = _guard23796 & _guard23797;
wire _guard23799 = _guard23793 | _guard23798;
wire _guard23800 = early_reset_static_par0_go_out;
wire _guard23801 = _guard23799 & _guard23800;
wire _guard23802 = fsm_out == 1'd0;
wire _guard23803 = cond_wire920_out;
wire _guard23804 = _guard23802 & _guard23803;
wire _guard23805 = fsm_out == 1'd0;
wire _guard23806 = _guard23804 & _guard23805;
wire _guard23807 = fsm_out == 1'd0;
wire _guard23808 = cond_wire922_out;
wire _guard23809 = _guard23807 & _guard23808;
wire _guard23810 = fsm_out == 1'd0;
wire _guard23811 = _guard23809 & _guard23810;
wire _guard23812 = _guard23806 | _guard23811;
wire _guard23813 = early_reset_static_par0_go_out;
wire _guard23814 = _guard23812 & _guard23813;
wire _guard23815 = fsm_out == 1'd0;
wire _guard23816 = cond_wire920_out;
wire _guard23817 = _guard23815 & _guard23816;
wire _guard23818 = fsm_out == 1'd0;
wire _guard23819 = _guard23817 & _guard23818;
wire _guard23820 = fsm_out == 1'd0;
wire _guard23821 = cond_wire922_out;
wire _guard23822 = _guard23820 & _guard23821;
wire _guard23823 = fsm_out == 1'd0;
wire _guard23824 = _guard23822 & _guard23823;
wire _guard23825 = _guard23819 | _guard23824;
wire _guard23826 = early_reset_static_par0_go_out;
wire _guard23827 = _guard23825 & _guard23826;
wire _guard23828 = cond_wire865_out;
wire _guard23829 = early_reset_static_par0_go_out;
wire _guard23830 = _guard23828 & _guard23829;
wire _guard23831 = cond_wire865_out;
wire _guard23832 = early_reset_static_par0_go_out;
wire _guard23833 = _guard23831 & _guard23832;
wire _guard23834 = cond_wire935_out;
wire _guard23835 = early_reset_static_par0_go_out;
wire _guard23836 = _guard23834 & _guard23835;
wire _guard23837 = cond_wire933_out;
wire _guard23838 = early_reset_static_par0_go_out;
wire _guard23839 = _guard23837 & _guard23838;
wire _guard23840 = fsm_out == 1'd0;
wire _guard23841 = cond_wire933_out;
wire _guard23842 = _guard23840 & _guard23841;
wire _guard23843 = fsm_out == 1'd0;
wire _guard23844 = _guard23842 & _guard23843;
wire _guard23845 = fsm_out == 1'd0;
wire _guard23846 = cond_wire935_out;
wire _guard23847 = _guard23845 & _guard23846;
wire _guard23848 = fsm_out == 1'd0;
wire _guard23849 = _guard23847 & _guard23848;
wire _guard23850 = _guard23844 | _guard23849;
wire _guard23851 = early_reset_static_par0_go_out;
wire _guard23852 = _guard23850 & _guard23851;
wire _guard23853 = fsm_out == 1'd0;
wire _guard23854 = cond_wire933_out;
wire _guard23855 = _guard23853 & _guard23854;
wire _guard23856 = fsm_out == 1'd0;
wire _guard23857 = _guard23855 & _guard23856;
wire _guard23858 = fsm_out == 1'd0;
wire _guard23859 = cond_wire935_out;
wire _guard23860 = _guard23858 & _guard23859;
wire _guard23861 = fsm_out == 1'd0;
wire _guard23862 = _guard23860 & _guard23861;
wire _guard23863 = _guard23857 | _guard23862;
wire _guard23864 = early_reset_static_par0_go_out;
wire _guard23865 = _guard23863 & _guard23864;
wire _guard23866 = fsm_out == 1'd0;
wire _guard23867 = cond_wire933_out;
wire _guard23868 = _guard23866 & _guard23867;
wire _guard23869 = fsm_out == 1'd0;
wire _guard23870 = _guard23868 & _guard23869;
wire _guard23871 = fsm_out == 1'd0;
wire _guard23872 = cond_wire935_out;
wire _guard23873 = _guard23871 & _guard23872;
wire _guard23874 = fsm_out == 1'd0;
wire _guard23875 = _guard23873 & _guard23874;
wire _guard23876 = _guard23870 | _guard23875;
wire _guard23877 = early_reset_static_par0_go_out;
wire _guard23878 = _guard23876 & _guard23877;
wire _guard23879 = cond_wire930_out;
wire _guard23880 = early_reset_static_par0_go_out;
wire _guard23881 = _guard23879 & _guard23880;
wire _guard23882 = cond_wire930_out;
wire _guard23883 = early_reset_static_par0_go_out;
wire _guard23884 = _guard23882 & _guard23883;
wire _guard23885 = cond_wire942_out;
wire _guard23886 = early_reset_static_par0_go_out;
wire _guard23887 = _guard23885 & _guard23886;
wire _guard23888 = cond_wire942_out;
wire _guard23889 = early_reset_static_par0_go_out;
wire _guard23890 = _guard23888 & _guard23889;
wire _guard23891 = cond_wire962_out;
wire _guard23892 = early_reset_static_par0_go_out;
wire _guard23893 = _guard23891 & _guard23892;
wire _guard23894 = cond_wire962_out;
wire _guard23895 = early_reset_static_par0_go_out;
wire _guard23896 = _guard23894 & _guard23895;
wire _guard23897 = cond_wire996_out;
wire _guard23898 = early_reset_static_par0_go_out;
wire _guard23899 = _guard23897 & _guard23898;
wire _guard23900 = cond_wire994_out;
wire _guard23901 = early_reset_static_par0_go_out;
wire _guard23902 = _guard23900 & _guard23901;
wire _guard23903 = fsm_out == 1'd0;
wire _guard23904 = cond_wire994_out;
wire _guard23905 = _guard23903 & _guard23904;
wire _guard23906 = fsm_out == 1'd0;
wire _guard23907 = _guard23905 & _guard23906;
wire _guard23908 = fsm_out == 1'd0;
wire _guard23909 = cond_wire996_out;
wire _guard23910 = _guard23908 & _guard23909;
wire _guard23911 = fsm_out == 1'd0;
wire _guard23912 = _guard23910 & _guard23911;
wire _guard23913 = _guard23907 | _guard23912;
wire _guard23914 = early_reset_static_par0_go_out;
wire _guard23915 = _guard23913 & _guard23914;
wire _guard23916 = fsm_out == 1'd0;
wire _guard23917 = cond_wire994_out;
wire _guard23918 = _guard23916 & _guard23917;
wire _guard23919 = fsm_out == 1'd0;
wire _guard23920 = _guard23918 & _guard23919;
wire _guard23921 = fsm_out == 1'd0;
wire _guard23922 = cond_wire996_out;
wire _guard23923 = _guard23921 & _guard23922;
wire _guard23924 = fsm_out == 1'd0;
wire _guard23925 = _guard23923 & _guard23924;
wire _guard23926 = _guard23920 | _guard23925;
wire _guard23927 = early_reset_static_par0_go_out;
wire _guard23928 = _guard23926 & _guard23927;
wire _guard23929 = fsm_out == 1'd0;
wire _guard23930 = cond_wire994_out;
wire _guard23931 = _guard23929 & _guard23930;
wire _guard23932 = fsm_out == 1'd0;
wire _guard23933 = _guard23931 & _guard23932;
wire _guard23934 = fsm_out == 1'd0;
wire _guard23935 = cond_wire996_out;
wire _guard23936 = _guard23934 & _guard23935;
wire _guard23937 = fsm_out == 1'd0;
wire _guard23938 = _guard23936 & _guard23937;
wire _guard23939 = _guard23933 | _guard23938;
wire _guard23940 = early_reset_static_par0_go_out;
wire _guard23941 = _guard23939 & _guard23940;
wire _guard23942 = cond_wire1012_out;
wire _guard23943 = early_reset_static_par0_go_out;
wire _guard23944 = _guard23942 & _guard23943;
wire _guard23945 = cond_wire1010_out;
wire _guard23946 = early_reset_static_par0_go_out;
wire _guard23947 = _guard23945 & _guard23946;
wire _guard23948 = fsm_out == 1'd0;
wire _guard23949 = cond_wire1010_out;
wire _guard23950 = _guard23948 & _guard23949;
wire _guard23951 = fsm_out == 1'd0;
wire _guard23952 = _guard23950 & _guard23951;
wire _guard23953 = fsm_out == 1'd0;
wire _guard23954 = cond_wire1012_out;
wire _guard23955 = _guard23953 & _guard23954;
wire _guard23956 = fsm_out == 1'd0;
wire _guard23957 = _guard23955 & _guard23956;
wire _guard23958 = _guard23952 | _guard23957;
wire _guard23959 = early_reset_static_par0_go_out;
wire _guard23960 = _guard23958 & _guard23959;
wire _guard23961 = fsm_out == 1'd0;
wire _guard23962 = cond_wire1010_out;
wire _guard23963 = _guard23961 & _guard23962;
wire _guard23964 = fsm_out == 1'd0;
wire _guard23965 = _guard23963 & _guard23964;
wire _guard23966 = fsm_out == 1'd0;
wire _guard23967 = cond_wire1012_out;
wire _guard23968 = _guard23966 & _guard23967;
wire _guard23969 = fsm_out == 1'd0;
wire _guard23970 = _guard23968 & _guard23969;
wire _guard23971 = _guard23965 | _guard23970;
wire _guard23972 = early_reset_static_par0_go_out;
wire _guard23973 = _guard23971 & _guard23972;
wire _guard23974 = fsm_out == 1'd0;
wire _guard23975 = cond_wire1010_out;
wire _guard23976 = _guard23974 & _guard23975;
wire _guard23977 = fsm_out == 1'd0;
wire _guard23978 = _guard23976 & _guard23977;
wire _guard23979 = fsm_out == 1'd0;
wire _guard23980 = cond_wire1012_out;
wire _guard23981 = _guard23979 & _guard23980;
wire _guard23982 = fsm_out == 1'd0;
wire _guard23983 = _guard23981 & _guard23982;
wire _guard23984 = _guard23978 | _guard23983;
wire _guard23985 = early_reset_static_par0_go_out;
wire _guard23986 = _guard23984 & _guard23985;
wire _guard23987 = cond_wire1032_out;
wire _guard23988 = early_reset_static_par0_go_out;
wire _guard23989 = _guard23987 & _guard23988;
wire _guard23990 = cond_wire1030_out;
wire _guard23991 = early_reset_static_par0_go_out;
wire _guard23992 = _guard23990 & _guard23991;
wire _guard23993 = fsm_out == 1'd0;
wire _guard23994 = cond_wire1030_out;
wire _guard23995 = _guard23993 & _guard23994;
wire _guard23996 = fsm_out == 1'd0;
wire _guard23997 = _guard23995 & _guard23996;
wire _guard23998 = fsm_out == 1'd0;
wire _guard23999 = cond_wire1032_out;
wire _guard24000 = _guard23998 & _guard23999;
wire _guard24001 = fsm_out == 1'd0;
wire _guard24002 = _guard24000 & _guard24001;
wire _guard24003 = _guard23997 | _guard24002;
wire _guard24004 = early_reset_static_par0_go_out;
wire _guard24005 = _guard24003 & _guard24004;
wire _guard24006 = fsm_out == 1'd0;
wire _guard24007 = cond_wire1030_out;
wire _guard24008 = _guard24006 & _guard24007;
wire _guard24009 = fsm_out == 1'd0;
wire _guard24010 = _guard24008 & _guard24009;
wire _guard24011 = fsm_out == 1'd0;
wire _guard24012 = cond_wire1032_out;
wire _guard24013 = _guard24011 & _guard24012;
wire _guard24014 = fsm_out == 1'd0;
wire _guard24015 = _guard24013 & _guard24014;
wire _guard24016 = _guard24010 | _guard24015;
wire _guard24017 = early_reset_static_par0_go_out;
wire _guard24018 = _guard24016 & _guard24017;
wire _guard24019 = fsm_out == 1'd0;
wire _guard24020 = cond_wire1030_out;
wire _guard24021 = _guard24019 & _guard24020;
wire _guard24022 = fsm_out == 1'd0;
wire _guard24023 = _guard24021 & _guard24022;
wire _guard24024 = fsm_out == 1'd0;
wire _guard24025 = cond_wire1032_out;
wire _guard24026 = _guard24024 & _guard24025;
wire _guard24027 = fsm_out == 1'd0;
wire _guard24028 = _guard24026 & _guard24027;
wire _guard24029 = _guard24023 | _guard24028;
wire _guard24030 = early_reset_static_par0_go_out;
wire _guard24031 = _guard24029 & _guard24030;
wire _guard24032 = cond_wire978_out;
wire _guard24033 = early_reset_static_par0_go_out;
wire _guard24034 = _guard24032 & _guard24033;
wire _guard24035 = cond_wire978_out;
wire _guard24036 = early_reset_static_par0_go_out;
wire _guard24037 = _guard24035 & _guard24036;
wire _guard24038 = cond_wire986_out;
wire _guard24039 = early_reset_static_par0_go_out;
wire _guard24040 = _guard24038 & _guard24039;
wire _guard24041 = cond_wire986_out;
wire _guard24042 = early_reset_static_par0_go_out;
wire _guard24043 = _guard24041 & _guard24042;
wire _guard24044 = cond_wire1047_out;
wire _guard24045 = early_reset_static_par0_go_out;
wire _guard24046 = _guard24044 & _guard24045;
wire _guard24047 = cond_wire1047_out;
wire _guard24048 = early_reset_static_par0_go_out;
wire _guard24049 = _guard24047 & _guard24048;
wire _guard24050 = cond_wire599_out;
wire _guard24051 = early_reset_static_par0_go_out;
wire _guard24052 = _guard24050 & _guard24051;
wire _guard24053 = cond_wire599_out;
wire _guard24054 = early_reset_static_par0_go_out;
wire _guard24055 = _guard24053 & _guard24054;
wire _guard24056 = fsm0_out == 6'd0;
wire _guard24057 = early_reset_static_seq_go_out;
wire _guard24058 = _guard24056 & _guard24057;
wire _guard24059 = early_reset_static_par0_go_out;
wire _guard24060 = _guard24058 | _guard24059;
wire _guard24061 = early_reset_static_par0_go_out;
wire _guard24062 = fsm0_out == 6'd0;
wire _guard24063 = early_reset_static_seq_go_out;
wire _guard24064 = _guard24062 & _guard24063;
wire _guard24065 = fsm0_out == 6'd0;
wire _guard24066 = early_reset_static_seq_go_out;
wire _guard24067 = _guard24065 & _guard24066;
wire _guard24068 = early_reset_static_par0_go_out;
wire _guard24069 = _guard24067 | _guard24068;
wire _guard24070 = early_reset_static_par0_go_out;
wire _guard24071 = fsm0_out == 6'd0;
wire _guard24072 = early_reset_static_seq_go_out;
wire _guard24073 = _guard24071 & _guard24072;
wire _guard24074 = early_reset_static_par0_go_out;
wire _guard24075 = early_reset_static_par0_go_out;
wire _guard24076 = early_reset_static_par0_go_out;
wire _guard24077 = early_reset_static_par0_go_out;
wire _guard24078 = early_reset_static_par0_go_out;
wire _guard24079 = early_reset_static_par0_go_out;
wire _guard24080 = early_reset_static_par0_go_out;
wire _guard24081 = early_reset_static_par0_go_out;
wire _guard24082 = early_reset_static_par0_go_out;
wire _guard24083 = early_reset_static_par0_go_out;
wire _guard24084 = early_reset_static_par0_go_out;
wire _guard24085 = early_reset_static_par0_go_out;
wire _guard24086 = fsm0_out == 6'd0;
wire _guard24087 = early_reset_static_seq_go_out;
wire _guard24088 = _guard24086 & _guard24087;
wire _guard24089 = early_reset_static_par0_go_out;
wire _guard24090 = _guard24088 | _guard24089;
wire _guard24091 = early_reset_static_par0_go_out;
wire _guard24092 = fsm0_out == 6'd0;
wire _guard24093 = early_reset_static_seq_go_out;
wire _guard24094 = _guard24092 & _guard24093;
wire _guard24095 = early_reset_static_par0_go_out;
wire _guard24096 = early_reset_static_par0_go_out;
wire _guard24097 = early_reset_static_par0_go_out;
wire _guard24098 = early_reset_static_par0_go_out;
wire _guard24099 = fsm0_out == 6'd0;
wire _guard24100 = early_reset_static_seq_go_out;
wire _guard24101 = _guard24099 & _guard24100;
wire _guard24102 = early_reset_static_par0_go_out;
wire _guard24103 = _guard24101 | _guard24102;
wire _guard24104 = early_reset_static_par0_go_out;
wire _guard24105 = fsm0_out == 6'd0;
wire _guard24106 = early_reset_static_seq_go_out;
wire _guard24107 = _guard24105 & _guard24106;
wire _guard24108 = fsm0_out == 6'd0;
wire _guard24109 = early_reset_static_seq_go_out;
wire _guard24110 = _guard24108 & _guard24109;
wire _guard24111 = early_reset_static_par0_go_out;
wire _guard24112 = _guard24110 | _guard24111;
wire _guard24113 = early_reset_static_par0_go_out;
wire _guard24114 = fsm0_out == 6'd0;
wire _guard24115 = early_reset_static_seq_go_out;
wire _guard24116 = _guard24114 & _guard24115;
wire _guard24117 = fsm0_out == 6'd0;
wire _guard24118 = early_reset_static_seq_go_out;
wire _guard24119 = _guard24117 & _guard24118;
wire _guard24120 = early_reset_static_par0_go_out;
wire _guard24121 = _guard24119 | _guard24120;
wire _guard24122 = fsm0_out == 6'd0;
wire _guard24123 = early_reset_static_seq_go_out;
wire _guard24124 = _guard24122 & _guard24123;
wire _guard24125 = early_reset_static_par0_go_out;
wire _guard24126 = fsm0_out == 6'd0;
wire _guard24127 = early_reset_static_seq_go_out;
wire _guard24128 = _guard24126 & _guard24127;
wire _guard24129 = early_reset_static_par0_go_out;
wire _guard24130 = _guard24128 | _guard24129;
wire _guard24131 = fsm0_out == 6'd0;
wire _guard24132 = early_reset_static_seq_go_out;
wire _guard24133 = _guard24131 & _guard24132;
wire _guard24134 = early_reset_static_par0_go_out;
wire _guard24135 = early_reset_static_par0_go_out;
wire _guard24136 = early_reset_static_par0_go_out;
wire _guard24137 = early_reset_static_par0_go_out;
wire _guard24138 = early_reset_static_par0_go_out;
wire _guard24139 = early_reset_static_par0_go_out;
wire _guard24140 = early_reset_static_par0_go_out;
wire _guard24141 = fsm0_out == 6'd0;
wire _guard24142 = early_reset_static_seq_go_out;
wire _guard24143 = _guard24141 & _guard24142;
wire _guard24144 = early_reset_static_par0_go_out;
wire _guard24145 = _guard24143 | _guard24144;
wire _guard24146 = early_reset_static_par0_go_out;
wire _guard24147 = fsm0_out == 6'd0;
wire _guard24148 = early_reset_static_seq_go_out;
wire _guard24149 = _guard24147 & _guard24148;
wire _guard24150 = fsm0_out == 6'd0;
wire _guard24151 = early_reset_static_seq_go_out;
wire _guard24152 = _guard24150 & _guard24151;
wire _guard24153 = early_reset_static_par0_go_out;
wire _guard24154 = _guard24152 | _guard24153;
wire _guard24155 = early_reset_static_par0_go_out;
wire _guard24156 = fsm0_out == 6'd0;
wire _guard24157 = early_reset_static_seq_go_out;
wire _guard24158 = _guard24156 & _guard24157;
wire _guard24159 = early_reset_static_par0_go_out;
wire _guard24160 = early_reset_static_par0_go_out;
wire _guard24161 = early_reset_static_par0_go_out;
wire _guard24162 = early_reset_static_par0_go_out;
wire _guard24163 = early_reset_static_par0_go_out;
wire _guard24164 = ~_guard0;
wire _guard24165 = early_reset_static_par0_go_out;
wire _guard24166 = _guard24164 & _guard24165;
wire _guard24167 = early_reset_static_par0_go_out;
wire _guard24168 = early_reset_static_par0_go_out;
wire _guard24169 = early_reset_static_par0_go_out;
wire _guard24170 = early_reset_static_par0_go_out;
wire _guard24171 = early_reset_static_par0_go_out;
wire _guard24172 = early_reset_static_par0_go_out;
wire _guard24173 = early_reset_static_par0_go_out;
wire _guard24174 = ~_guard0;
wire _guard24175 = early_reset_static_par0_go_out;
wire _guard24176 = _guard24174 & _guard24175;
wire _guard24177 = ~_guard0;
wire _guard24178 = early_reset_static_par0_go_out;
wire _guard24179 = _guard24177 & _guard24178;
wire _guard24180 = early_reset_static_par0_go_out;
wire _guard24181 = early_reset_static_par0_go_out;
wire _guard24182 = early_reset_static_par0_go_out;
wire _guard24183 = ~_guard0;
wire _guard24184 = early_reset_static_par0_go_out;
wire _guard24185 = _guard24183 & _guard24184;
wire _guard24186 = early_reset_static_par0_go_out;
wire _guard24187 = early_reset_static_par0_go_out;
wire _guard24188 = early_reset_static_par0_go_out;
wire _guard24189 = early_reset_static_par0_go_out;
wire _guard24190 = ~_guard0;
wire _guard24191 = early_reset_static_par0_go_out;
wire _guard24192 = _guard24190 & _guard24191;
wire _guard24193 = early_reset_static_par0_go_out;
wire _guard24194 = ~_guard0;
wire _guard24195 = early_reset_static_par0_go_out;
wire _guard24196 = _guard24194 & _guard24195;
wire _guard24197 = ~_guard0;
wire _guard24198 = early_reset_static_par0_go_out;
wire _guard24199 = _guard24197 & _guard24198;
wire _guard24200 = early_reset_static_par0_go_out;
wire _guard24201 = ~_guard0;
wire _guard24202 = early_reset_static_par0_go_out;
wire _guard24203 = _guard24201 & _guard24202;
wire _guard24204 = early_reset_static_par0_go_out;
wire _guard24205 = ~_guard0;
wire _guard24206 = early_reset_static_par0_go_out;
wire _guard24207 = _guard24205 & _guard24206;
wire _guard24208 = early_reset_static_par0_go_out;
wire _guard24209 = early_reset_static_par0_go_out;
wire _guard24210 = early_reset_static_par0_go_out;
wire _guard24211 = early_reset_static_par0_go_out;
wire _guard24212 = ~_guard0;
wire _guard24213 = early_reset_static_par0_go_out;
wire _guard24214 = _guard24212 & _guard24213;
wire _guard24215 = early_reset_static_par0_go_out;
wire _guard24216 = early_reset_static_par0_go_out;
wire _guard24217 = early_reset_static_par0_go_out;
wire _guard24218 = early_reset_static_par0_go_out;
wire _guard24219 = early_reset_static_par0_go_out;
wire _guard24220 = ~_guard0;
wire _guard24221 = early_reset_static_par0_go_out;
wire _guard24222 = _guard24220 & _guard24221;
wire _guard24223 = early_reset_static_par0_go_out;
wire _guard24224 = early_reset_static_par0_go_out;
wire _guard24225 = early_reset_static_par0_go_out;
wire _guard24226 = ~_guard0;
wire _guard24227 = early_reset_static_par0_go_out;
wire _guard24228 = _guard24226 & _guard24227;
wire _guard24229 = ~_guard0;
wire _guard24230 = early_reset_static_par0_go_out;
wire _guard24231 = _guard24229 & _guard24230;
wire _guard24232 = early_reset_static_par0_go_out;
wire _guard24233 = ~_guard0;
wire _guard24234 = early_reset_static_par0_go_out;
wire _guard24235 = _guard24233 & _guard24234;
wire _guard24236 = early_reset_static_par0_go_out;
wire _guard24237 = early_reset_static_par0_go_out;
wire _guard24238 = early_reset_static_par0_go_out;
wire _guard24239 = early_reset_static_par0_go_out;
wire _guard24240 = early_reset_static_par0_go_out;
wire _guard24241 = early_reset_static_par0_go_out;
wire _guard24242 = ~_guard0;
wire _guard24243 = early_reset_static_par0_go_out;
wire _guard24244 = _guard24242 & _guard24243;
wire _guard24245 = ~_guard0;
wire _guard24246 = early_reset_static_par0_go_out;
wire _guard24247 = _guard24245 & _guard24246;
wire _guard24248 = early_reset_static_par0_go_out;
wire _guard24249 = early_reset_static_par0_go_out;
wire _guard24250 = early_reset_static_par0_go_out;
wire _guard24251 = early_reset_static_par0_go_out;
wire _guard24252 = early_reset_static_par0_go_out;
wire _guard24253 = ~_guard0;
wire _guard24254 = early_reset_static_par0_go_out;
wire _guard24255 = _guard24253 & _guard24254;
wire _guard24256 = early_reset_static_par0_go_out;
wire _guard24257 = early_reset_static_par0_go_out;
wire _guard24258 = early_reset_static_par0_go_out;
wire _guard24259 = ~_guard0;
wire _guard24260 = early_reset_static_par0_go_out;
wire _guard24261 = _guard24259 & _guard24260;
wire _guard24262 = early_reset_static_par0_go_out;
wire _guard24263 = early_reset_static_par0_go_out;
wire _guard24264 = early_reset_static_par0_go_out;
wire _guard24265 = ~_guard0;
wire _guard24266 = early_reset_static_par0_go_out;
wire _guard24267 = _guard24265 & _guard24266;
wire _guard24268 = early_reset_static_par0_go_out;
wire _guard24269 = early_reset_static_par0_go_out;
wire _guard24270 = ~_guard0;
wire _guard24271 = early_reset_static_par0_go_out;
wire _guard24272 = _guard24270 & _guard24271;
wire _guard24273 = early_reset_static_par0_go_out;
wire _guard24274 = early_reset_static_par0_go_out;
wire _guard24275 = early_reset_static_par0_go_out;
wire _guard24276 = ~_guard0;
wire _guard24277 = early_reset_static_par0_go_out;
wire _guard24278 = _guard24276 & _guard24277;
wire _guard24279 = early_reset_static_par0_go_out;
wire _guard24280 = early_reset_static_par0_go_out;
wire _guard24281 = early_reset_static_par0_go_out;
wire _guard24282 = early_reset_static_par0_go_out;
wire _guard24283 = early_reset_static_par0_go_out;
wire _guard24284 = early_reset_static_par0_go_out;
wire _guard24285 = early_reset_static_par0_go_out;
wire _guard24286 = early_reset_static_par0_go_out;
wire _guard24287 = early_reset_static_par0_go_out;
wire _guard24288 = early_reset_static_par0_go_out;
wire _guard24289 = early_reset_static_par0_go_out;
wire _guard24290 = early_reset_static_par0_go_out;
wire _guard24291 = early_reset_static_par0_go_out;
wire _guard24292 = early_reset_static_par0_go_out;
wire _guard24293 = early_reset_static_par0_go_out;
wire _guard24294 = early_reset_static_par0_go_out;
wire _guard24295 = early_reset_static_par0_go_out;
wire _guard24296 = early_reset_static_par0_go_out;
wire _guard24297 = early_reset_static_par0_go_out;
wire _guard24298 = early_reset_static_par0_go_out;
wire _guard24299 = early_reset_static_par0_go_out;
wire _guard24300 = early_reset_static_par0_go_out;
wire _guard24301 = early_reset_static_par0_go_out;
wire _guard24302 = ~_guard0;
wire _guard24303 = early_reset_static_par0_go_out;
wire _guard24304 = _guard24302 & _guard24303;
wire _guard24305 = early_reset_static_par0_go_out;
wire _guard24306 = early_reset_static_par0_go_out;
wire _guard24307 = early_reset_static_par0_go_out;
wire _guard24308 = ~_guard0;
wire _guard24309 = early_reset_static_par0_go_out;
wire _guard24310 = _guard24308 & _guard24309;
wire _guard24311 = early_reset_static_par0_go_out;
wire _guard24312 = ~_guard0;
wire _guard24313 = early_reset_static_par0_go_out;
wire _guard24314 = _guard24312 & _guard24313;
wire _guard24315 = early_reset_static_par0_go_out;
wire _guard24316 = ~_guard0;
wire _guard24317 = early_reset_static_par0_go_out;
wire _guard24318 = _guard24316 & _guard24317;
wire _guard24319 = ~_guard0;
wire _guard24320 = early_reset_static_par0_go_out;
wire _guard24321 = _guard24319 & _guard24320;
wire _guard24322 = early_reset_static_par0_go_out;
wire _guard24323 = early_reset_static_par0_go_out;
wire _guard24324 = ~_guard0;
wire _guard24325 = early_reset_static_par0_go_out;
wire _guard24326 = _guard24324 & _guard24325;
wire _guard24327 = early_reset_static_par0_go_out;
wire _guard24328 = ~_guard0;
wire _guard24329 = early_reset_static_par0_go_out;
wire _guard24330 = _guard24328 & _guard24329;
wire _guard24331 = ~_guard0;
wire _guard24332 = early_reset_static_par0_go_out;
wire _guard24333 = _guard24331 & _guard24332;
wire _guard24334 = early_reset_static_par0_go_out;
wire _guard24335 = early_reset_static_par0_go_out;
wire _guard24336 = ~_guard0;
wire _guard24337 = early_reset_static_par0_go_out;
wire _guard24338 = _guard24336 & _guard24337;
wire _guard24339 = ~_guard0;
wire _guard24340 = early_reset_static_par0_go_out;
wire _guard24341 = _guard24339 & _guard24340;
wire _guard24342 = early_reset_static_par0_go_out;
wire _guard24343 = early_reset_static_par0_go_out;
wire _guard24344 = early_reset_static_par0_go_out;
wire _guard24345 = ~_guard0;
wire _guard24346 = early_reset_static_par0_go_out;
wire _guard24347 = _guard24345 & _guard24346;
wire _guard24348 = early_reset_static_par0_go_out;
wire _guard24349 = early_reset_static_par0_go_out;
wire _guard24350 = early_reset_static_par0_go_out;
wire _guard24351 = early_reset_static_par0_go_out;
wire _guard24352 = ~_guard0;
wire _guard24353 = early_reset_static_par0_go_out;
wire _guard24354 = _guard24352 & _guard24353;
wire _guard24355 = early_reset_static_par0_go_out;
wire _guard24356 = ~_guard0;
wire _guard24357 = early_reset_static_par0_go_out;
wire _guard24358 = _guard24356 & _guard24357;
wire _guard24359 = early_reset_static_par0_go_out;
wire _guard24360 = early_reset_static_par0_go_out;
wire _guard24361 = early_reset_static_par0_go_out;
wire _guard24362 = ~_guard0;
wire _guard24363 = early_reset_static_par0_go_out;
wire _guard24364 = _guard24362 & _guard24363;
wire _guard24365 = ~_guard0;
wire _guard24366 = early_reset_static_par0_go_out;
wire _guard24367 = _guard24365 & _guard24366;
wire _guard24368 = early_reset_static_par0_go_out;
wire _guard24369 = early_reset_static_par0_go_out;
wire _guard24370 = early_reset_static_par0_go_out;
wire _guard24371 = early_reset_static_par0_go_out;
wire _guard24372 = early_reset_static_par0_go_out;
wire _guard24373 = ~_guard0;
wire _guard24374 = early_reset_static_par0_go_out;
wire _guard24375 = _guard24373 & _guard24374;
wire _guard24376 = early_reset_static_par0_go_out;
wire _guard24377 = early_reset_static_par0_go_out;
wire _guard24378 = early_reset_static_par0_go_out;
wire _guard24379 = early_reset_static_par0_go_out;
wire _guard24380 = early_reset_static_par0_go_out;
wire _guard24381 = early_reset_static_par0_go_out;
wire _guard24382 = ~_guard0;
wire _guard24383 = early_reset_static_par0_go_out;
wire _guard24384 = _guard24382 & _guard24383;
wire _guard24385 = early_reset_static_par0_go_out;
wire _guard24386 = ~_guard0;
wire _guard24387 = early_reset_static_par0_go_out;
wire _guard24388 = _guard24386 & _guard24387;
wire _guard24389 = early_reset_static_par0_go_out;
wire _guard24390 = ~_guard0;
wire _guard24391 = early_reset_static_par0_go_out;
wire _guard24392 = _guard24390 & _guard24391;
wire _guard24393 = early_reset_static_par0_go_out;
wire _guard24394 = early_reset_static_par0_go_out;
wire _guard24395 = early_reset_static_par0_go_out;
wire _guard24396 = early_reset_static_par0_go_out;
wire _guard24397 = ~_guard0;
wire _guard24398 = early_reset_static_par0_go_out;
wire _guard24399 = _guard24397 & _guard24398;
wire _guard24400 = early_reset_static_par0_go_out;
wire _guard24401 = early_reset_static_par0_go_out;
wire _guard24402 = ~_guard0;
wire _guard24403 = early_reset_static_par0_go_out;
wire _guard24404 = _guard24402 & _guard24403;
wire _guard24405 = early_reset_static_par0_go_out;
wire _guard24406 = ~_guard0;
wire _guard24407 = early_reset_static_par0_go_out;
wire _guard24408 = _guard24406 & _guard24407;
wire _guard24409 = early_reset_static_par0_go_out;
wire _guard24410 = early_reset_static_par0_go_out;
wire _guard24411 = early_reset_static_par0_go_out;
wire _guard24412 = early_reset_static_par0_go_out;
wire _guard24413 = ~_guard0;
wire _guard24414 = early_reset_static_par0_go_out;
wire _guard24415 = _guard24413 & _guard24414;
wire _guard24416 = early_reset_static_par0_go_out;
wire _guard24417 = ~_guard0;
wire _guard24418 = early_reset_static_par0_go_out;
wire _guard24419 = _guard24417 & _guard24418;
wire _guard24420 = early_reset_static_par0_go_out;
wire _guard24421 = early_reset_static_par0_go_out;
wire _guard24422 = ~_guard0;
wire _guard24423 = early_reset_static_par0_go_out;
wire _guard24424 = _guard24422 & _guard24423;
wire _guard24425 = early_reset_static_par0_go_out;
wire _guard24426 = early_reset_static_par0_go_out;
wire _guard24427 = ~_guard0;
wire _guard24428 = early_reset_static_par0_go_out;
wire _guard24429 = _guard24427 & _guard24428;
wire _guard24430 = early_reset_static_par0_go_out;
wire _guard24431 = early_reset_static_par0_go_out;
wire _guard24432 = early_reset_static_par0_go_out;
wire _guard24433 = early_reset_static_par0_go_out;
wire _guard24434 = early_reset_static_par0_go_out;
wire _guard24435 = early_reset_static_par0_go_out;
wire _guard24436 = ~_guard0;
wire _guard24437 = early_reset_static_par0_go_out;
wire _guard24438 = _guard24436 & _guard24437;
wire _guard24439 = early_reset_static_par0_go_out;
wire _guard24440 = ~_guard0;
wire _guard24441 = early_reset_static_par0_go_out;
wire _guard24442 = _guard24440 & _guard24441;
wire _guard24443 = early_reset_static_par0_go_out;
wire _guard24444 = ~_guard0;
wire _guard24445 = early_reset_static_par0_go_out;
wire _guard24446 = _guard24444 & _guard24445;
wire _guard24447 = early_reset_static_par0_go_out;
wire _guard24448 = early_reset_static_par0_go_out;
wire _guard24449 = early_reset_static_par0_go_out;
wire _guard24450 = ~_guard0;
wire _guard24451 = early_reset_static_par0_go_out;
wire _guard24452 = _guard24450 & _guard24451;
wire _guard24453 = early_reset_static_par0_go_out;
wire _guard24454 = ~_guard0;
wire _guard24455 = early_reset_static_par0_go_out;
wire _guard24456 = _guard24454 & _guard24455;
wire _guard24457 = ~_guard0;
wire _guard24458 = early_reset_static_par0_go_out;
wire _guard24459 = _guard24457 & _guard24458;
wire _guard24460 = early_reset_static_par0_go_out;
wire _guard24461 = ~_guard0;
wire _guard24462 = early_reset_static_par0_go_out;
wire _guard24463 = _guard24461 & _guard24462;
wire _guard24464 = early_reset_static_par0_go_out;
wire _guard24465 = early_reset_static_par0_go_out;
wire _guard24466 = early_reset_static_par0_go_out;
wire _guard24467 = ~_guard0;
wire _guard24468 = early_reset_static_par0_go_out;
wire _guard24469 = _guard24467 & _guard24468;
wire _guard24470 = early_reset_static_par0_go_out;
wire _guard24471 = ~_guard0;
wire _guard24472 = early_reset_static_par0_go_out;
wire _guard24473 = _guard24471 & _guard24472;
wire _guard24474 = early_reset_static_par0_go_out;
wire _guard24475 = ~_guard0;
wire _guard24476 = early_reset_static_par0_go_out;
wire _guard24477 = _guard24475 & _guard24476;
wire _guard24478 = early_reset_static_par0_go_out;
wire _guard24479 = early_reset_static_par0_go_out;
wire _guard24480 = ~_guard0;
wire _guard24481 = early_reset_static_par0_go_out;
wire _guard24482 = _guard24480 & _guard24481;
wire _guard24483 = ~_guard0;
wire _guard24484 = early_reset_static_par0_go_out;
wire _guard24485 = _guard24483 & _guard24484;
wire _guard24486 = early_reset_static_par0_go_out;
wire _guard24487 = ~_guard0;
wire _guard24488 = early_reset_static_par0_go_out;
wire _guard24489 = _guard24487 & _guard24488;
wire _guard24490 = early_reset_static_par0_go_out;
wire _guard24491 = ~_guard0;
wire _guard24492 = early_reset_static_par0_go_out;
wire _guard24493 = _guard24491 & _guard24492;
wire _guard24494 = early_reset_static_par0_go_out;
wire _guard24495 = early_reset_static_par0_go_out;
wire _guard24496 = ~_guard0;
wire _guard24497 = early_reset_static_par0_go_out;
wire _guard24498 = _guard24496 & _guard24497;
wire _guard24499 = early_reset_static_par0_go_out;
wire _guard24500 = early_reset_static_par0_go_out;
wire _guard24501 = early_reset_static_par0_go_out;
wire _guard24502 = early_reset_static_par0_go_out;
wire _guard24503 = early_reset_static_par0_go_out;
wire _guard24504 = early_reset_static_par0_go_out;
wire _guard24505 = ~_guard0;
wire _guard24506 = early_reset_static_par0_go_out;
wire _guard24507 = _guard24505 & _guard24506;
wire _guard24508 = early_reset_static_par0_go_out;
wire _guard24509 = early_reset_static_par0_go_out;
wire _guard24510 = early_reset_static_par0_go_out;
wire _guard24511 = early_reset_static_par0_go_out;
wire _guard24512 = ~_guard0;
wire _guard24513 = early_reset_static_par0_go_out;
wire _guard24514 = _guard24512 & _guard24513;
wire _guard24515 = early_reset_static_par0_go_out;
wire _guard24516 = early_reset_static_par0_go_out;
wire _guard24517 = early_reset_static_par0_go_out;
wire _guard24518 = early_reset_static_par0_go_out;
wire _guard24519 = early_reset_static_par0_go_out;
wire _guard24520 = early_reset_static_par0_go_out;
wire _guard24521 = ~_guard0;
wire _guard24522 = early_reset_static_par0_go_out;
wire _guard24523 = _guard24521 & _guard24522;
wire _guard24524 = early_reset_static_par0_go_out;
wire _guard24525 = early_reset_static_par0_go_out;
wire _guard24526 = early_reset_static_par0_go_out;
wire _guard24527 = early_reset_static_par0_go_out;
wire _guard24528 = ~_guard0;
wire _guard24529 = early_reset_static_par0_go_out;
wire _guard24530 = _guard24528 & _guard24529;
wire _guard24531 = early_reset_static_par0_go_out;
wire _guard24532 = early_reset_static_par0_go_out;
wire _guard24533 = ~_guard0;
wire _guard24534 = early_reset_static_par0_go_out;
wire _guard24535 = _guard24533 & _guard24534;
wire _guard24536 = early_reset_static_par0_go_out;
wire _guard24537 = early_reset_static_par0_go_out;
wire _guard24538 = early_reset_static_par0_go_out;
wire _guard24539 = early_reset_static_par0_go_out;
wire _guard24540 = early_reset_static_par0_go_out;
wire _guard24541 = ~_guard0;
wire _guard24542 = early_reset_static_par0_go_out;
wire _guard24543 = _guard24541 & _guard24542;
wire _guard24544 = early_reset_static_par0_go_out;
wire _guard24545 = early_reset_static_par0_go_out;
wire _guard24546 = ~_guard0;
wire _guard24547 = early_reset_static_par0_go_out;
wire _guard24548 = _guard24546 & _guard24547;
wire _guard24549 = early_reset_static_par0_go_out;
wire _guard24550 = ~_guard0;
wire _guard24551 = early_reset_static_par0_go_out;
wire _guard24552 = _guard24550 & _guard24551;
wire _guard24553 = early_reset_static_par0_go_out;
wire _guard24554 = early_reset_static_par0_go_out;
wire _guard24555 = early_reset_static_par0_go_out;
wire _guard24556 = ~_guard0;
wire _guard24557 = early_reset_static_par0_go_out;
wire _guard24558 = _guard24556 & _guard24557;
wire _guard24559 = early_reset_static_par0_go_out;
wire _guard24560 = ~_guard0;
wire _guard24561 = early_reset_static_par0_go_out;
wire _guard24562 = _guard24560 & _guard24561;
wire _guard24563 = early_reset_static_par0_go_out;
wire _guard24564 = early_reset_static_par0_go_out;
wire _guard24565 = early_reset_static_par0_go_out;
wire _guard24566 = early_reset_static_par0_go_out;
wire _guard24567 = early_reset_static_par0_go_out;
wire _guard24568 = early_reset_static_par0_go_out;
wire _guard24569 = ~_guard0;
wire _guard24570 = early_reset_static_par0_go_out;
wire _guard24571 = _guard24569 & _guard24570;
wire _guard24572 = early_reset_static_par0_go_out;
wire _guard24573 = early_reset_static_par0_go_out;
wire _guard24574 = early_reset_static_par0_go_out;
wire _guard24575 = early_reset_static_par0_go_out;
wire _guard24576 = ~_guard0;
wire _guard24577 = early_reset_static_par0_go_out;
wire _guard24578 = _guard24576 & _guard24577;
wire _guard24579 = ~_guard0;
wire _guard24580 = early_reset_static_par0_go_out;
wire _guard24581 = _guard24579 & _guard24580;
wire _guard24582 = early_reset_static_par0_go_out;
wire _guard24583 = early_reset_static_par0_go_out;
wire _guard24584 = early_reset_static_par0_go_out;
wire _guard24585 = early_reset_static_par0_go_out;
wire _guard24586 = early_reset_static_par0_go_out;
wire _guard24587 = early_reset_static_par0_go_out;
wire _guard24588 = early_reset_static_par0_go_out;
wire _guard24589 = early_reset_static_par0_go_out;
wire _guard24590 = early_reset_static_par0_go_out;
wire _guard24591 = early_reset_static_par0_go_out;
wire _guard24592 = early_reset_static_par0_go_out;
wire _guard24593 = early_reset_static_par0_go_out;
wire _guard24594 = early_reset_static_par0_go_out;
wire _guard24595 = cond_wire1_out;
wire _guard24596 = early_reset_static_par0_go_out;
wire _guard24597 = _guard24595 & _guard24596;
wire _guard24598 = cond_wire1_out;
wire _guard24599 = early_reset_static_par0_go_out;
wire _guard24600 = _guard24598 & _guard24599;
wire _guard24601 = cond_wire34_out;
wire _guard24602 = early_reset_static_par0_go_out;
wire _guard24603 = _guard24601 & _guard24602;
wire _guard24604 = cond_wire34_out;
wire _guard24605 = early_reset_static_par0_go_out;
wire _guard24606 = _guard24604 & _guard24605;
wire _guard24607 = cond_wire51_out;
wire _guard24608 = early_reset_static_par0_go_out;
wire _guard24609 = _guard24607 & _guard24608;
wire _guard24610 = cond_wire51_out;
wire _guard24611 = early_reset_static_par0_go_out;
wire _guard24612 = _guard24610 & _guard24611;
wire _guard24613 = cond_wire67_out;
wire _guard24614 = early_reset_static_par0_go_out;
wire _guard24615 = _guard24613 & _guard24614;
wire _guard24616 = cond_wire65_out;
wire _guard24617 = early_reset_static_par0_go_out;
wire _guard24618 = _guard24616 & _guard24617;
wire _guard24619 = fsm_out == 1'd0;
wire _guard24620 = cond_wire65_out;
wire _guard24621 = _guard24619 & _guard24620;
wire _guard24622 = fsm_out == 1'd0;
wire _guard24623 = _guard24621 & _guard24622;
wire _guard24624 = fsm_out == 1'd0;
wire _guard24625 = cond_wire67_out;
wire _guard24626 = _guard24624 & _guard24625;
wire _guard24627 = fsm_out == 1'd0;
wire _guard24628 = _guard24626 & _guard24627;
wire _guard24629 = _guard24623 | _guard24628;
wire _guard24630 = early_reset_static_par0_go_out;
wire _guard24631 = _guard24629 & _guard24630;
wire _guard24632 = fsm_out == 1'd0;
wire _guard24633 = cond_wire65_out;
wire _guard24634 = _guard24632 & _guard24633;
wire _guard24635 = fsm_out == 1'd0;
wire _guard24636 = _guard24634 & _guard24635;
wire _guard24637 = fsm_out == 1'd0;
wire _guard24638 = cond_wire67_out;
wire _guard24639 = _guard24637 & _guard24638;
wire _guard24640 = fsm_out == 1'd0;
wire _guard24641 = _guard24639 & _guard24640;
wire _guard24642 = _guard24636 | _guard24641;
wire _guard24643 = early_reset_static_par0_go_out;
wire _guard24644 = _guard24642 & _guard24643;
wire _guard24645 = fsm_out == 1'd0;
wire _guard24646 = cond_wire65_out;
wire _guard24647 = _guard24645 & _guard24646;
wire _guard24648 = fsm_out == 1'd0;
wire _guard24649 = _guard24647 & _guard24648;
wire _guard24650 = fsm_out == 1'd0;
wire _guard24651 = cond_wire67_out;
wire _guard24652 = _guard24650 & _guard24651;
wire _guard24653 = fsm_out == 1'd0;
wire _guard24654 = _guard24652 & _guard24653;
wire _guard24655 = _guard24649 | _guard24654;
wire _guard24656 = early_reset_static_par0_go_out;
wire _guard24657 = _guard24655 & _guard24656;
wire _guard24658 = cond_wire64_out;
wire _guard24659 = early_reset_static_par0_go_out;
wire _guard24660 = _guard24658 & _guard24659;
wire _guard24661 = cond_wire64_out;
wire _guard24662 = early_reset_static_par0_go_out;
wire _guard24663 = _guard24661 & _guard24662;
wire _guard24664 = cond_wire71_out;
wire _guard24665 = early_reset_static_par0_go_out;
wire _guard24666 = _guard24664 & _guard24665;
wire _guard24667 = cond_wire71_out;
wire _guard24668 = early_reset_static_par0_go_out;
wire _guard24669 = _guard24667 & _guard24668;
wire _guard24670 = cond_wire105_out;
wire _guard24671 = early_reset_static_par0_go_out;
wire _guard24672 = _guard24670 & _guard24671;
wire _guard24673 = cond_wire105_out;
wire _guard24674 = early_reset_static_par0_go_out;
wire _guard24675 = _guard24673 & _guard24674;
wire _guard24676 = cond_wire122_out;
wire _guard24677 = early_reset_static_par0_go_out;
wire _guard24678 = _guard24676 & _guard24677;
wire _guard24679 = cond_wire120_out;
wire _guard24680 = early_reset_static_par0_go_out;
wire _guard24681 = _guard24679 & _guard24680;
wire _guard24682 = fsm_out == 1'd0;
wire _guard24683 = cond_wire120_out;
wire _guard24684 = _guard24682 & _guard24683;
wire _guard24685 = fsm_out == 1'd0;
wire _guard24686 = _guard24684 & _guard24685;
wire _guard24687 = fsm_out == 1'd0;
wire _guard24688 = cond_wire122_out;
wire _guard24689 = _guard24687 & _guard24688;
wire _guard24690 = fsm_out == 1'd0;
wire _guard24691 = _guard24689 & _guard24690;
wire _guard24692 = _guard24686 | _guard24691;
wire _guard24693 = early_reset_static_par0_go_out;
wire _guard24694 = _guard24692 & _guard24693;
wire _guard24695 = fsm_out == 1'd0;
wire _guard24696 = cond_wire120_out;
wire _guard24697 = _guard24695 & _guard24696;
wire _guard24698 = fsm_out == 1'd0;
wire _guard24699 = _guard24697 & _guard24698;
wire _guard24700 = fsm_out == 1'd0;
wire _guard24701 = cond_wire122_out;
wire _guard24702 = _guard24700 & _guard24701;
wire _guard24703 = fsm_out == 1'd0;
wire _guard24704 = _guard24702 & _guard24703;
wire _guard24705 = _guard24699 | _guard24704;
wire _guard24706 = early_reset_static_par0_go_out;
wire _guard24707 = _guard24705 & _guard24706;
wire _guard24708 = fsm_out == 1'd0;
wire _guard24709 = cond_wire120_out;
wire _guard24710 = _guard24708 & _guard24709;
wire _guard24711 = fsm_out == 1'd0;
wire _guard24712 = _guard24710 & _guard24711;
wire _guard24713 = fsm_out == 1'd0;
wire _guard24714 = cond_wire122_out;
wire _guard24715 = _guard24713 & _guard24714;
wire _guard24716 = fsm_out == 1'd0;
wire _guard24717 = _guard24715 & _guard24716;
wire _guard24718 = _guard24712 | _guard24717;
wire _guard24719 = early_reset_static_par0_go_out;
wire _guard24720 = _guard24718 & _guard24719;
wire _guard24721 = cond_wire138_out;
wire _guard24722 = early_reset_static_par0_go_out;
wire _guard24723 = _guard24721 & _guard24722;
wire _guard24724 = cond_wire136_out;
wire _guard24725 = early_reset_static_par0_go_out;
wire _guard24726 = _guard24724 & _guard24725;
wire _guard24727 = fsm_out == 1'd0;
wire _guard24728 = cond_wire136_out;
wire _guard24729 = _guard24727 & _guard24728;
wire _guard24730 = fsm_out == 1'd0;
wire _guard24731 = _guard24729 & _guard24730;
wire _guard24732 = fsm_out == 1'd0;
wire _guard24733 = cond_wire138_out;
wire _guard24734 = _guard24732 & _guard24733;
wire _guard24735 = fsm_out == 1'd0;
wire _guard24736 = _guard24734 & _guard24735;
wire _guard24737 = _guard24731 | _guard24736;
wire _guard24738 = early_reset_static_par0_go_out;
wire _guard24739 = _guard24737 & _guard24738;
wire _guard24740 = fsm_out == 1'd0;
wire _guard24741 = cond_wire136_out;
wire _guard24742 = _guard24740 & _guard24741;
wire _guard24743 = fsm_out == 1'd0;
wire _guard24744 = _guard24742 & _guard24743;
wire _guard24745 = fsm_out == 1'd0;
wire _guard24746 = cond_wire138_out;
wire _guard24747 = _guard24745 & _guard24746;
wire _guard24748 = fsm_out == 1'd0;
wire _guard24749 = _guard24747 & _guard24748;
wire _guard24750 = _guard24744 | _guard24749;
wire _guard24751 = early_reset_static_par0_go_out;
wire _guard24752 = _guard24750 & _guard24751;
wire _guard24753 = fsm_out == 1'd0;
wire _guard24754 = cond_wire136_out;
wire _guard24755 = _guard24753 & _guard24754;
wire _guard24756 = fsm_out == 1'd0;
wire _guard24757 = _guard24755 & _guard24756;
wire _guard24758 = fsm_out == 1'd0;
wire _guard24759 = cond_wire138_out;
wire _guard24760 = _guard24758 & _guard24759;
wire _guard24761 = fsm_out == 1'd0;
wire _guard24762 = _guard24760 & _guard24761;
wire _guard24763 = _guard24757 | _guard24762;
wire _guard24764 = early_reset_static_par0_go_out;
wire _guard24765 = _guard24763 & _guard24764;
wire _guard24766 = cond_wire155_out;
wire _guard24767 = early_reset_static_par0_go_out;
wire _guard24768 = _guard24766 & _guard24767;
wire _guard24769 = cond_wire153_out;
wire _guard24770 = early_reset_static_par0_go_out;
wire _guard24771 = _guard24769 & _guard24770;
wire _guard24772 = fsm_out == 1'd0;
wire _guard24773 = cond_wire153_out;
wire _guard24774 = _guard24772 & _guard24773;
wire _guard24775 = fsm_out == 1'd0;
wire _guard24776 = _guard24774 & _guard24775;
wire _guard24777 = fsm_out == 1'd0;
wire _guard24778 = cond_wire155_out;
wire _guard24779 = _guard24777 & _guard24778;
wire _guard24780 = fsm_out == 1'd0;
wire _guard24781 = _guard24779 & _guard24780;
wire _guard24782 = _guard24776 | _guard24781;
wire _guard24783 = early_reset_static_par0_go_out;
wire _guard24784 = _guard24782 & _guard24783;
wire _guard24785 = fsm_out == 1'd0;
wire _guard24786 = cond_wire153_out;
wire _guard24787 = _guard24785 & _guard24786;
wire _guard24788 = fsm_out == 1'd0;
wire _guard24789 = _guard24787 & _guard24788;
wire _guard24790 = fsm_out == 1'd0;
wire _guard24791 = cond_wire155_out;
wire _guard24792 = _guard24790 & _guard24791;
wire _guard24793 = fsm_out == 1'd0;
wire _guard24794 = _guard24792 & _guard24793;
wire _guard24795 = _guard24789 | _guard24794;
wire _guard24796 = early_reset_static_par0_go_out;
wire _guard24797 = _guard24795 & _guard24796;
wire _guard24798 = fsm_out == 1'd0;
wire _guard24799 = cond_wire153_out;
wire _guard24800 = _guard24798 & _guard24799;
wire _guard24801 = fsm_out == 1'd0;
wire _guard24802 = _guard24800 & _guard24801;
wire _guard24803 = fsm_out == 1'd0;
wire _guard24804 = cond_wire155_out;
wire _guard24805 = _guard24803 & _guard24804;
wire _guard24806 = fsm_out == 1'd0;
wire _guard24807 = _guard24805 & _guard24806;
wire _guard24808 = _guard24802 | _guard24807;
wire _guard24809 = early_reset_static_par0_go_out;
wire _guard24810 = _guard24808 & _guard24809;
wire _guard24811 = cond_wire183_out;
wire _guard24812 = early_reset_static_par0_go_out;
wire _guard24813 = _guard24811 & _guard24812;
wire _guard24814 = cond_wire181_out;
wire _guard24815 = early_reset_static_par0_go_out;
wire _guard24816 = _guard24814 & _guard24815;
wire _guard24817 = fsm_out == 1'd0;
wire _guard24818 = cond_wire181_out;
wire _guard24819 = _guard24817 & _guard24818;
wire _guard24820 = fsm_out == 1'd0;
wire _guard24821 = _guard24819 & _guard24820;
wire _guard24822 = fsm_out == 1'd0;
wire _guard24823 = cond_wire183_out;
wire _guard24824 = _guard24822 & _guard24823;
wire _guard24825 = fsm_out == 1'd0;
wire _guard24826 = _guard24824 & _guard24825;
wire _guard24827 = _guard24821 | _guard24826;
wire _guard24828 = early_reset_static_par0_go_out;
wire _guard24829 = _guard24827 & _guard24828;
wire _guard24830 = fsm_out == 1'd0;
wire _guard24831 = cond_wire181_out;
wire _guard24832 = _guard24830 & _guard24831;
wire _guard24833 = fsm_out == 1'd0;
wire _guard24834 = _guard24832 & _guard24833;
wire _guard24835 = fsm_out == 1'd0;
wire _guard24836 = cond_wire183_out;
wire _guard24837 = _guard24835 & _guard24836;
wire _guard24838 = fsm_out == 1'd0;
wire _guard24839 = _guard24837 & _guard24838;
wire _guard24840 = _guard24834 | _guard24839;
wire _guard24841 = early_reset_static_par0_go_out;
wire _guard24842 = _guard24840 & _guard24841;
wire _guard24843 = fsm_out == 1'd0;
wire _guard24844 = cond_wire181_out;
wire _guard24845 = _guard24843 & _guard24844;
wire _guard24846 = fsm_out == 1'd0;
wire _guard24847 = _guard24845 & _guard24846;
wire _guard24848 = fsm_out == 1'd0;
wire _guard24849 = cond_wire183_out;
wire _guard24850 = _guard24848 & _guard24849;
wire _guard24851 = fsm_out == 1'd0;
wire _guard24852 = _guard24850 & _guard24851;
wire _guard24853 = _guard24847 | _guard24852;
wire _guard24854 = early_reset_static_par0_go_out;
wire _guard24855 = _guard24853 & _guard24854;
wire _guard24856 = cond_wire117_out;
wire _guard24857 = early_reset_static_par0_go_out;
wire _guard24858 = _guard24856 & _guard24857;
wire _guard24859 = cond_wire117_out;
wire _guard24860 = early_reset_static_par0_go_out;
wire _guard24861 = _guard24859 & _guard24860;
wire _guard24862 = cond_wire187_out;
wire _guard24863 = early_reset_static_par0_go_out;
wire _guard24864 = _guard24862 & _guard24863;
wire _guard24865 = cond_wire185_out;
wire _guard24866 = early_reset_static_par0_go_out;
wire _guard24867 = _guard24865 & _guard24866;
wire _guard24868 = fsm_out == 1'd0;
wire _guard24869 = cond_wire185_out;
wire _guard24870 = _guard24868 & _guard24869;
wire _guard24871 = fsm_out == 1'd0;
wire _guard24872 = _guard24870 & _guard24871;
wire _guard24873 = fsm_out == 1'd0;
wire _guard24874 = cond_wire187_out;
wire _guard24875 = _guard24873 & _guard24874;
wire _guard24876 = fsm_out == 1'd0;
wire _guard24877 = _guard24875 & _guard24876;
wire _guard24878 = _guard24872 | _guard24877;
wire _guard24879 = early_reset_static_par0_go_out;
wire _guard24880 = _guard24878 & _guard24879;
wire _guard24881 = fsm_out == 1'd0;
wire _guard24882 = cond_wire185_out;
wire _guard24883 = _guard24881 & _guard24882;
wire _guard24884 = fsm_out == 1'd0;
wire _guard24885 = _guard24883 & _guard24884;
wire _guard24886 = fsm_out == 1'd0;
wire _guard24887 = cond_wire187_out;
wire _guard24888 = _guard24886 & _guard24887;
wire _guard24889 = fsm_out == 1'd0;
wire _guard24890 = _guard24888 & _guard24889;
wire _guard24891 = _guard24885 | _guard24890;
wire _guard24892 = early_reset_static_par0_go_out;
wire _guard24893 = _guard24891 & _guard24892;
wire _guard24894 = fsm_out == 1'd0;
wire _guard24895 = cond_wire185_out;
wire _guard24896 = _guard24894 & _guard24895;
wire _guard24897 = fsm_out == 1'd0;
wire _guard24898 = _guard24896 & _guard24897;
wire _guard24899 = fsm_out == 1'd0;
wire _guard24900 = cond_wire187_out;
wire _guard24901 = _guard24899 & _guard24900;
wire _guard24902 = fsm_out == 1'd0;
wire _guard24903 = _guard24901 & _guard24902;
wire _guard24904 = _guard24898 | _guard24903;
wire _guard24905 = early_reset_static_par0_go_out;
wire _guard24906 = _guard24904 & _guard24905;
wire _guard24907 = cond_wire194_out;
wire _guard24908 = early_reset_static_par0_go_out;
wire _guard24909 = _guard24907 & _guard24908;
wire _guard24910 = cond_wire194_out;
wire _guard24911 = early_reset_static_par0_go_out;
wire _guard24912 = _guard24910 & _guard24911;
wire _guard24913 = cond_wire281_out;
wire _guard24914 = early_reset_static_par0_go_out;
wire _guard24915 = _guard24913 & _guard24914;
wire _guard24916 = cond_wire279_out;
wire _guard24917 = early_reset_static_par0_go_out;
wire _guard24918 = _guard24916 & _guard24917;
wire _guard24919 = fsm_out == 1'd0;
wire _guard24920 = cond_wire279_out;
wire _guard24921 = _guard24919 & _guard24920;
wire _guard24922 = fsm_out == 1'd0;
wire _guard24923 = _guard24921 & _guard24922;
wire _guard24924 = fsm_out == 1'd0;
wire _guard24925 = cond_wire281_out;
wire _guard24926 = _guard24924 & _guard24925;
wire _guard24927 = fsm_out == 1'd0;
wire _guard24928 = _guard24926 & _guard24927;
wire _guard24929 = _guard24923 | _guard24928;
wire _guard24930 = early_reset_static_par0_go_out;
wire _guard24931 = _guard24929 & _guard24930;
wire _guard24932 = fsm_out == 1'd0;
wire _guard24933 = cond_wire279_out;
wire _guard24934 = _guard24932 & _guard24933;
wire _guard24935 = fsm_out == 1'd0;
wire _guard24936 = _guard24934 & _guard24935;
wire _guard24937 = fsm_out == 1'd0;
wire _guard24938 = cond_wire281_out;
wire _guard24939 = _guard24937 & _guard24938;
wire _guard24940 = fsm_out == 1'd0;
wire _guard24941 = _guard24939 & _guard24940;
wire _guard24942 = _guard24936 | _guard24941;
wire _guard24943 = early_reset_static_par0_go_out;
wire _guard24944 = _guard24942 & _guard24943;
wire _guard24945 = fsm_out == 1'd0;
wire _guard24946 = cond_wire279_out;
wire _guard24947 = _guard24945 & _guard24946;
wire _guard24948 = fsm_out == 1'd0;
wire _guard24949 = _guard24947 & _guard24948;
wire _guard24950 = fsm_out == 1'd0;
wire _guard24951 = cond_wire281_out;
wire _guard24952 = _guard24950 & _guard24951;
wire _guard24953 = fsm_out == 1'd0;
wire _guard24954 = _guard24952 & _guard24953;
wire _guard24955 = _guard24949 | _guard24954;
wire _guard24956 = early_reset_static_par0_go_out;
wire _guard24957 = _guard24955 & _guard24956;
wire _guard24958 = cond_wire284_out;
wire _guard24959 = early_reset_static_par0_go_out;
wire _guard24960 = _guard24958 & _guard24959;
wire _guard24961 = cond_wire284_out;
wire _guard24962 = early_reset_static_par0_go_out;
wire _guard24963 = _guard24961 & _guard24962;
wire _guard24964 = cond_wire251_out;
wire _guard24965 = early_reset_static_par0_go_out;
wire _guard24966 = _guard24964 & _guard24965;
wire _guard24967 = cond_wire251_out;
wire _guard24968 = early_reset_static_par0_go_out;
wire _guard24969 = _guard24967 & _guard24968;
wire _guard24970 = cond_wire320_out;
wire _guard24971 = early_reset_static_par0_go_out;
wire _guard24972 = _guard24970 & _guard24971;
wire _guard24973 = cond_wire320_out;
wire _guard24974 = early_reset_static_par0_go_out;
wire _guard24975 = _guard24973 & _guard24974;
wire _guard24976 = cond_wire324_out;
wire _guard24977 = early_reset_static_par0_go_out;
wire _guard24978 = _guard24976 & _guard24977;
wire _guard24979 = cond_wire324_out;
wire _guard24980 = early_reset_static_par0_go_out;
wire _guard24981 = _guard24979 & _guard24980;
wire _guard24982 = cond_wire271_out;
wire _guard24983 = early_reset_static_par0_go_out;
wire _guard24984 = _guard24982 & _guard24983;
wire _guard24985 = cond_wire271_out;
wire _guard24986 = early_reset_static_par0_go_out;
wire _guard24987 = _guard24985 & _guard24986;
wire _guard24988 = cond_wire390_out;
wire _guard24989 = early_reset_static_par0_go_out;
wire _guard24990 = _guard24988 & _guard24989;
wire _guard24991 = cond_wire388_out;
wire _guard24992 = early_reset_static_par0_go_out;
wire _guard24993 = _guard24991 & _guard24992;
wire _guard24994 = fsm_out == 1'd0;
wire _guard24995 = cond_wire388_out;
wire _guard24996 = _guard24994 & _guard24995;
wire _guard24997 = fsm_out == 1'd0;
wire _guard24998 = _guard24996 & _guard24997;
wire _guard24999 = fsm_out == 1'd0;
wire _guard25000 = cond_wire390_out;
wire _guard25001 = _guard24999 & _guard25000;
wire _guard25002 = fsm_out == 1'd0;
wire _guard25003 = _guard25001 & _guard25002;
wire _guard25004 = _guard24998 | _guard25003;
wire _guard25005 = early_reset_static_par0_go_out;
wire _guard25006 = _guard25004 & _guard25005;
wire _guard25007 = fsm_out == 1'd0;
wire _guard25008 = cond_wire388_out;
wire _guard25009 = _guard25007 & _guard25008;
wire _guard25010 = fsm_out == 1'd0;
wire _guard25011 = _guard25009 & _guard25010;
wire _guard25012 = fsm_out == 1'd0;
wire _guard25013 = cond_wire390_out;
wire _guard25014 = _guard25012 & _guard25013;
wire _guard25015 = fsm_out == 1'd0;
wire _guard25016 = _guard25014 & _guard25015;
wire _guard25017 = _guard25011 | _guard25016;
wire _guard25018 = early_reset_static_par0_go_out;
wire _guard25019 = _guard25017 & _guard25018;
wire _guard25020 = fsm_out == 1'd0;
wire _guard25021 = cond_wire388_out;
wire _guard25022 = _guard25020 & _guard25021;
wire _guard25023 = fsm_out == 1'd0;
wire _guard25024 = _guard25022 & _guard25023;
wire _guard25025 = fsm_out == 1'd0;
wire _guard25026 = cond_wire390_out;
wire _guard25027 = _guard25025 & _guard25026;
wire _guard25028 = fsm_out == 1'd0;
wire _guard25029 = _guard25027 & _guard25028;
wire _guard25030 = _guard25024 | _guard25029;
wire _guard25031 = early_reset_static_par0_go_out;
wire _guard25032 = _guard25030 & _guard25031;
wire _guard25033 = cond_wire414_out;
wire _guard25034 = early_reset_static_par0_go_out;
wire _guard25035 = _guard25033 & _guard25034;
wire _guard25036 = cond_wire414_out;
wire _guard25037 = early_reset_static_par0_go_out;
wire _guard25038 = _guard25036 & _guard25037;
wire _guard25039 = cond_wire443_out;
wire _guard25040 = early_reset_static_par0_go_out;
wire _guard25041 = _guard25039 & _guard25040;
wire _guard25042 = cond_wire441_out;
wire _guard25043 = early_reset_static_par0_go_out;
wire _guard25044 = _guard25042 & _guard25043;
wire _guard25045 = fsm_out == 1'd0;
wire _guard25046 = cond_wire441_out;
wire _guard25047 = _guard25045 & _guard25046;
wire _guard25048 = fsm_out == 1'd0;
wire _guard25049 = _guard25047 & _guard25048;
wire _guard25050 = fsm_out == 1'd0;
wire _guard25051 = cond_wire443_out;
wire _guard25052 = _guard25050 & _guard25051;
wire _guard25053 = fsm_out == 1'd0;
wire _guard25054 = _guard25052 & _guard25053;
wire _guard25055 = _guard25049 | _guard25054;
wire _guard25056 = early_reset_static_par0_go_out;
wire _guard25057 = _guard25055 & _guard25056;
wire _guard25058 = fsm_out == 1'd0;
wire _guard25059 = cond_wire441_out;
wire _guard25060 = _guard25058 & _guard25059;
wire _guard25061 = fsm_out == 1'd0;
wire _guard25062 = _guard25060 & _guard25061;
wire _guard25063 = fsm_out == 1'd0;
wire _guard25064 = cond_wire443_out;
wire _guard25065 = _guard25063 & _guard25064;
wire _guard25066 = fsm_out == 1'd0;
wire _guard25067 = _guard25065 & _guard25066;
wire _guard25068 = _guard25062 | _guard25067;
wire _guard25069 = early_reset_static_par0_go_out;
wire _guard25070 = _guard25068 & _guard25069;
wire _guard25071 = fsm_out == 1'd0;
wire _guard25072 = cond_wire441_out;
wire _guard25073 = _guard25071 & _guard25072;
wire _guard25074 = fsm_out == 1'd0;
wire _guard25075 = _guard25073 & _guard25074;
wire _guard25076 = fsm_out == 1'd0;
wire _guard25077 = cond_wire443_out;
wire _guard25078 = _guard25076 & _guard25077;
wire _guard25079 = fsm_out == 1'd0;
wire _guard25080 = _guard25078 & _guard25079;
wire _guard25081 = _guard25075 | _guard25080;
wire _guard25082 = early_reset_static_par0_go_out;
wire _guard25083 = _guard25081 & _guard25082;
wire _guard25084 = cond_wire381_out;
wire _guard25085 = early_reset_static_par0_go_out;
wire _guard25086 = _guard25084 & _guard25085;
wire _guard25087 = cond_wire381_out;
wire _guard25088 = early_reset_static_par0_go_out;
wire _guard25089 = _guard25087 & _guard25088;
wire _guard25090 = cond_wire511_out;
wire _guard25091 = early_reset_static_par0_go_out;
wire _guard25092 = _guard25090 & _guard25091;
wire _guard25093 = cond_wire511_out;
wire _guard25094 = early_reset_static_par0_go_out;
wire _guard25095 = _guard25093 & _guard25094;
wire _guard25096 = cond_wire454_out;
wire _guard25097 = early_reset_static_par0_go_out;
wire _guard25098 = _guard25096 & _guard25097;
wire _guard25099 = cond_wire454_out;
wire _guard25100 = early_reset_static_par0_go_out;
wire _guard25101 = _guard25099 & _guard25100;
wire _guard25102 = cond_wire475_out;
wire _guard25103 = early_reset_static_par0_go_out;
wire _guard25104 = _guard25102 & _guard25103;
wire _guard25105 = cond_wire475_out;
wire _guard25106 = early_reset_static_par0_go_out;
wire _guard25107 = _guard25105 & _guard25106;
wire _guard25108 = cond_wire565_out;
wire _guard25109 = early_reset_static_par0_go_out;
wire _guard25110 = _guard25108 & _guard25109;
wire _guard25111 = cond_wire563_out;
wire _guard25112 = early_reset_static_par0_go_out;
wire _guard25113 = _guard25111 & _guard25112;
wire _guard25114 = fsm_out == 1'd0;
wire _guard25115 = cond_wire563_out;
wire _guard25116 = _guard25114 & _guard25115;
wire _guard25117 = fsm_out == 1'd0;
wire _guard25118 = _guard25116 & _guard25117;
wire _guard25119 = fsm_out == 1'd0;
wire _guard25120 = cond_wire565_out;
wire _guard25121 = _guard25119 & _guard25120;
wire _guard25122 = fsm_out == 1'd0;
wire _guard25123 = _guard25121 & _guard25122;
wire _guard25124 = _guard25118 | _guard25123;
wire _guard25125 = early_reset_static_par0_go_out;
wire _guard25126 = _guard25124 & _guard25125;
wire _guard25127 = fsm_out == 1'd0;
wire _guard25128 = cond_wire563_out;
wire _guard25129 = _guard25127 & _guard25128;
wire _guard25130 = fsm_out == 1'd0;
wire _guard25131 = _guard25129 & _guard25130;
wire _guard25132 = fsm_out == 1'd0;
wire _guard25133 = cond_wire565_out;
wire _guard25134 = _guard25132 & _guard25133;
wire _guard25135 = fsm_out == 1'd0;
wire _guard25136 = _guard25134 & _guard25135;
wire _guard25137 = _guard25131 | _guard25136;
wire _guard25138 = early_reset_static_par0_go_out;
wire _guard25139 = _guard25137 & _guard25138;
wire _guard25140 = fsm_out == 1'd0;
wire _guard25141 = cond_wire563_out;
wire _guard25142 = _guard25140 & _guard25141;
wire _guard25143 = fsm_out == 1'd0;
wire _guard25144 = _guard25142 & _guard25143;
wire _guard25145 = fsm_out == 1'd0;
wire _guard25146 = cond_wire565_out;
wire _guard25147 = _guard25145 & _guard25146;
wire _guard25148 = fsm_out == 1'd0;
wire _guard25149 = _guard25147 & _guard25148;
wire _guard25150 = _guard25144 | _guard25149;
wire _guard25151 = early_reset_static_par0_go_out;
wire _guard25152 = _guard25150 & _guard25151;
wire _guard25153 = cond_wire569_out;
wire _guard25154 = early_reset_static_par0_go_out;
wire _guard25155 = _guard25153 & _guard25154;
wire _guard25156 = cond_wire567_out;
wire _guard25157 = early_reset_static_par0_go_out;
wire _guard25158 = _guard25156 & _guard25157;
wire _guard25159 = fsm_out == 1'd0;
wire _guard25160 = cond_wire567_out;
wire _guard25161 = _guard25159 & _guard25160;
wire _guard25162 = fsm_out == 1'd0;
wire _guard25163 = _guard25161 & _guard25162;
wire _guard25164 = fsm_out == 1'd0;
wire _guard25165 = cond_wire569_out;
wire _guard25166 = _guard25164 & _guard25165;
wire _guard25167 = fsm_out == 1'd0;
wire _guard25168 = _guard25166 & _guard25167;
wire _guard25169 = _guard25163 | _guard25168;
wire _guard25170 = early_reset_static_par0_go_out;
wire _guard25171 = _guard25169 & _guard25170;
wire _guard25172 = fsm_out == 1'd0;
wire _guard25173 = cond_wire567_out;
wire _guard25174 = _guard25172 & _guard25173;
wire _guard25175 = fsm_out == 1'd0;
wire _guard25176 = _guard25174 & _guard25175;
wire _guard25177 = fsm_out == 1'd0;
wire _guard25178 = cond_wire569_out;
wire _guard25179 = _guard25177 & _guard25178;
wire _guard25180 = fsm_out == 1'd0;
wire _guard25181 = _guard25179 & _guard25180;
wire _guard25182 = _guard25176 | _guard25181;
wire _guard25183 = early_reset_static_par0_go_out;
wire _guard25184 = _guard25182 & _guard25183;
wire _guard25185 = fsm_out == 1'd0;
wire _guard25186 = cond_wire567_out;
wire _guard25187 = _guard25185 & _guard25186;
wire _guard25188 = fsm_out == 1'd0;
wire _guard25189 = _guard25187 & _guard25188;
wire _guard25190 = fsm_out == 1'd0;
wire _guard25191 = cond_wire569_out;
wire _guard25192 = _guard25190 & _guard25191;
wire _guard25193 = fsm_out == 1'd0;
wire _guard25194 = _guard25192 & _guard25193;
wire _guard25195 = _guard25189 | _guard25194;
wire _guard25196 = early_reset_static_par0_go_out;
wire _guard25197 = _guard25195 & _guard25196;
wire _guard25198 = cond_wire536_out;
wire _guard25199 = early_reset_static_par0_go_out;
wire _guard25200 = _guard25198 & _guard25199;
wire _guard25201 = cond_wire536_out;
wire _guard25202 = early_reset_static_par0_go_out;
wire _guard25203 = _guard25201 & _guard25202;
wire _guard25204 = cond_wire621_out;
wire _guard25205 = early_reset_static_par0_go_out;
wire _guard25206 = _guard25204 & _guard25205;
wire _guard25207 = cond_wire621_out;
wire _guard25208 = early_reset_static_par0_go_out;
wire _guard25209 = _guard25207 & _guard25208;
wire _guard25210 = cond_wire568_out;
wire _guard25211 = early_reset_static_par0_go_out;
wire _guard25212 = _guard25210 & _guard25211;
wire _guard25213 = cond_wire568_out;
wire _guard25214 = early_reset_static_par0_go_out;
wire _guard25215 = _guard25213 & _guard25214;
wire _guard25216 = cond_wire694_out;
wire _guard25217 = early_reset_static_par0_go_out;
wire _guard25218 = _guard25216 & _guard25217;
wire _guard25219 = cond_wire694_out;
wire _guard25220 = early_reset_static_par0_go_out;
wire _guard25221 = _guard25219 & _guard25220;
wire _guard25222 = cond_wire729_out;
wire _guard25223 = early_reset_static_par0_go_out;
wire _guard25224 = _guard25222 & _guard25223;
wire _guard25225 = cond_wire729_out;
wire _guard25226 = early_reset_static_par0_go_out;
wire _guard25227 = _guard25225 & _guard25226;
wire _guard25228 = cond_wire805_out;
wire _guard25229 = early_reset_static_par0_go_out;
wire _guard25230 = _guard25228 & _guard25229;
wire _guard25231 = cond_wire803_out;
wire _guard25232 = early_reset_static_par0_go_out;
wire _guard25233 = _guard25231 & _guard25232;
wire _guard25234 = fsm_out == 1'd0;
wire _guard25235 = cond_wire803_out;
wire _guard25236 = _guard25234 & _guard25235;
wire _guard25237 = fsm_out == 1'd0;
wire _guard25238 = _guard25236 & _guard25237;
wire _guard25239 = fsm_out == 1'd0;
wire _guard25240 = cond_wire805_out;
wire _guard25241 = _guard25239 & _guard25240;
wire _guard25242 = fsm_out == 1'd0;
wire _guard25243 = _guard25241 & _guard25242;
wire _guard25244 = _guard25238 | _guard25243;
wire _guard25245 = early_reset_static_par0_go_out;
wire _guard25246 = _guard25244 & _guard25245;
wire _guard25247 = fsm_out == 1'd0;
wire _guard25248 = cond_wire803_out;
wire _guard25249 = _guard25247 & _guard25248;
wire _guard25250 = fsm_out == 1'd0;
wire _guard25251 = _guard25249 & _guard25250;
wire _guard25252 = fsm_out == 1'd0;
wire _guard25253 = cond_wire805_out;
wire _guard25254 = _guard25252 & _guard25253;
wire _guard25255 = fsm_out == 1'd0;
wire _guard25256 = _guard25254 & _guard25255;
wire _guard25257 = _guard25251 | _guard25256;
wire _guard25258 = early_reset_static_par0_go_out;
wire _guard25259 = _guard25257 & _guard25258;
wire _guard25260 = fsm_out == 1'd0;
wire _guard25261 = cond_wire803_out;
wire _guard25262 = _guard25260 & _guard25261;
wire _guard25263 = fsm_out == 1'd0;
wire _guard25264 = _guard25262 & _guard25263;
wire _guard25265 = fsm_out == 1'd0;
wire _guard25266 = cond_wire805_out;
wire _guard25267 = _guard25265 & _guard25266;
wire _guard25268 = fsm_out == 1'd0;
wire _guard25269 = _guard25267 & _guard25268;
wire _guard25270 = _guard25264 | _guard25269;
wire _guard25271 = early_reset_static_par0_go_out;
wire _guard25272 = _guard25270 & _guard25271;
wire _guard25273 = cond_wire829_out;
wire _guard25274 = early_reset_static_par0_go_out;
wire _guard25275 = _guard25273 & _guard25274;
wire _guard25276 = cond_wire827_out;
wire _guard25277 = early_reset_static_par0_go_out;
wire _guard25278 = _guard25276 & _guard25277;
wire _guard25279 = fsm_out == 1'd0;
wire _guard25280 = cond_wire827_out;
wire _guard25281 = _guard25279 & _guard25280;
wire _guard25282 = fsm_out == 1'd0;
wire _guard25283 = _guard25281 & _guard25282;
wire _guard25284 = fsm_out == 1'd0;
wire _guard25285 = cond_wire829_out;
wire _guard25286 = _guard25284 & _guard25285;
wire _guard25287 = fsm_out == 1'd0;
wire _guard25288 = _guard25286 & _guard25287;
wire _guard25289 = _guard25283 | _guard25288;
wire _guard25290 = early_reset_static_par0_go_out;
wire _guard25291 = _guard25289 & _guard25290;
wire _guard25292 = fsm_out == 1'd0;
wire _guard25293 = cond_wire827_out;
wire _guard25294 = _guard25292 & _guard25293;
wire _guard25295 = fsm_out == 1'd0;
wire _guard25296 = _guard25294 & _guard25295;
wire _guard25297 = fsm_out == 1'd0;
wire _guard25298 = cond_wire829_out;
wire _guard25299 = _guard25297 & _guard25298;
wire _guard25300 = fsm_out == 1'd0;
wire _guard25301 = _guard25299 & _guard25300;
wire _guard25302 = _guard25296 | _guard25301;
wire _guard25303 = early_reset_static_par0_go_out;
wire _guard25304 = _guard25302 & _guard25303;
wire _guard25305 = fsm_out == 1'd0;
wire _guard25306 = cond_wire827_out;
wire _guard25307 = _guard25305 & _guard25306;
wire _guard25308 = fsm_out == 1'd0;
wire _guard25309 = _guard25307 & _guard25308;
wire _guard25310 = fsm_out == 1'd0;
wire _guard25311 = cond_wire829_out;
wire _guard25312 = _guard25310 & _guard25311;
wire _guard25313 = fsm_out == 1'd0;
wire _guard25314 = _guard25312 & _guard25313;
wire _guard25315 = _guard25309 | _guard25314;
wire _guard25316 = early_reset_static_par0_go_out;
wire _guard25317 = _guard25315 & _guard25316;
wire _guard25318 = cond_wire767_out;
wire _guard25319 = early_reset_static_par0_go_out;
wire _guard25320 = _guard25318 & _guard25319;
wire _guard25321 = cond_wire767_out;
wire _guard25322 = early_reset_static_par0_go_out;
wire _guard25323 = _guard25321 & _guard25322;
wire _guard25324 = cond_wire853_out;
wire _guard25325 = early_reset_static_par0_go_out;
wire _guard25326 = _guard25324 & _guard25325;
wire _guard25327 = cond_wire851_out;
wire _guard25328 = early_reset_static_par0_go_out;
wire _guard25329 = _guard25327 & _guard25328;
wire _guard25330 = fsm_out == 1'd0;
wire _guard25331 = cond_wire851_out;
wire _guard25332 = _guard25330 & _guard25331;
wire _guard25333 = fsm_out == 1'd0;
wire _guard25334 = _guard25332 & _guard25333;
wire _guard25335 = fsm_out == 1'd0;
wire _guard25336 = cond_wire853_out;
wire _guard25337 = _guard25335 & _guard25336;
wire _guard25338 = fsm_out == 1'd0;
wire _guard25339 = _guard25337 & _guard25338;
wire _guard25340 = _guard25334 | _guard25339;
wire _guard25341 = early_reset_static_par0_go_out;
wire _guard25342 = _guard25340 & _guard25341;
wire _guard25343 = fsm_out == 1'd0;
wire _guard25344 = cond_wire851_out;
wire _guard25345 = _guard25343 & _guard25344;
wire _guard25346 = fsm_out == 1'd0;
wire _guard25347 = _guard25345 & _guard25346;
wire _guard25348 = fsm_out == 1'd0;
wire _guard25349 = cond_wire853_out;
wire _guard25350 = _guard25348 & _guard25349;
wire _guard25351 = fsm_out == 1'd0;
wire _guard25352 = _guard25350 & _guard25351;
wire _guard25353 = _guard25347 | _guard25352;
wire _guard25354 = early_reset_static_par0_go_out;
wire _guard25355 = _guard25353 & _guard25354;
wire _guard25356 = fsm_out == 1'd0;
wire _guard25357 = cond_wire851_out;
wire _guard25358 = _guard25356 & _guard25357;
wire _guard25359 = fsm_out == 1'd0;
wire _guard25360 = _guard25358 & _guard25359;
wire _guard25361 = fsm_out == 1'd0;
wire _guard25362 = cond_wire853_out;
wire _guard25363 = _guard25361 & _guard25362;
wire _guard25364 = fsm_out == 1'd0;
wire _guard25365 = _guard25363 & _guard25364;
wire _guard25366 = _guard25360 | _guard25365;
wire _guard25367 = early_reset_static_par0_go_out;
wire _guard25368 = _guard25366 & _guard25367;
wire _guard25369 = cond_wire870_out;
wire _guard25370 = early_reset_static_par0_go_out;
wire _guard25371 = _guard25369 & _guard25370;
wire _guard25372 = cond_wire868_out;
wire _guard25373 = early_reset_static_par0_go_out;
wire _guard25374 = _guard25372 & _guard25373;
wire _guard25375 = fsm_out == 1'd0;
wire _guard25376 = cond_wire868_out;
wire _guard25377 = _guard25375 & _guard25376;
wire _guard25378 = fsm_out == 1'd0;
wire _guard25379 = _guard25377 & _guard25378;
wire _guard25380 = fsm_out == 1'd0;
wire _guard25381 = cond_wire870_out;
wire _guard25382 = _guard25380 & _guard25381;
wire _guard25383 = fsm_out == 1'd0;
wire _guard25384 = _guard25382 & _guard25383;
wire _guard25385 = _guard25379 | _guard25384;
wire _guard25386 = early_reset_static_par0_go_out;
wire _guard25387 = _guard25385 & _guard25386;
wire _guard25388 = fsm_out == 1'd0;
wire _guard25389 = cond_wire868_out;
wire _guard25390 = _guard25388 & _guard25389;
wire _guard25391 = fsm_out == 1'd0;
wire _guard25392 = _guard25390 & _guard25391;
wire _guard25393 = fsm_out == 1'd0;
wire _guard25394 = cond_wire870_out;
wire _guard25395 = _guard25393 & _guard25394;
wire _guard25396 = fsm_out == 1'd0;
wire _guard25397 = _guard25395 & _guard25396;
wire _guard25398 = _guard25392 | _guard25397;
wire _guard25399 = early_reset_static_par0_go_out;
wire _guard25400 = _guard25398 & _guard25399;
wire _guard25401 = fsm_out == 1'd0;
wire _guard25402 = cond_wire868_out;
wire _guard25403 = _guard25401 & _guard25402;
wire _guard25404 = fsm_out == 1'd0;
wire _guard25405 = _guard25403 & _guard25404;
wire _guard25406 = fsm_out == 1'd0;
wire _guard25407 = cond_wire870_out;
wire _guard25408 = _guard25406 & _guard25407;
wire _guard25409 = fsm_out == 1'd0;
wire _guard25410 = _guard25408 & _guard25409;
wire _guard25411 = _guard25405 | _guard25410;
wire _guard25412 = early_reset_static_par0_go_out;
wire _guard25413 = _guard25411 & _guard25412;
wire _guard25414 = cond_wire804_out;
wire _guard25415 = early_reset_static_par0_go_out;
wire _guard25416 = _guard25414 & _guard25415;
wire _guard25417 = cond_wire804_out;
wire _guard25418 = early_reset_static_par0_go_out;
wire _guard25419 = _guard25417 & _guard25418;
wire _guard25420 = cond_wire905_out;
wire _guard25421 = early_reset_static_par0_go_out;
wire _guard25422 = _guard25420 & _guard25421;
wire _guard25423 = cond_wire905_out;
wire _guard25424 = early_reset_static_par0_go_out;
wire _guard25425 = _guard25423 & _guard25424;
wire _guard25426 = cond_wire901_out;
wire _guard25427 = early_reset_static_par0_go_out;
wire _guard25428 = _guard25426 & _guard25427;
wire _guard25429 = cond_wire901_out;
wire _guard25430 = early_reset_static_par0_go_out;
wire _guard25431 = _guard25429 & _guard25430;
wire _guard25432 = cond_wire971_out;
wire _guard25433 = early_reset_static_par0_go_out;
wire _guard25434 = _guard25432 & _guard25433;
wire _guard25435 = cond_wire969_out;
wire _guard25436 = early_reset_static_par0_go_out;
wire _guard25437 = _guard25435 & _guard25436;
wire _guard25438 = fsm_out == 1'd0;
wire _guard25439 = cond_wire969_out;
wire _guard25440 = _guard25438 & _guard25439;
wire _guard25441 = fsm_out == 1'd0;
wire _guard25442 = _guard25440 & _guard25441;
wire _guard25443 = fsm_out == 1'd0;
wire _guard25444 = cond_wire971_out;
wire _guard25445 = _guard25443 & _guard25444;
wire _guard25446 = fsm_out == 1'd0;
wire _guard25447 = _guard25445 & _guard25446;
wire _guard25448 = _guard25442 | _guard25447;
wire _guard25449 = early_reset_static_par0_go_out;
wire _guard25450 = _guard25448 & _guard25449;
wire _guard25451 = fsm_out == 1'd0;
wire _guard25452 = cond_wire969_out;
wire _guard25453 = _guard25451 & _guard25452;
wire _guard25454 = fsm_out == 1'd0;
wire _guard25455 = _guard25453 & _guard25454;
wire _guard25456 = fsm_out == 1'd0;
wire _guard25457 = cond_wire971_out;
wire _guard25458 = _guard25456 & _guard25457;
wire _guard25459 = fsm_out == 1'd0;
wire _guard25460 = _guard25458 & _guard25459;
wire _guard25461 = _guard25455 | _guard25460;
wire _guard25462 = early_reset_static_par0_go_out;
wire _guard25463 = _guard25461 & _guard25462;
wire _guard25464 = fsm_out == 1'd0;
wire _guard25465 = cond_wire969_out;
wire _guard25466 = _guard25464 & _guard25465;
wire _guard25467 = fsm_out == 1'd0;
wire _guard25468 = _guard25466 & _guard25467;
wire _guard25469 = fsm_out == 1'd0;
wire _guard25470 = cond_wire971_out;
wire _guard25471 = _guard25469 & _guard25470;
wire _guard25472 = fsm_out == 1'd0;
wire _guard25473 = _guard25471 & _guard25472;
wire _guard25474 = _guard25468 | _guard25473;
wire _guard25475 = early_reset_static_par0_go_out;
wire _guard25476 = _guard25474 & _guard25475;
wire _guard25477 = cond_wire913_out;
wire _guard25478 = early_reset_static_par0_go_out;
wire _guard25479 = _guard25477 & _guard25478;
wire _guard25480 = cond_wire913_out;
wire _guard25481 = early_reset_static_par0_go_out;
wire _guard25482 = _guard25480 & _guard25481;
wire _guard25483 = cond_wire999_out;
wire _guard25484 = early_reset_static_par0_go_out;
wire _guard25485 = _guard25483 & _guard25484;
wire _guard25486 = cond_wire999_out;
wire _guard25487 = early_reset_static_par0_go_out;
wire _guard25488 = _guard25486 & _guard25487;
wire _guard25489 = cond_wire1024_out;
wire _guard25490 = early_reset_static_par0_go_out;
wire _guard25491 = _guard25489 & _guard25490;
wire _guard25492 = cond_wire1022_out;
wire _guard25493 = early_reset_static_par0_go_out;
wire _guard25494 = _guard25492 & _guard25493;
wire _guard25495 = fsm_out == 1'd0;
wire _guard25496 = cond_wire1022_out;
wire _guard25497 = _guard25495 & _guard25496;
wire _guard25498 = fsm_out == 1'd0;
wire _guard25499 = _guard25497 & _guard25498;
wire _guard25500 = fsm_out == 1'd0;
wire _guard25501 = cond_wire1024_out;
wire _guard25502 = _guard25500 & _guard25501;
wire _guard25503 = fsm_out == 1'd0;
wire _guard25504 = _guard25502 & _guard25503;
wire _guard25505 = _guard25499 | _guard25504;
wire _guard25506 = early_reset_static_par0_go_out;
wire _guard25507 = _guard25505 & _guard25506;
wire _guard25508 = fsm_out == 1'd0;
wire _guard25509 = cond_wire1022_out;
wire _guard25510 = _guard25508 & _guard25509;
wire _guard25511 = fsm_out == 1'd0;
wire _guard25512 = _guard25510 & _guard25511;
wire _guard25513 = fsm_out == 1'd0;
wire _guard25514 = cond_wire1024_out;
wire _guard25515 = _guard25513 & _guard25514;
wire _guard25516 = fsm_out == 1'd0;
wire _guard25517 = _guard25515 & _guard25516;
wire _guard25518 = _guard25512 | _guard25517;
wire _guard25519 = early_reset_static_par0_go_out;
wire _guard25520 = _guard25518 & _guard25519;
wire _guard25521 = fsm_out == 1'd0;
wire _guard25522 = cond_wire1022_out;
wire _guard25523 = _guard25521 & _guard25522;
wire _guard25524 = fsm_out == 1'd0;
wire _guard25525 = _guard25523 & _guard25524;
wire _guard25526 = fsm_out == 1'd0;
wire _guard25527 = cond_wire1024_out;
wire _guard25528 = _guard25526 & _guard25527;
wire _guard25529 = fsm_out == 1'd0;
wire _guard25530 = _guard25528 & _guard25529;
wire _guard25531 = _guard25525 | _guard25530;
wire _guard25532 = early_reset_static_par0_go_out;
wire _guard25533 = _guard25531 & _guard25532;
wire _guard25534 = cond_wire958_out;
wire _guard25535 = early_reset_static_par0_go_out;
wire _guard25536 = _guard25534 & _guard25535;
wire _guard25537 = cond_wire958_out;
wire _guard25538 = early_reset_static_par0_go_out;
wire _guard25539 = _guard25537 & _guard25538;
wire _guard25540 = cond_wire1019_out;
wire _guard25541 = early_reset_static_par0_go_out;
wire _guard25542 = _guard25540 & _guard25541;
wire _guard25543 = cond_wire1019_out;
wire _guard25544 = early_reset_static_par0_go_out;
wire _guard25545 = _guard25543 & _guard25544;
wire _guard25546 = cond_wire1035_out;
wire _guard25547 = early_reset_static_par0_go_out;
wire _guard25548 = _guard25546 & _guard25547;
wire _guard25549 = cond_wire1035_out;
wire _guard25550 = early_reset_static_par0_go_out;
wire _guard25551 = _guard25549 & _guard25550;
wire _guard25552 = cond_wire1039_out;
wire _guard25553 = early_reset_static_par0_go_out;
wire _guard25554 = _guard25552 & _guard25553;
wire _guard25555 = cond_wire1039_out;
wire _guard25556 = early_reset_static_par0_go_out;
wire _guard25557 = _guard25555 & _guard25556;
wire _guard25558 = cond_wire39_out;
wire _guard25559 = early_reset_static_par0_go_out;
wire _guard25560 = _guard25558 & _guard25559;
wire _guard25561 = cond_wire39_out;
wire _guard25562 = early_reset_static_par0_go_out;
wire _guard25563 = _guard25561 & _guard25562;
wire _guard25564 = cond_wire144_out;
wire _guard25565 = early_reset_static_par0_go_out;
wire _guard25566 = _guard25564 & _guard25565;
wire _guard25567 = cond_wire144_out;
wire _guard25568 = early_reset_static_par0_go_out;
wire _guard25569 = _guard25567 & _guard25568;
wire _guard25570 = fsm0_out == 6'd0;
wire _guard25571 = early_reset_static_seq_go_out;
wire _guard25572 = _guard25570 & _guard25571;
wire _guard25573 = cond_wire339_out;
wire _guard25574 = early_reset_static_par0_go_out;
wire _guard25575 = _guard25573 & _guard25574;
wire _guard25576 = _guard25572 | _guard25575;
wire _guard25577 = fsm0_out == 6'd0;
wire _guard25578 = early_reset_static_seq_go_out;
wire _guard25579 = _guard25577 & _guard25578;
wire _guard25580 = cond_wire339_out;
wire _guard25581 = early_reset_static_par0_go_out;
wire _guard25582 = _guard25580 & _guard25581;
wire _guard25583 = cond_wire404_out;
wire _guard25584 = early_reset_static_par0_go_out;
wire _guard25585 = _guard25583 & _guard25584;
wire _guard25586 = cond_wire404_out;
wire _guard25587 = early_reset_static_par0_go_out;
wire _guard25588 = _guard25586 & _guard25587;
wire _guard25589 = fsm0_out == 6'd0;
wire _guard25590 = early_reset_static_seq_go_out;
wire _guard25591 = _guard25589 & _guard25590;
wire _guard25592 = cond_wire534_out;
wire _guard25593 = early_reset_static_par0_go_out;
wire _guard25594 = _guard25592 & _guard25593;
wire _guard25595 = _guard25591 | _guard25594;
wire _guard25596 = fsm0_out == 6'd0;
wire _guard25597 = early_reset_static_seq_go_out;
wire _guard25598 = _guard25596 & _guard25597;
wire _guard25599 = cond_wire534_out;
wire _guard25600 = early_reset_static_par0_go_out;
wire _guard25601 = _guard25599 & _guard25600;
wire _guard25602 = early_reset_static_par0_go_out;
wire _guard25603 = early_reset_static_par0_go_out;
wire _guard25604 = early_reset_static_par0_go_out;
wire _guard25605 = early_reset_static_par0_go_out;
wire _guard25606 = early_reset_static_par0_go_out;
wire _guard25607 = early_reset_static_par0_go_out;
wire _guard25608 = early_reset_static_par0_go_out;
wire _guard25609 = early_reset_static_par0_go_out;
wire _guard25610 = early_reset_static_par0_go_out;
wire _guard25611 = early_reset_static_par0_go_out;
wire _guard25612 = fsm0_out == 6'd0;
wire _guard25613 = early_reset_static_seq_go_out;
wire _guard25614 = _guard25612 & _guard25613;
wire _guard25615 = early_reset_static_par0_go_out;
wire _guard25616 = _guard25614 | _guard25615;
wire _guard25617 = early_reset_static_par0_go_out;
wire _guard25618 = fsm0_out == 6'd0;
wire _guard25619 = early_reset_static_seq_go_out;
wire _guard25620 = _guard25618 & _guard25619;
wire _guard25621 = early_reset_static_par0_go_out;
wire _guard25622 = early_reset_static_par0_go_out;
wire _guard25623 = early_reset_static_par0_go_out;
wire _guard25624 = early_reset_static_par0_go_out;
wire _guard25625 = fsm0_out == 6'd0;
wire _guard25626 = early_reset_static_seq_go_out;
wire _guard25627 = _guard25625 & _guard25626;
wire _guard25628 = early_reset_static_par0_go_out;
wire _guard25629 = _guard25627 | _guard25628;
wire _guard25630 = early_reset_static_par0_go_out;
wire _guard25631 = fsm0_out == 6'd0;
wire _guard25632 = early_reset_static_seq_go_out;
wire _guard25633 = _guard25631 & _guard25632;
wire _guard25634 = early_reset_static_par0_go_out;
wire _guard25635 = early_reset_static_par0_go_out;
wire _guard25636 = fsm0_out == 6'd0;
wire _guard25637 = early_reset_static_seq_go_out;
wire _guard25638 = _guard25636 & _guard25637;
wire _guard25639 = early_reset_static_par0_go_out;
wire _guard25640 = _guard25638 | _guard25639;
wire _guard25641 = fsm0_out == 6'd0;
wire _guard25642 = early_reset_static_seq_go_out;
wire _guard25643 = _guard25641 & _guard25642;
wire _guard25644 = early_reset_static_par0_go_out;
wire _guard25645 = fsm0_out == 6'd0;
wire _guard25646 = early_reset_static_seq_go_out;
wire _guard25647 = _guard25645 & _guard25646;
wire _guard25648 = early_reset_static_par0_go_out;
wire _guard25649 = _guard25647 | _guard25648;
wire _guard25650 = fsm0_out == 6'd0;
wire _guard25651 = early_reset_static_seq_go_out;
wire _guard25652 = _guard25650 & _guard25651;
wire _guard25653 = early_reset_static_par0_go_out;
wire _guard25654 = early_reset_static_par0_go_out;
wire _guard25655 = early_reset_static_par0_go_out;
wire _guard25656 = early_reset_static_par0_go_out;
wire _guard25657 = early_reset_static_par0_go_out;
wire _guard25658 = fsm0_out == 6'd0;
wire _guard25659 = early_reset_static_seq_go_out;
wire _guard25660 = _guard25658 & _guard25659;
wire _guard25661 = early_reset_static_par0_go_out;
wire _guard25662 = _guard25660 | _guard25661;
wire _guard25663 = early_reset_static_par0_go_out;
wire _guard25664 = fsm0_out == 6'd0;
wire _guard25665 = early_reset_static_seq_go_out;
wire _guard25666 = _guard25664 & _guard25665;
wire _guard25667 = early_reset_static_par0_go_out;
wire _guard25668 = ~_guard0;
wire _guard25669 = early_reset_static_par0_go_out;
wire _guard25670 = _guard25668 & _guard25669;
wire _guard25671 = early_reset_static_par0_go_out;
wire _guard25672 = ~_guard0;
wire _guard25673 = early_reset_static_par0_go_out;
wire _guard25674 = _guard25672 & _guard25673;
wire _guard25675 = early_reset_static_par0_go_out;
wire _guard25676 = early_reset_static_par0_go_out;
wire _guard25677 = early_reset_static_par0_go_out;
wire _guard25678 = early_reset_static_par0_go_out;
wire _guard25679 = early_reset_static_par0_go_out;
wire _guard25680 = ~_guard0;
wire _guard25681 = early_reset_static_par0_go_out;
wire _guard25682 = _guard25680 & _guard25681;
wire _guard25683 = early_reset_static_par0_go_out;
wire _guard25684 = early_reset_static_par0_go_out;
wire _guard25685 = early_reset_static_par0_go_out;
wire _guard25686 = ~_guard0;
wire _guard25687 = early_reset_static_par0_go_out;
wire _guard25688 = _guard25686 & _guard25687;
wire _guard25689 = early_reset_static_par0_go_out;
wire _guard25690 = ~_guard0;
wire _guard25691 = early_reset_static_par0_go_out;
wire _guard25692 = _guard25690 & _guard25691;
wire _guard25693 = early_reset_static_par0_go_out;
wire _guard25694 = early_reset_static_par0_go_out;
wire _guard25695 = early_reset_static_par0_go_out;
wire _guard25696 = ~_guard0;
wire _guard25697 = early_reset_static_par0_go_out;
wire _guard25698 = _guard25696 & _guard25697;
wire _guard25699 = early_reset_static_par0_go_out;
wire _guard25700 = early_reset_static_par0_go_out;
wire _guard25701 = ~_guard0;
wire _guard25702 = early_reset_static_par0_go_out;
wire _guard25703 = _guard25701 & _guard25702;
wire _guard25704 = early_reset_static_par0_go_out;
wire _guard25705 = early_reset_static_par0_go_out;
wire _guard25706 = early_reset_static_par0_go_out;
wire _guard25707 = early_reset_static_par0_go_out;
wire _guard25708 = early_reset_static_par0_go_out;
wire _guard25709 = ~_guard0;
wire _guard25710 = early_reset_static_par0_go_out;
wire _guard25711 = _guard25709 & _guard25710;
wire _guard25712 = early_reset_static_par0_go_out;
wire _guard25713 = ~_guard0;
wire _guard25714 = early_reset_static_par0_go_out;
wire _guard25715 = _guard25713 & _guard25714;
wire _guard25716 = early_reset_static_par0_go_out;
wire _guard25717 = early_reset_static_par0_go_out;
wire _guard25718 = ~_guard0;
wire _guard25719 = early_reset_static_par0_go_out;
wire _guard25720 = _guard25718 & _guard25719;
wire _guard25721 = ~_guard0;
wire _guard25722 = early_reset_static_par0_go_out;
wire _guard25723 = _guard25721 & _guard25722;
wire _guard25724 = early_reset_static_par0_go_out;
wire _guard25725 = early_reset_static_par0_go_out;
wire _guard25726 = early_reset_static_par0_go_out;
wire _guard25727 = ~_guard0;
wire _guard25728 = early_reset_static_par0_go_out;
wire _guard25729 = _guard25727 & _guard25728;
wire _guard25730 = early_reset_static_par0_go_out;
wire _guard25731 = ~_guard0;
wire _guard25732 = early_reset_static_par0_go_out;
wire _guard25733 = _guard25731 & _guard25732;
wire _guard25734 = early_reset_static_par0_go_out;
wire _guard25735 = ~_guard0;
wire _guard25736 = early_reset_static_par0_go_out;
wire _guard25737 = _guard25735 & _guard25736;
wire _guard25738 = early_reset_static_par0_go_out;
wire _guard25739 = ~_guard0;
wire _guard25740 = early_reset_static_par0_go_out;
wire _guard25741 = _guard25739 & _guard25740;
wire _guard25742 = early_reset_static_par0_go_out;
wire _guard25743 = ~_guard0;
wire _guard25744 = early_reset_static_par0_go_out;
wire _guard25745 = _guard25743 & _guard25744;
wire _guard25746 = early_reset_static_par0_go_out;
wire _guard25747 = early_reset_static_par0_go_out;
wire _guard25748 = early_reset_static_par0_go_out;
wire _guard25749 = early_reset_static_par0_go_out;
wire _guard25750 = early_reset_static_par0_go_out;
wire _guard25751 = early_reset_static_par0_go_out;
wire _guard25752 = ~_guard0;
wire _guard25753 = early_reset_static_par0_go_out;
wire _guard25754 = _guard25752 & _guard25753;
wire _guard25755 = ~_guard0;
wire _guard25756 = early_reset_static_par0_go_out;
wire _guard25757 = _guard25755 & _guard25756;
wire _guard25758 = early_reset_static_par0_go_out;
wire _guard25759 = early_reset_static_par0_go_out;
wire _guard25760 = early_reset_static_par0_go_out;
wire _guard25761 = early_reset_static_par0_go_out;
wire _guard25762 = early_reset_static_par0_go_out;
wire _guard25763 = ~_guard0;
wire _guard25764 = early_reset_static_par0_go_out;
wire _guard25765 = _guard25763 & _guard25764;
wire _guard25766 = early_reset_static_par0_go_out;
wire _guard25767 = early_reset_static_par0_go_out;
wire _guard25768 = ~_guard0;
wire _guard25769 = early_reset_static_par0_go_out;
wire _guard25770 = _guard25768 & _guard25769;
wire _guard25771 = ~_guard0;
wire _guard25772 = early_reset_static_par0_go_out;
wire _guard25773 = _guard25771 & _guard25772;
wire _guard25774 = early_reset_static_par0_go_out;
wire _guard25775 = early_reset_static_par0_go_out;
wire _guard25776 = early_reset_static_par0_go_out;
wire _guard25777 = early_reset_static_par0_go_out;
wire _guard25778 = ~_guard0;
wire _guard25779 = early_reset_static_par0_go_out;
wire _guard25780 = _guard25778 & _guard25779;
wire _guard25781 = early_reset_static_par0_go_out;
wire _guard25782 = early_reset_static_par0_go_out;
wire _guard25783 = early_reset_static_par0_go_out;
wire _guard25784 = ~_guard0;
wire _guard25785 = early_reset_static_par0_go_out;
wire _guard25786 = _guard25784 & _guard25785;
wire _guard25787 = early_reset_static_par0_go_out;
wire _guard25788 = ~_guard0;
wire _guard25789 = early_reset_static_par0_go_out;
wire _guard25790 = _guard25788 & _guard25789;
wire _guard25791 = ~_guard0;
wire _guard25792 = early_reset_static_par0_go_out;
wire _guard25793 = _guard25791 & _guard25792;
wire _guard25794 = early_reset_static_par0_go_out;
wire _guard25795 = early_reset_static_par0_go_out;
wire _guard25796 = early_reset_static_par0_go_out;
wire _guard25797 = ~_guard0;
wire _guard25798 = early_reset_static_par0_go_out;
wire _guard25799 = _guard25797 & _guard25798;
wire _guard25800 = early_reset_static_par0_go_out;
wire _guard25801 = ~_guard0;
wire _guard25802 = early_reset_static_par0_go_out;
wire _guard25803 = _guard25801 & _guard25802;
wire _guard25804 = early_reset_static_par0_go_out;
wire _guard25805 = ~_guard0;
wire _guard25806 = early_reset_static_par0_go_out;
wire _guard25807 = _guard25805 & _guard25806;
wire _guard25808 = early_reset_static_par0_go_out;
wire _guard25809 = early_reset_static_par0_go_out;
wire _guard25810 = ~_guard0;
wire _guard25811 = early_reset_static_par0_go_out;
wire _guard25812 = _guard25810 & _guard25811;
wire _guard25813 = early_reset_static_par0_go_out;
wire _guard25814 = early_reset_static_par0_go_out;
wire _guard25815 = early_reset_static_par0_go_out;
wire _guard25816 = early_reset_static_par0_go_out;
wire _guard25817 = ~_guard0;
wire _guard25818 = early_reset_static_par0_go_out;
wire _guard25819 = _guard25817 & _guard25818;
wire _guard25820 = early_reset_static_par0_go_out;
wire _guard25821 = early_reset_static_par0_go_out;
wire _guard25822 = ~_guard0;
wire _guard25823 = early_reset_static_par0_go_out;
wire _guard25824 = _guard25822 & _guard25823;
wire _guard25825 = early_reset_static_par0_go_out;
wire _guard25826 = ~_guard0;
wire _guard25827 = early_reset_static_par0_go_out;
wire _guard25828 = _guard25826 & _guard25827;
wire _guard25829 = early_reset_static_par0_go_out;
wire _guard25830 = ~_guard0;
wire _guard25831 = early_reset_static_par0_go_out;
wire _guard25832 = _guard25830 & _guard25831;
wire _guard25833 = ~_guard0;
wire _guard25834 = early_reset_static_par0_go_out;
wire _guard25835 = _guard25833 & _guard25834;
wire _guard25836 = early_reset_static_par0_go_out;
wire _guard25837 = ~_guard0;
wire _guard25838 = early_reset_static_par0_go_out;
wire _guard25839 = _guard25837 & _guard25838;
wire _guard25840 = early_reset_static_par0_go_out;
wire _guard25841 = ~_guard0;
wire _guard25842 = early_reset_static_par0_go_out;
wire _guard25843 = _guard25841 & _guard25842;
wire _guard25844 = early_reset_static_par0_go_out;
wire _guard25845 = ~_guard0;
wire _guard25846 = early_reset_static_par0_go_out;
wire _guard25847 = _guard25845 & _guard25846;
wire _guard25848 = early_reset_static_par0_go_out;
wire _guard25849 = early_reset_static_par0_go_out;
wire _guard25850 = ~_guard0;
wire _guard25851 = early_reset_static_par0_go_out;
wire _guard25852 = _guard25850 & _guard25851;
wire _guard25853 = ~_guard0;
wire _guard25854 = early_reset_static_par0_go_out;
wire _guard25855 = _guard25853 & _guard25854;
wire _guard25856 = early_reset_static_par0_go_out;
wire _guard25857 = early_reset_static_par0_go_out;
wire _guard25858 = early_reset_static_par0_go_out;
wire _guard25859 = ~_guard0;
wire _guard25860 = early_reset_static_par0_go_out;
wire _guard25861 = _guard25859 & _guard25860;
wire _guard25862 = early_reset_static_par0_go_out;
wire _guard25863 = early_reset_static_par0_go_out;
wire _guard25864 = early_reset_static_par0_go_out;
wire _guard25865 = early_reset_static_par0_go_out;
wire _guard25866 = early_reset_static_par0_go_out;
wire _guard25867 = early_reset_static_par0_go_out;
wire _guard25868 = early_reset_static_par0_go_out;
wire _guard25869 = early_reset_static_par0_go_out;
wire _guard25870 = early_reset_static_par0_go_out;
wire _guard25871 = early_reset_static_par0_go_out;
wire _guard25872 = ~_guard0;
wire _guard25873 = early_reset_static_par0_go_out;
wire _guard25874 = _guard25872 & _guard25873;
wire _guard25875 = early_reset_static_par0_go_out;
wire _guard25876 = early_reset_static_par0_go_out;
wire _guard25877 = early_reset_static_par0_go_out;
wire _guard25878 = early_reset_static_par0_go_out;
wire _guard25879 = early_reset_static_par0_go_out;
wire _guard25880 = ~_guard0;
wire _guard25881 = early_reset_static_par0_go_out;
wire _guard25882 = _guard25880 & _guard25881;
wire _guard25883 = early_reset_static_par0_go_out;
wire _guard25884 = early_reset_static_par0_go_out;
wire _guard25885 = early_reset_static_par0_go_out;
wire _guard25886 = early_reset_static_par0_go_out;
wire _guard25887 = ~_guard0;
wire _guard25888 = early_reset_static_par0_go_out;
wire _guard25889 = _guard25887 & _guard25888;
wire _guard25890 = early_reset_static_par0_go_out;
wire _guard25891 = early_reset_static_par0_go_out;
wire _guard25892 = early_reset_static_par0_go_out;
wire _guard25893 = early_reset_static_par0_go_out;
wire _guard25894 = early_reset_static_par0_go_out;
wire _guard25895 = ~_guard0;
wire _guard25896 = early_reset_static_par0_go_out;
wire _guard25897 = _guard25895 & _guard25896;
wire _guard25898 = early_reset_static_par0_go_out;
wire _guard25899 = early_reset_static_par0_go_out;
wire _guard25900 = early_reset_static_par0_go_out;
wire _guard25901 = early_reset_static_par0_go_out;
wire _guard25902 = early_reset_static_par0_go_out;
wire _guard25903 = ~_guard0;
wire _guard25904 = early_reset_static_par0_go_out;
wire _guard25905 = _guard25903 & _guard25904;
wire _guard25906 = early_reset_static_par0_go_out;
wire _guard25907 = ~_guard0;
wire _guard25908 = early_reset_static_par0_go_out;
wire _guard25909 = _guard25907 & _guard25908;
wire _guard25910 = early_reset_static_par0_go_out;
wire _guard25911 = ~_guard0;
wire _guard25912 = early_reset_static_par0_go_out;
wire _guard25913 = _guard25911 & _guard25912;
wire _guard25914 = early_reset_static_par0_go_out;
wire _guard25915 = early_reset_static_par0_go_out;
wire _guard25916 = early_reset_static_par0_go_out;
wire _guard25917 = ~_guard0;
wire _guard25918 = early_reset_static_par0_go_out;
wire _guard25919 = _guard25917 & _guard25918;
wire _guard25920 = early_reset_static_par0_go_out;
wire _guard25921 = early_reset_static_par0_go_out;
wire _guard25922 = early_reset_static_par0_go_out;
wire _guard25923 = early_reset_static_par0_go_out;
wire _guard25924 = early_reset_static_par0_go_out;
wire _guard25925 = early_reset_static_par0_go_out;
wire _guard25926 = ~_guard0;
wire _guard25927 = early_reset_static_par0_go_out;
wire _guard25928 = _guard25926 & _guard25927;
wire _guard25929 = early_reset_static_par0_go_out;
wire _guard25930 = early_reset_static_par0_go_out;
wire _guard25931 = early_reset_static_par0_go_out;
wire _guard25932 = ~_guard0;
wire _guard25933 = early_reset_static_par0_go_out;
wire _guard25934 = _guard25932 & _guard25933;
wire _guard25935 = ~_guard0;
wire _guard25936 = early_reset_static_par0_go_out;
wire _guard25937 = _guard25935 & _guard25936;
wire _guard25938 = early_reset_static_par0_go_out;
wire _guard25939 = ~_guard0;
wire _guard25940 = early_reset_static_par0_go_out;
wire _guard25941 = _guard25939 & _guard25940;
wire _guard25942 = early_reset_static_par0_go_out;
wire _guard25943 = ~_guard0;
wire _guard25944 = early_reset_static_par0_go_out;
wire _guard25945 = _guard25943 & _guard25944;
wire _guard25946 = early_reset_static_par0_go_out;
wire _guard25947 = ~_guard0;
wire _guard25948 = early_reset_static_par0_go_out;
wire _guard25949 = _guard25947 & _guard25948;
wire _guard25950 = early_reset_static_par0_go_out;
wire _guard25951 = ~_guard0;
wire _guard25952 = early_reset_static_par0_go_out;
wire _guard25953 = _guard25951 & _guard25952;
wire _guard25954 = early_reset_static_par0_go_out;
wire _guard25955 = early_reset_static_par0_go_out;
wire _guard25956 = early_reset_static_par0_go_out;
wire _guard25957 = early_reset_static_par0_go_out;
wire _guard25958 = ~_guard0;
wire _guard25959 = early_reset_static_par0_go_out;
wire _guard25960 = _guard25958 & _guard25959;
wire _guard25961 = early_reset_static_par0_go_out;
wire _guard25962 = early_reset_static_par0_go_out;
wire _guard25963 = early_reset_static_par0_go_out;
wire _guard25964 = ~_guard0;
wire _guard25965 = early_reset_static_par0_go_out;
wire _guard25966 = _guard25964 & _guard25965;
wire _guard25967 = early_reset_static_par0_go_out;
wire _guard25968 = ~_guard0;
wire _guard25969 = early_reset_static_par0_go_out;
wire _guard25970 = _guard25968 & _guard25969;
wire _guard25971 = early_reset_static_par0_go_out;
wire _guard25972 = ~_guard0;
wire _guard25973 = early_reset_static_par0_go_out;
wire _guard25974 = _guard25972 & _guard25973;
wire _guard25975 = ~_guard0;
wire _guard25976 = early_reset_static_par0_go_out;
wire _guard25977 = _guard25975 & _guard25976;
wire _guard25978 = early_reset_static_par0_go_out;
wire _guard25979 = early_reset_static_par0_go_out;
wire _guard25980 = early_reset_static_par0_go_out;
wire _guard25981 = early_reset_static_par0_go_out;
wire _guard25982 = ~_guard0;
wire _guard25983 = early_reset_static_par0_go_out;
wire _guard25984 = _guard25982 & _guard25983;
wire _guard25985 = early_reset_static_par0_go_out;
wire _guard25986 = early_reset_static_par0_go_out;
wire _guard25987 = early_reset_static_par0_go_out;
wire _guard25988 = early_reset_static_par0_go_out;
wire _guard25989 = ~_guard0;
wire _guard25990 = early_reset_static_par0_go_out;
wire _guard25991 = _guard25989 & _guard25990;
wire _guard25992 = early_reset_static_par0_go_out;
wire _guard25993 = early_reset_static_par0_go_out;
wire _guard25994 = ~_guard0;
wire _guard25995 = early_reset_static_par0_go_out;
wire _guard25996 = _guard25994 & _guard25995;
wire _guard25997 = ~_guard0;
wire _guard25998 = early_reset_static_par0_go_out;
wire _guard25999 = _guard25997 & _guard25998;
wire _guard26000 = early_reset_static_par0_go_out;
wire _guard26001 = early_reset_static_par0_go_out;
wire _guard26002 = early_reset_static_par0_go_out;
wire _guard26003 = early_reset_static_par0_go_out;
wire _guard26004 = early_reset_static_par0_go_out;
wire _guard26005 = early_reset_static_par0_go_out;
wire _guard26006 = early_reset_static_par0_go_out;
wire _guard26007 = ~_guard0;
wire _guard26008 = early_reset_static_par0_go_out;
wire _guard26009 = _guard26007 & _guard26008;
wire _guard26010 = early_reset_static_par0_go_out;
wire _guard26011 = early_reset_static_par0_go_out;
wire _guard26012 = early_reset_static_par0_go_out;
wire _guard26013 = ~_guard0;
wire _guard26014 = early_reset_static_par0_go_out;
wire _guard26015 = _guard26013 & _guard26014;
wire _guard26016 = early_reset_static_par0_go_out;
wire _guard26017 = ~_guard0;
wire _guard26018 = early_reset_static_par0_go_out;
wire _guard26019 = _guard26017 & _guard26018;
wire _guard26020 = early_reset_static_par0_go_out;
wire _guard26021 = ~_guard0;
wire _guard26022 = early_reset_static_par0_go_out;
wire _guard26023 = _guard26021 & _guard26022;
wire _guard26024 = early_reset_static_par0_go_out;
wire _guard26025 = early_reset_static_par0_go_out;
wire _guard26026 = early_reset_static_par0_go_out;
wire _guard26027 = early_reset_static_par0_go_out;
wire _guard26028 = early_reset_static_par0_go_out;
wire _guard26029 = early_reset_static_par0_go_out;
wire _guard26030 = early_reset_static_par0_go_out;
wire _guard26031 = early_reset_static_par0_go_out;
wire _guard26032 = early_reset_static_par0_go_out;
wire _guard26033 = early_reset_static_par0_go_out;
wire _guard26034 = early_reset_static_par0_go_out;
wire _guard26035 = early_reset_static_par0_go_out;
wire _guard26036 = ~_guard0;
wire _guard26037 = early_reset_static_par0_go_out;
wire _guard26038 = _guard26036 & _guard26037;
wire _guard26039 = early_reset_static_par0_go_out;
wire _guard26040 = early_reset_static_par0_go_out;
assign pe_1_4_mul_ready =
  _guard3 ? 1'd1 :
  _guard6 ? 1'd0 :
  1'd0;
assign pe_1_4_clk = clk;
assign pe_1_4_top =
  _guard19 ? top_1_4_out :
  32'd0;
assign pe_1_4_left =
  _guard32 ? left_1_4_out :
  32'd0;
assign pe_1_4_reset = reset;
assign pe_1_4_go = _guard45;
assign pe_1_7_mul_ready =
  _guard48 ? 1'd1 :
  _guard51 ? 1'd0 :
  1'd0;
assign pe_1_7_clk = clk;
assign pe_1_7_top =
  _guard64 ? top_1_7_out :
  32'd0;
assign pe_1_7_left =
  _guard77 ? left_1_7_out :
  32'd0;
assign pe_1_7_reset = reset;
assign pe_1_7_go = _guard90;
assign left_1_13_write_en = _guard93;
assign left_1_13_clk = clk;
assign left_1_13_reset = reset;
assign left_1_13_in = left_1_12_out;
assign top_2_4_write_en = _guard99;
assign top_2_4_clk = clk;
assign top_2_4_reset = reset;
assign top_2_4_in = top_1_4_out;
assign left_2_4_write_en = _guard105;
assign left_2_4_clk = clk;
assign left_2_4_reset = reset;
assign left_2_4_in = left_2_3_out;
assign pe_2_12_mul_ready =
  _guard111 ? 1'd1 :
  _guard114 ? 1'd0 :
  1'd0;
assign pe_2_12_clk = clk;
assign pe_2_12_top =
  _guard127 ? top_2_12_out :
  32'd0;
assign pe_2_12_left =
  _guard140 ? left_2_12_out :
  32'd0;
assign pe_2_12_reset = reset;
assign pe_2_12_go = _guard153;
assign top_3_5_write_en = _guard156;
assign top_3_5_clk = clk;
assign top_3_5_reset = reset;
assign top_3_5_in = top_2_5_out;
assign top_3_6_write_en = _guard162;
assign top_3_6_clk = clk;
assign top_3_6_reset = reset;
assign top_3_6_in = top_2_6_out;
assign pe_3_8_mul_ready =
  _guard168 ? 1'd1 :
  _guard171 ? 1'd0 :
  1'd0;
assign pe_3_8_clk = clk;
assign pe_3_8_top =
  _guard184 ? top_3_8_out :
  32'd0;
assign pe_3_8_left =
  _guard197 ? left_3_8_out :
  32'd0;
assign pe_3_8_reset = reset;
assign pe_3_8_go = _guard210;
assign left_4_0_write_en = _guard213;
assign left_4_0_clk = clk;
assign left_4_0_reset = reset;
assign left_4_0_in = l4_read_data;
assign top_4_4_write_en = _guard219;
assign top_4_4_clk = clk;
assign top_4_4_reset = reset;
assign top_4_4_in = top_3_4_out;
assign pe_4_9_mul_ready =
  _guard225 ? 1'd1 :
  _guard228 ? 1'd0 :
  1'd0;
assign pe_4_9_clk = clk;
assign pe_4_9_top =
  _guard241 ? top_4_9_out :
  32'd0;
assign pe_4_9_left =
  _guard254 ? left_4_9_out :
  32'd0;
assign pe_4_9_reset = reset;
assign pe_4_9_go = _guard267;
assign pe_5_2_mul_ready =
  _guard270 ? 1'd1 :
  _guard273 ? 1'd0 :
  1'd0;
assign pe_5_2_clk = clk;
assign pe_5_2_top =
  _guard286 ? top_5_2_out :
  32'd0;
assign pe_5_2_left =
  _guard299 ? left_5_2_out :
  32'd0;
assign pe_5_2_reset = reset;
assign pe_5_2_go = _guard312;
assign top_5_8_write_en = _guard315;
assign top_5_8_clk = clk;
assign top_5_8_reset = reset;
assign top_5_8_in = top_4_8_out;
assign top_6_1_write_en = _guard321;
assign top_6_1_clk = clk;
assign top_6_1_reset = reset;
assign top_6_1_in = top_5_1_out;
assign left_6_2_write_en = _guard327;
assign left_6_2_clk = clk;
assign left_6_2_reset = reset;
assign left_6_2_in = left_6_1_out;
assign top_6_3_write_en = _guard333;
assign top_6_3_clk = clk;
assign top_6_3_reset = reset;
assign top_6_3_in = top_5_3_out;
assign left_6_4_write_en = _guard339;
assign left_6_4_clk = clk;
assign left_6_4_reset = reset;
assign left_6_4_in = left_6_3_out;
assign top_6_13_write_en = _guard345;
assign top_6_13_clk = clk;
assign top_6_13_reset = reset;
assign top_6_13_in = top_5_13_out;
assign top_7_0_write_en = _guard351;
assign top_7_0_clk = clk;
assign top_7_0_reset = reset;
assign top_7_0_in = top_6_0_out;
assign pe_7_9_mul_ready =
  _guard357 ? 1'd1 :
  _guard360 ? 1'd0 :
  1'd0;
assign pe_7_9_clk = clk;
assign pe_7_9_top =
  _guard373 ? top_7_9_out :
  32'd0;
assign pe_7_9_left =
  _guard386 ? left_7_9_out :
  32'd0;
assign pe_7_9_reset = reset;
assign pe_7_9_go = _guard399;
assign left_7_14_write_en = _guard402;
assign left_7_14_clk = clk;
assign left_7_14_reset = reset;
assign left_7_14_in = left_7_13_out;
assign top_8_4_write_en = _guard408;
assign top_8_4_clk = clk;
assign top_8_4_reset = reset;
assign top_8_4_in = top_7_4_out;
assign left_8_11_write_en = _guard414;
assign left_8_11_clk = clk;
assign left_8_11_reset = reset;
assign left_8_11_in = left_8_10_out;
assign left_9_5_write_en = _guard420;
assign left_9_5_clk = clk;
assign left_9_5_reset = reset;
assign left_9_5_in = left_9_4_out;
assign pe_9_15_mul_ready =
  _guard426 ? 1'd1 :
  _guard429 ? 1'd0 :
  1'd0;
assign pe_9_15_clk = clk;
assign pe_9_15_top =
  _guard442 ? top_9_15_out :
  32'd0;
assign pe_9_15_left =
  _guard455 ? left_9_15_out :
  32'd0;
assign pe_9_15_reset = reset;
assign pe_9_15_go = _guard468;
assign pe_10_5_mul_ready =
  _guard471 ? 1'd1 :
  _guard474 ? 1'd0 :
  1'd0;
assign pe_10_5_clk = clk;
assign pe_10_5_top =
  _guard487 ? top_10_5_out :
  32'd0;
assign pe_10_5_left =
  _guard500 ? left_10_5_out :
  32'd0;
assign pe_10_5_reset = reset;
assign pe_10_5_go = _guard513;
assign top_10_8_write_en = _guard516;
assign top_10_8_clk = clk;
assign top_10_8_reset = reset;
assign top_10_8_in = top_9_8_out;
assign top_10_13_write_en = _guard522;
assign top_10_13_clk = clk;
assign top_10_13_reset = reset;
assign top_10_13_in = top_9_13_out;
assign top_11_15_write_en = _guard528;
assign top_11_15_clk = clk;
assign top_11_15_reset = reset;
assign top_11_15_in = top_10_15_out;
assign top_12_3_write_en = _guard534;
assign top_12_3_clk = clk;
assign top_12_3_reset = reset;
assign top_12_3_in = top_11_3_out;
assign left_12_4_write_en = _guard540;
assign left_12_4_clk = clk;
assign left_12_4_reset = reset;
assign left_12_4_in = left_12_3_out;
assign pe_12_10_mul_ready =
  _guard546 ? 1'd1 :
  _guard549 ? 1'd0 :
  1'd0;
assign pe_12_10_clk = clk;
assign pe_12_10_top =
  _guard562 ? top_12_10_out :
  32'd0;
assign pe_12_10_left =
  _guard575 ? left_12_10_out :
  32'd0;
assign pe_12_10_reset = reset;
assign pe_12_10_go = _guard588;
assign left_13_2_write_en = _guard591;
assign left_13_2_clk = clk;
assign left_13_2_reset = reset;
assign left_13_2_in = left_13_1_out;
assign top_13_7_write_en = _guard597;
assign top_13_7_clk = clk;
assign top_13_7_reset = reset;
assign top_13_7_in = top_12_7_out;
assign top_13_12_write_en = _guard603;
assign top_13_12_clk = clk;
assign top_13_12_reset = reset;
assign top_13_12_in = top_12_12_out;
assign pe_13_14_mul_ready =
  _guard609 ? 1'd1 :
  _guard612 ? 1'd0 :
  1'd0;
assign pe_13_14_clk = clk;
assign pe_13_14_top =
  _guard625 ? top_13_14_out :
  32'd0;
assign pe_13_14_left =
  _guard638 ? left_13_14_out :
  32'd0;
assign pe_13_14_reset = reset;
assign pe_13_14_go = _guard651;
assign top_14_0_write_en = _guard654;
assign top_14_0_clk = clk;
assign top_14_0_reset = reset;
assign top_14_0_in = top_13_0_out;
assign top_14_15_write_en = _guard660;
assign top_14_15_clk = clk;
assign top_14_15_reset = reset;
assign top_14_15_in = top_13_15_out;
assign top_15_0_write_en = _guard666;
assign top_15_0_clk = clk;
assign top_15_0_reset = reset;
assign top_15_0_in = top_14_0_out;
assign top_15_7_write_en = _guard672;
assign top_15_7_clk = clk;
assign top_15_7_reset = reset;
assign top_15_7_in = top_14_7_out;
assign t3_add_left = 5'd1;
assign t3_add_right = t3_idx_out;
assign t15_idx_write_en = _guard688;
assign t15_idx_clk = clk;
assign t15_idx_reset = reset;
assign t15_idx_in =
  _guard691 ? 5'd0 :
  _guard694 ? t15_add_out :
  'x;
assign l1_add_left = 5'd1;
assign l1_add_right = l1_idx_out;
assign l12_idx_write_en = _guard707;
assign l12_idx_clk = clk;
assign l12_idx_reset = reset;
assign l12_idx_in =
  _guard710 ? 5'd0 :
  _guard713 ? l12_add_out :
  'x;
assign l13_idx_write_en = _guard720;
assign l13_idx_clk = clk;
assign l13_idx_reset = reset;
assign l13_idx_in =
  _guard723 ? 5'd0 :
  _guard726 ? l13_add_out :
  'x;
assign index_ge_30_left = idx_add_out;
assign index_ge_30_right = 6'd30;
assign idx_between_35_51_comb_left = index_ge_35_out;
assign idx_between_35_51_comb_right = index_lt_51_out;
assign idx_between_17_21_comb_left = index_ge_17_out;
assign idx_between_17_21_comb_right = index_lt_21_out;
assign idx_between_41_42_comb_left = index_ge_41_out;
assign idx_between_41_42_comb_right = index_lt_42_out;
assign idx_between_1_17_reg_write_en = _guard739;
assign idx_between_1_17_reg_clk = clk;
assign idx_between_1_17_reg_reset = reset;
assign idx_between_1_17_reg_in =
  _guard740 ? idx_between_1_17_comb_out :
  _guard743 ? 1'd0 :
  'x;
assign idx_between_42_43_reg_write_en = _guard748;
assign idx_between_42_43_reg_clk = clk;
assign idx_between_42_43_reg_reset = reset;
assign idx_between_42_43_reg_in =
  _guard751 ? 1'd0 :
  _guard752 ? idx_between_42_43_comb_out :
  'x;
assign idx_between_29_45_comb_left = index_ge_29_out;
assign idx_between_29_45_comb_right = index_lt_45_out;
assign idx_between_30_34_comb_left = index_ge_30_out;
assign idx_between_30_34_comb_right = index_lt_34_out;
assign idx_between_7_23_reg_write_en = _guard761;
assign idx_between_7_23_reg_clk = clk;
assign idx_between_7_23_reg_reset = reset;
assign idx_between_7_23_reg_in =
  _guard762 ? idx_between_7_23_comb_out :
  _guard765 ? 1'd0 :
  'x;
assign idx_between_21_25_comb_left = index_ge_21_out;
assign idx_between_21_25_comb_right = index_lt_25_out;
assign idx_between_45_46_comb_left = index_ge_45_out;
assign idx_between_45_46_comb_right = index_lt_46_out;
assign idx_between_32_48_comb_left = index_ge_32_out;
assign idx_between_32_48_comb_right = index_lt_48_out;
assign index_lt_5_left = idx_add_out;
assign index_lt_5_right = 6'd5;
assign idx_between_24_25_comb_left = index_ge_24_out;
assign idx_between_24_25_comb_right = index_lt_25_out;
assign idx_between_11_27_reg_write_en = _guard780;
assign idx_between_11_27_reg_clk = clk;
assign idx_between_11_27_reg_reset = reset;
assign idx_between_11_27_reg_in =
  _guard781 ? idx_between_11_27_comb_out :
  _guard784 ? 1'd0 :
  'x;
assign idx_between_3_7_reg_write_en = _guard789;
assign idx_between_3_7_reg_clk = clk;
assign idx_between_3_7_reg_reset = reset;
assign idx_between_3_7_reg_in =
  _guard790 ? idx_between_3_7_comb_out :
  _guard793 ? 1'd0 :
  'x;
assign index_ge_15_left = idx_add_out;
assign index_ge_15_right = 6'd15;
assign idx_between_19_23_reg_write_en = _guard800;
assign idx_between_19_23_reg_clk = clk;
assign idx_between_19_23_reg_reset = reset;
assign idx_between_19_23_reg_in =
  _guard801 ? idx_between_19_23_comb_out :
  _guard804 ? 1'd0 :
  'x;
assign idx_between_15_19_reg_write_en = _guard809;
assign idx_between_15_19_reg_clk = clk;
assign idx_between_15_19_reg_reset = reset;
assign idx_between_15_19_reg_in =
  _guard810 ? idx_between_15_19_comb_out :
  _guard813 ? 1'd0 :
  'x;
assign idx_between_34_35_reg_write_en = _guard818;
assign idx_between_34_35_reg_clk = clk;
assign idx_between_34_35_reg_reset = reset;
assign idx_between_34_35_reg_in =
  _guard819 ? idx_between_34_35_comb_out :
  _guard822 ? 1'd0 :
  'x;
assign cond_wire3_in =
  _guard823 ? idx_between_21_22_reg_out :
  _guard826 ? cond3_out :
  1'd0;
assign cond_wire30_in =
  _guard829 ? cond30_out :
  _guard830 ? idx_between_7_11_reg_out :
  1'd0;
assign cond_wire38_in =
  _guard831 ? idx_between_28_29_reg_out :
  _guard834 ? cond38_out :
  1'd0;
assign cond_wire39_in =
  _guard835 ? idx_between_8_24_reg_out :
  _guard838 ? cond39_out :
  1'd0;
assign cond_wire47_in =
  _guard839 ? idx_between_14_30_reg_out :
  _guard842 ? cond47_out :
  1'd0;
assign cond53_write_en = _guard843;
assign cond53_clk = clk;
assign cond53_reset = reset;
assign cond53_in =
  _guard844 ? idx_between_31_32_reg_out :
  1'd0;
assign cond_wire54_in =
  _guard845 ? idx_between_11_27_reg_out :
  _guard848 ? cond54_out :
  1'd0;
assign cond65_write_en = _guard849;
assign cond65_clk = clk;
assign cond65_reset = reset;
assign cond65_in =
  _guard850 ? idx_between_14_18_reg_out :
  1'd0;
assign cond70_write_en = _guard851;
assign cond70_clk = clk;
assign cond70_reset = reset;
assign cond70_in =
  _guard852 ? idx_between_15_19_reg_out :
  1'd0;
assign cond71_write_en = _guard853;
assign cond71_clk = clk;
assign cond71_reset = reset;
assign cond71_in =
  _guard854 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire89_in =
  _guard857 ? cond89_out :
  _guard858 ? idx_between_4_20_reg_out :
  1'd0;
assign cond_wire90_in =
  _guard861 ? cond90_out :
  _guard862 ? idx_between_8_24_reg_out :
  1'd0;
assign cond_wire103_in =
  _guard865 ? cond103_out :
  _guard866 ? idx_between_27_28_reg_out :
  1'd0;
assign cond_wire131_in =
  _guard867 ? idx_between_34_35_reg_out :
  _guard870 ? cond131_out :
  1'd0;
assign cond_wire164_in =
  _guard873 ? cond164_out :
  _guard874 ? idx_between_27_28_reg_out :
  1'd0;
assign cond167_write_en = _guard875;
assign cond167_clk = clk;
assign cond167_reset = reset;
assign cond167_in =
  _guard876 ? idx_between_12_28_reg_out :
  1'd0;
assign cond181_write_en = _guard877;
assign cond181_clk = clk;
assign cond181_reset = reset;
assign cond181_in =
  _guard878 ? idx_between_12_16_reg_out :
  1'd0;
assign cond_wire185_in =
  _guard879 ? idx_between_13_17_reg_out :
  _guard882 ? cond185_out :
  1'd0;
assign cond_wire193_in =
  _guard883 ? idx_between_15_19_reg_out :
  _guard886 ? cond193_out :
  1'd0;
assign cond202_write_en = _guard887;
assign cond202_clk = clk;
assign cond202_reset = reset;
assign cond202_in =
  _guard888 ? idx_between_17_33_reg_out :
  1'd0;
assign cond_wire204_in =
  _guard891 ? cond204_out :
  _guard892 ? idx_between_37_38_reg_out :
  1'd0;
assign cond_wire224_in =
  _guard893 ? idx_between_11_27_reg_out :
  _guard896 ? cond224_out :
  1'd0;
assign cond227_write_en = _guard897;
assign cond227_clk = clk;
assign cond227_reset = reset;
assign cond227_in =
  _guard898 ? idx_between_8_24_reg_out :
  1'd0;
assign cond230_write_en = _guard899;
assign cond230_clk = clk;
assign cond230_reset = reset;
assign cond230_in =
  _guard900 ? idx_between_9_13_reg_out :
  1'd0;
assign cond_wire234_in =
  _guard901 ? idx_between_10_14_reg_out :
  _guard904 ? cond234_out :
  1'd0;
assign cond239_write_en = _guard905;
assign cond239_clk = clk;
assign cond239_reset = reset;
assign cond239_in =
  _guard906 ? idx_between_11_27_reg_out :
  1'd0;
assign cond_wire240_in =
  _guard909 ? cond240_out :
  _guard910 ? idx_between_15_31_reg_out :
  1'd0;
assign cond263_write_en = _guard911;
assign cond263_clk = clk;
assign cond263_reset = reset;
assign cond263_in =
  _guard912 ? idx_between_17_33_reg_out :
  1'd0;
assign cond281_write_en = _guard913;
assign cond281_clk = clk;
assign cond281_reset = reset;
assign cond281_in =
  _guard914 ? idx_between_10_26_reg_out :
  1'd0;
assign cond287_write_en = _guard915;
assign cond287_clk = clk;
assign cond287_reset = reset;
assign cond287_in =
  _guard916 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire291_in =
  _guard919 ? cond291_out :
  _guard920 ? idx_between_9_13_reg_out :
  1'd0;
assign cond_wire302_in =
  _guard923 ? cond302_out :
  _guard924 ? idx_between_31_32_reg_out :
  1'd0;
assign cond_wire305_in =
  _guard925 ? idx_between_16_32_reg_out :
  _guard928 ? cond305_out :
  1'd0;
assign cond_wire316_in =
  _guard931 ? cond316_out :
  _guard932 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire324_in =
  _guard933 ? idx_between_17_33_reg_out :
  _guard936 ? cond324_out :
  1'd0;
assign cond_wire336_in =
  _guard937 ? idx_between_20_36_reg_out :
  _guard940 ? cond336_out :
  1'd0;
assign cond_wire338_in =
  _guard941 ? idx_between_40_41_reg_out :
  _guard944 ? cond338_out :
  1'd0;
assign cond340_write_en = _guard945;
assign cond340_clk = clk;
assign cond340_reset = reset;
assign cond340_in =
  _guard946 ? idx_between_6_10_reg_out :
  1'd0;
assign cond342_write_en = _guard947;
assign cond342_clk = clk;
assign cond342_reset = reset;
assign cond342_in =
  _guard948 ? idx_between_10_26_reg_out :
  1'd0;
assign cond350_write_en = _guard949;
assign cond350_clk = clk;
assign cond350_reset = reset;
assign cond350_in =
  _guard950 ? idx_between_12_28_reg_out :
  1'd0;
assign cond356_write_en = _guard951;
assign cond356_clk = clk;
assign cond356_reset = reset;
assign cond356_in =
  _guard952 ? idx_between_10_14_reg_out :
  1'd0;
assign cond375_write_en = _guard953;
assign cond375_clk = clk;
assign cond375_reset = reset;
assign cond375_in =
  _guard954 ? idx_between_34_35_reg_out :
  1'd0;
assign cond_wire380_in =
  _guard955 ? idx_between_16_20_reg_out :
  _guard958 ? cond380_out :
  1'd0;
assign cond_wire394_in =
  _guard959 ? idx_between_23_39_reg_out :
  _guard962 ? cond394_out :
  1'd0;
assign cond_wire399_in =
  _guard963 ? idx_between_40_41_reg_out :
  _guard966 ? cond399_out :
  1'd0;
assign cond_wire403_in =
  _guard967 ? idx_between_41_42_reg_out :
  _guard970 ? cond403_out :
  1'd0;
assign cond_wire411_in =
  _guard973 ? cond411_out :
  _guard974 ? idx_between_12_28_reg_out :
  1'd0;
assign cond420_write_en = _guard975;
assign cond420_clk = clk;
assign cond420_reset = reset;
assign cond420_in =
  _guard976 ? idx_between_30_31_reg_out :
  1'd0;
assign cond_wire422_in =
  _guard977 ? idx_between_11_27_reg_out :
  _guard980 ? cond422_out :
  1'd0;
assign cond_wire425_in =
  _guard981 ? idx_between_12_16_reg_out :
  _guard984 ? cond425_out :
  1'd0;
assign cond435_write_en = _guard985;
assign cond435_clk = clk;
assign cond435_reset = reset;
assign cond435_in =
  _guard986 ? idx_between_18_34_reg_out :
  1'd0;
assign cond_wire462_in =
  _guard989 ? cond462_out :
  _guard990 ? idx_between_21_37_reg_out :
  1'd0;
assign cond463_write_en = _guard991;
assign cond463_clk = clk;
assign cond463_reset = reset;
assign cond463_in =
  _guard992 ? idx_between_25_41_reg_out :
  1'd0;
assign cond_wire471_in =
  _guard995 ? cond471_out :
  _guard996 ? idx_between_8_24_reg_out :
  1'd0;
assign cond476_write_en = _guard997;
assign cond476_clk = clk;
assign cond476_reset = reset;
assign cond476_in =
  _guard998 ? idx_between_13_29_reg_out :
  1'd0;
assign cond495_write_en = _guard999;
assign cond495_clk = clk;
assign cond495_reset = reset;
assign cond495_in =
  _guard1000 ? idx_between_14_30_reg_out :
  1'd0;
assign cond499_write_en = _guard1001;
assign cond499_clk = clk;
assign cond499_reset = reset;
assign cond499_in =
  _guard1002 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire505_in =
  _guard1003 ? idx_between_36_37_reg_out :
  _guard1006 ? cond505_out :
  1'd0;
assign cond_wire512_in =
  _guard1007 ? idx_between_22_38_reg_out :
  _guard1010 ? cond512_out :
  1'd0;
assign cond518_write_en = _guard1011;
assign cond518_clk = clk;
assign cond518_reset = reset;
assign cond518_in =
  _guard1012 ? idx_between_20_24_reg_out :
  1'd0;
assign cond_wire520_in =
  _guard1015 ? cond520_out :
  _guard1016 ? idx_between_24_40_reg_out :
  1'd0;
assign cond_wire523_in =
  _guard1019 ? cond523_out :
  _guard1020 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire542_in =
  _guard1023 ? cond542_out :
  _guard1024 ? idx_between_30_31_reg_out :
  1'd0;
assign cond554_write_en = _guard1025;
assign cond554_clk = clk;
assign cond554_reset = reset;
assign cond554_in =
  _guard1026 ? idx_between_33_34_reg_out :
  1'd0;
assign cond_wire578_in =
  _guard1029 ? cond578_out :
  _guard1030 ? idx_between_39_40_reg_out :
  1'd0;
assign cond_wire579_in =
  _guard1031 ? idx_between_20_24_reg_out :
  _guard1034 ? cond579_out :
  1'd0;
assign cond581_write_en = _guard1035;
assign cond581_clk = clk;
assign cond581_reset = reset;
assign cond581_in =
  _guard1036 ? idx_between_24_40_reg_out :
  1'd0;
assign cond_wire581_in =
  _guard1039 ? cond581_out :
  _guard1040 ? idx_between_24_40_reg_out :
  1'd0;
assign cond_wire582_in =
  _guard1043 ? cond582_out :
  _guard1044 ? idx_between_40_41_reg_out :
  1'd0;
assign cond_wire589_in =
  _guard1047 ? cond589_out :
  _guard1048 ? idx_between_26_42_reg_out :
  1'd0;
assign cond_wire591_in =
  _guard1049 ? idx_between_23_27_reg_out :
  _guard1052 ? cond591_out :
  1'd0;
assign cond_wire630_in =
  _guard1053 ? idx_between_21_37_reg_out :
  _guard1056 ? cond630_out :
  1'd0;
assign cond667_write_en = _guard1057;
assign cond667_clk = clk;
assign cond667_reset = reset;
assign cond667_in =
  _guard1058 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire680_in =
  _guard1059 ? idx_between_34_35_reg_out :
  _guard1062 ? cond680_out :
  1'd0;
assign cond708_write_en = _guard1063;
assign cond708_clk = clk;
assign cond708_reset = reset;
assign cond708_in =
  _guard1064 ? idx_between_41_42_reg_out :
  1'd0;
assign cond743_write_en = _guard1065;
assign cond743_clk = clk;
assign cond743_reset = reset;
assign cond743_in =
  _guard1066 ? idx_between_15_31_reg_out :
  1'd0;
assign cond760_write_en = _guard1067;
assign cond760_clk = clk;
assign cond760_reset = reset;
assign cond760_in =
  _guard1068 ? idx_between_23_39_reg_out :
  1'd0;
assign cond763_write_en = _guard1069;
assign cond763_clk = clk;
assign cond763_reset = reset;
assign cond763_in =
  _guard1070 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire765_in =
  _guard1073 ? cond765_out :
  _guard1074 ? idx_between_40_41_reg_out :
  1'd0;
assign cond767_write_en = _guard1075;
assign cond767_clk = clk;
assign cond767_reset = reset;
assign cond767_in =
  _guard1076 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire768_in =
  _guard1079 ? cond768_out :
  _guard1080 ? idx_between_25_41_reg_out :
  1'd0;
assign cond792_write_en = _guard1081;
assign cond792_clk = clk;
assign cond792_reset = reset;
assign cond792_in =
  _guard1082 ? idx_between_31_47_reg_out :
  1'd0;
assign cond_wire794_in =
  _guard1085 ? cond794_out :
  _guard1086 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire799_in =
  _guard1089 ? cond799_out :
  _guard1090 ? idx_between_14_18_reg_out :
  1'd0;
assign cond_wire803_in =
  _guard1091 ? idx_between_15_19_reg_out :
  _guard1094 ? cond803_out :
  1'd0;
assign cond804_write_en = _guard1095;
assign cond804_clk = clk;
assign cond804_reset = reset;
assign cond804_in =
  _guard1096 ? idx_between_15_31_reg_out :
  1'd0;
assign cond822_write_en = _guard1097;
assign cond822_clk = clk;
assign cond822_reset = reset;
assign cond822_in =
  _guard1098 ? idx_between_39_40_reg_out :
  1'd0;
assign cond829_write_en = _guard1099;
assign cond829_clk = clk;
assign cond829_reset = reset;
assign cond829_in =
  _guard1100 ? idx_between_25_41_reg_out :
  1'd0;
assign cond_wire854_in =
  _guard1101 ? idx_between_47_48_reg_out :
  _guard1104 ? cond854_out :
  1'd0;
assign cond_wire857_in =
  _guard1105 ? idx_between_32_48_reg_out :
  _guard1108 ? cond857_out :
  1'd0;
assign cond861_write_en = _guard1109;
assign cond861_clk = clk;
assign cond861_reset = reset;
assign cond861_in =
  _guard1110 ? idx_between_14_30_reg_out :
  1'd0;
assign cond_wire863_in =
  _guard1111 ? idx_between_34_35_reg_out :
  _guard1114 ? cond863_out :
  1'd0;
assign cond_wire881_in =
  _guard1115 ? idx_between_19_35_reg_out :
  _guard1118 ? cond881_out :
  1'd0;
assign cond_wire886_in =
  _guard1119 ? idx_between_24_40_reg_out :
  _guard1122 ? cond886_out :
  1'd0;
assign cond899_write_en = _guard1123;
assign cond899_clk = clk;
assign cond899_reset = reset;
assign cond899_in =
  _guard1124 ? idx_between_43_44_reg_out :
  1'd0;
assign cond_wire905_in =
  _guard1125 ? idx_between_25_41_reg_out :
  _guard1128 ? cond905_out :
  1'd0;
assign cond_wire908_in =
  _guard1131 ? cond908_out :
  _guard1132 ? idx_between_26_30_reg_out :
  1'd0;
assign cond_wire927_in =
  _guard1135 ? cond927_out :
  _guard1136 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire928_in =
  _guard1137 ? idx_between_35_36_reg_out :
  _guard1140 ? cond928_out :
  1'd0;
assign cond_wire932_in =
  _guard1143 ? cond932_out :
  _guard1144 ? idx_between_36_37_reg_out :
  1'd0;
assign cond_wire939_in =
  _guard1147 ? cond939_out :
  _guard1148 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire941_in =
  _guard1149 ? idx_between_19_23_reg_out :
  _guard1152 ? cond941_out :
  1'd0;
assign cond944_write_en = _guard1153;
assign cond944_clk = clk;
assign cond944_reset = reset;
assign cond944_in =
  _guard1154 ? idx_between_39_40_reg_out :
  1'd0;
assign cond_wire949_in =
  _guard1157 ? cond949_out :
  _guard1158 ? idx_between_21_25_reg_out :
  1'd0;
assign cond955_write_en = _guard1159;
assign cond955_clk = clk;
assign cond955_reset = reset;
assign cond955_in =
  _guard1160 ? idx_between_26_42_reg_out :
  1'd0;
assign cond957_write_en = _guard1161;
assign cond957_clk = clk;
assign cond957_reset = reset;
assign cond957_in =
  _guard1162 ? idx_between_23_27_reg_out :
  1'd0;
assign cond977_write_en = _guard1163;
assign cond977_clk = clk;
assign cond977_reset = reset;
assign cond977_in =
  _guard1164 ? idx_between_28_32_reg_out :
  1'd0;
assign cond987_write_en = _guard1165;
assign cond987_clk = clk;
assign cond987_reset = reset;
assign cond987_in =
  _guard1166 ? idx_between_34_50_reg_out :
  1'd0;
assign cond996_write_en = _guard1167;
assign cond996_clk = clk;
assign cond996_reset = reset;
assign cond996_in =
  _guard1168 ? idx_between_21_37_reg_out :
  1'd0;
assign cond1005_write_en = _guard1169;
assign cond1005_clk = clk;
assign cond1005_reset = reset;
assign cond1005_in =
  _guard1170 ? idx_between_39_40_reg_out :
  1'd0;
assign cond_wire1011_in =
  _guard1171 ? idx_between_21_37_reg_out :
  _guard1174 ? cond1011_out :
  1'd0;
assign cond_wire1026_in =
  _guard1175 ? idx_between_25_29_reg_out :
  _guard1178 ? cond1026_out :
  1'd0;
assign cond_wire1030_in =
  _guard1179 ? idx_between_26_30_reg_out :
  _guard1182 ? cond1030_out :
  1'd0;
assign cond_wire1036_in =
  _guard1183 ? idx_between_31_47_reg_out :
  _guard1186 ? cond1036_out :
  1'd0;
assign cond_wire1040_in =
  _guard1187 ? idx_between_32_48_reg_out :
  _guard1190 ? cond1040_out :
  1'd0;
assign cond_wire1046_in =
  _guard1191 ? idx_between_30_34_reg_out :
  _guard1194 ? cond1046_out :
  1'd0;
assign cond_wire1047_in =
  _guard1195 ? idx_between_30_46_reg_out :
  _guard1198 ? cond1047_out :
  1'd0;
assign left_0_3_write_en = _guard1201;
assign left_0_3_clk = clk;
assign left_0_3_reset = reset;
assign left_0_3_in = left_0_2_out;
assign left_0_4_write_en = _guard1207;
assign left_0_4_clk = clk;
assign left_0_4_reset = reset;
assign left_0_4_in = left_0_3_out;
assign pe_0_10_mul_ready =
  _guard1213 ? 1'd1 :
  _guard1216 ? 1'd0 :
  1'd0;
assign pe_0_10_clk = clk;
assign pe_0_10_top =
  _guard1229 ? top_0_10_out :
  32'd0;
assign pe_0_10_left =
  _guard1242 ? left_0_10_out :
  32'd0;
assign pe_0_10_reset = reset;
assign pe_0_10_go = _guard1255;
assign top_1_0_write_en = _guard1258;
assign top_1_0_clk = clk;
assign top_1_0_reset = reset;
assign top_1_0_in = top_0_0_out;
assign pe_1_2_mul_ready =
  _guard1264 ? 1'd1 :
  _guard1267 ? 1'd0 :
  1'd0;
assign pe_1_2_clk = clk;
assign pe_1_2_top =
  _guard1280 ? top_1_2_out :
  32'd0;
assign pe_1_2_left =
  _guard1293 ? left_1_2_out :
  32'd0;
assign pe_1_2_reset = reset;
assign pe_1_2_go = _guard1306;
assign pe_1_3_mul_ready =
  _guard1309 ? 1'd1 :
  _guard1312 ? 1'd0 :
  1'd0;
assign pe_1_3_clk = clk;
assign pe_1_3_top =
  _guard1325 ? top_1_3_out :
  32'd0;
assign pe_1_3_left =
  _guard1338 ? left_1_3_out :
  32'd0;
assign pe_1_3_reset = reset;
assign pe_1_3_go = _guard1351;
assign left_1_3_write_en = _guard1354;
assign left_1_3_clk = clk;
assign left_1_3_reset = reset;
assign left_1_3_in = left_1_2_out;
assign top_1_13_write_en = _guard1360;
assign top_1_13_clk = clk;
assign top_1_13_reset = reset;
assign top_1_13_in = top_0_13_out;
assign left_1_14_write_en = _guard1366;
assign left_1_14_clk = clk;
assign left_1_14_reset = reset;
assign left_1_14_in = left_1_13_out;
assign left_2_6_write_en = _guard1372;
assign left_2_6_clk = clk;
assign left_2_6_reset = reset;
assign left_2_6_in = left_2_5_out;
assign left_2_8_write_en = _guard1378;
assign left_2_8_clk = clk;
assign left_2_8_reset = reset;
assign left_2_8_in = left_2_7_out;
assign pe_2_11_mul_ready =
  _guard1384 ? 1'd1 :
  _guard1387 ? 1'd0 :
  1'd0;
assign pe_2_11_clk = clk;
assign pe_2_11_top =
  _guard1400 ? top_2_11_out :
  32'd0;
assign pe_2_11_left =
  _guard1413 ? left_2_11_out :
  32'd0;
assign pe_2_11_reset = reset;
assign pe_2_11_go = _guard1426;
assign top_4_7_write_en = _guard1429;
assign top_4_7_clk = clk;
assign top_4_7_reset = reset;
assign top_4_7_in = top_3_7_out;
assign left_5_1_write_en = _guard1435;
assign left_5_1_clk = clk;
assign left_5_1_reset = reset;
assign left_5_1_in = left_5_0_out;
assign left_5_3_write_en = _guard1441;
assign left_5_3_clk = clk;
assign left_5_3_reset = reset;
assign left_5_3_in = left_5_2_out;
assign pe_5_8_mul_ready =
  _guard1447 ? 1'd1 :
  _guard1450 ? 1'd0 :
  1'd0;
assign pe_5_8_clk = clk;
assign pe_5_8_top =
  _guard1463 ? top_5_8_out :
  32'd0;
assign pe_5_8_left =
  _guard1476 ? left_5_8_out :
  32'd0;
assign pe_5_8_reset = reset;
assign pe_5_8_go = _guard1489;
assign pe_5_13_mul_ready =
  _guard1492 ? 1'd1 :
  _guard1495 ? 1'd0 :
  1'd0;
assign pe_5_13_clk = clk;
assign pe_5_13_top =
  _guard1508 ? top_5_13_out :
  32'd0;
assign pe_5_13_left =
  _guard1521 ? left_5_13_out :
  32'd0;
assign pe_5_13_reset = reset;
assign pe_5_13_go = _guard1534;
assign top_5_14_write_en = _guard1537;
assign top_5_14_clk = clk;
assign top_5_14_reset = reset;
assign top_5_14_in = top_4_14_out;
assign pe_6_4_mul_ready =
  _guard1543 ? 1'd1 :
  _guard1546 ? 1'd0 :
  1'd0;
assign pe_6_4_clk = clk;
assign pe_6_4_top =
  _guard1559 ? top_6_4_out :
  32'd0;
assign pe_6_4_left =
  _guard1572 ? left_6_4_out :
  32'd0;
assign pe_6_4_reset = reset;
assign pe_6_4_go = _guard1585;
assign top_6_7_write_en = _guard1588;
assign top_6_7_clk = clk;
assign top_6_7_reset = reset;
assign top_6_7_in = top_5_7_out;
assign left_6_12_write_en = _guard1594;
assign left_6_12_clk = clk;
assign left_6_12_reset = reset;
assign left_6_12_in = left_6_11_out;
assign pe_7_3_mul_ready =
  _guard1600 ? 1'd1 :
  _guard1603 ? 1'd0 :
  1'd0;
assign pe_7_3_clk = clk;
assign pe_7_3_top =
  _guard1616 ? top_7_3_out :
  32'd0;
assign pe_7_3_left =
  _guard1629 ? left_7_3_out :
  32'd0;
assign pe_7_3_reset = reset;
assign pe_7_3_go = _guard1642;
assign left_7_4_write_en = _guard1645;
assign left_7_4_clk = clk;
assign left_7_4_reset = reset;
assign left_7_4_in = left_7_3_out;
assign left_7_6_write_en = _guard1651;
assign left_7_6_clk = clk;
assign left_7_6_reset = reset;
assign left_7_6_in = left_7_5_out;
assign top_7_7_write_en = _guard1657;
assign top_7_7_clk = clk;
assign top_7_7_reset = reset;
assign top_7_7_in = top_6_7_out;
assign left_7_9_write_en = _guard1663;
assign left_7_9_clk = clk;
assign left_7_9_reset = reset;
assign left_7_9_in = left_7_8_out;
assign top_8_2_write_en = _guard1669;
assign top_8_2_clk = clk;
assign top_8_2_reset = reset;
assign top_8_2_in = top_7_2_out;
assign pe_8_6_mul_ready =
  _guard1675 ? 1'd1 :
  _guard1678 ? 1'd0 :
  1'd0;
assign pe_8_6_clk = clk;
assign pe_8_6_top =
  _guard1691 ? top_8_6_out :
  32'd0;
assign pe_8_6_left =
  _guard1704 ? left_8_6_out :
  32'd0;
assign pe_8_6_reset = reset;
assign pe_8_6_go = _guard1717;
assign top_8_6_write_en = _guard1720;
assign top_8_6_clk = clk;
assign top_8_6_reset = reset;
assign top_8_6_in = top_7_6_out;
assign top_8_10_write_en = _guard1726;
assign top_8_10_clk = clk;
assign top_8_10_reset = reset;
assign top_8_10_in = top_7_10_out;
assign left_8_14_write_en = _guard1732;
assign left_8_14_clk = clk;
assign left_8_14_reset = reset;
assign left_8_14_in = left_8_13_out;
assign left_8_15_write_en = _guard1738;
assign left_8_15_clk = clk;
assign left_8_15_reset = reset;
assign left_8_15_in = left_8_14_out;
assign pe_9_3_mul_ready =
  _guard1744 ? 1'd1 :
  _guard1747 ? 1'd0 :
  1'd0;
assign pe_9_3_clk = clk;
assign pe_9_3_top =
  _guard1760 ? top_9_3_out :
  32'd0;
assign pe_9_3_left =
  _guard1773 ? left_9_3_out :
  32'd0;
assign pe_9_3_reset = reset;
assign pe_9_3_go = _guard1786;
assign pe_9_11_mul_ready =
  _guard1789 ? 1'd1 :
  _guard1792 ? 1'd0 :
  1'd0;
assign pe_9_11_clk = clk;
assign pe_9_11_top =
  _guard1805 ? top_9_11_out :
  32'd0;
assign pe_9_11_left =
  _guard1818 ? left_9_11_out :
  32'd0;
assign pe_9_11_reset = reset;
assign pe_9_11_go = _guard1831;
assign left_9_13_write_en = _guard1834;
assign left_9_13_clk = clk;
assign left_9_13_reset = reset;
assign left_9_13_in = left_9_12_out;
assign top_9_14_write_en = _guard1840;
assign top_9_14_clk = clk;
assign top_9_14_reset = reset;
assign top_9_14_in = top_8_14_out;
assign left_10_0_write_en = _guard1846;
assign left_10_0_clk = clk;
assign left_10_0_reset = reset;
assign left_10_0_in = l10_read_data;
assign left_10_4_write_en = _guard1852;
assign left_10_4_clk = clk;
assign left_10_4_reset = reset;
assign left_10_4_in = left_10_3_out;
assign top_10_7_write_en = _guard1858;
assign top_10_7_clk = clk;
assign top_10_7_reset = reset;
assign top_10_7_in = top_9_7_out;
assign left_11_2_write_en = _guard1864;
assign left_11_2_clk = clk;
assign left_11_2_reset = reset;
assign left_11_2_in = left_11_1_out;
assign pe_11_5_mul_ready =
  _guard1870 ? 1'd1 :
  _guard1873 ? 1'd0 :
  1'd0;
assign pe_11_5_clk = clk;
assign pe_11_5_top =
  _guard1886 ? top_11_5_out :
  32'd0;
assign pe_11_5_left =
  _guard1899 ? left_11_5_out :
  32'd0;
assign pe_11_5_reset = reset;
assign pe_11_5_go = _guard1912;
assign left_11_5_write_en = _guard1915;
assign left_11_5_clk = clk;
assign left_11_5_reset = reset;
assign left_11_5_in = left_11_4_out;
assign left_11_10_write_en = _guard1921;
assign left_11_10_clk = clk;
assign left_11_10_reset = reset;
assign left_11_10_in = left_11_9_out;
assign pe_11_12_mul_ready =
  _guard1927 ? 1'd1 :
  _guard1930 ? 1'd0 :
  1'd0;
assign pe_11_12_clk = clk;
assign pe_11_12_top =
  _guard1943 ? top_11_12_out :
  32'd0;
assign pe_11_12_left =
  _guard1956 ? left_11_12_out :
  32'd0;
assign pe_11_12_reset = reset;
assign pe_11_12_go = _guard1969;
assign left_12_10_write_en = _guard1972;
assign left_12_10_clk = clk;
assign left_12_10_reset = reset;
assign left_12_10_in = left_12_9_out;
assign left_13_9_write_en = _guard1978;
assign left_13_9_clk = clk;
assign left_13_9_reset = reset;
assign left_13_9_in = left_13_8_out;
assign pe_13_10_mul_ready =
  _guard1984 ? 1'd1 :
  _guard1987 ? 1'd0 :
  1'd0;
assign pe_13_10_clk = clk;
assign pe_13_10_top =
  _guard2000 ? top_13_10_out :
  32'd0;
assign pe_13_10_left =
  _guard2013 ? left_13_10_out :
  32'd0;
assign pe_13_10_reset = reset;
assign pe_13_10_go = _guard2026;
assign top_15_1_write_en = _guard2029;
assign top_15_1_clk = clk;
assign top_15_1_reset = reset;
assign top_15_1_in = top_14_1_out;
assign t8_idx_write_en = _guard2039;
assign t8_idx_clk = clk;
assign t8_idx_reset = reset;
assign t8_idx_in =
  _guard2042 ? 5'd0 :
  _guard2045 ? t8_add_out :
  'x;
assign t11_idx_write_en = _guard2052;
assign t11_idx_clk = clk;
assign t11_idx_reset = reset;
assign t11_idx_in =
  _guard2055 ? 5'd0 :
  _guard2058 ? t11_add_out :
  'x;
assign l3_idx_write_en = _guard2065;
assign l3_idx_clk = clk;
assign l3_idx_reset = reset;
assign l3_idx_in =
  _guard2068 ? l3_add_out :
  _guard2071 ? 5'd0 :
  'x;
assign l7_idx_write_en = _guard2078;
assign l7_idx_clk = clk;
assign l7_idx_reset = reset;
assign l7_idx_in =
  _guard2081 ? 5'd0 :
  _guard2084 ? l7_add_out :
  'x;
assign l10_idx_write_en = _guard2091;
assign l10_idx_clk = clk;
assign l10_idx_reset = reset;
assign l10_idx_in =
  _guard2094 ? 5'd0 :
  _guard2097 ? l10_add_out :
  'x;
assign idx_between_30_46_reg_write_en = _guard2102;
assign idx_between_30_46_reg_clk = clk;
assign idx_between_30_46_reg_reset = reset;
assign idx_between_30_46_reg_in =
  _guard2103 ? idx_between_30_46_comb_out :
  _guard2106 ? 1'd0 :
  'x;
assign index_lt_17_left = idx_add_out;
assign index_lt_17_right = 6'd17;
assign index_ge_42_left = idx_add_out;
assign index_ge_42_right = 6'd42;
assign index_lt_34_left = idx_add_out;
assign index_lt_34_right = 6'd34;
assign idx_between_27_31_comb_left = index_ge_27_out;
assign idx_between_27_31_comb_right = index_lt_31_out;
assign index_ge_51_left = idx_add_out;
assign index_ge_51_right = 6'd51;
assign index_ge_14_left = idx_add_out;
assign index_ge_14_right = 6'd14;
assign idx_between_28_32_comb_left = index_ge_28_out;
assign idx_between_28_32_comb_right = index_lt_32_out;
assign idx_between_6_22_reg_write_en = _guard2125;
assign idx_between_6_22_reg_clk = clk;
assign idx_between_6_22_reg_reset = reset;
assign idx_between_6_22_reg_in =
  _guard2126 ? idx_between_6_22_comb_out :
  _guard2129 ? 1'd0 :
  'x;
assign idx_between_34_50_comb_left = index_ge_34_out;
assign idx_between_34_50_comb_right = index_lt_50_out;
assign idx_between_25_26_reg_write_en = _guard2136;
assign idx_between_25_26_reg_clk = clk;
assign idx_between_25_26_reg_reset = reset;
assign idx_between_25_26_reg_in =
  _guard2139 ? 1'd0 :
  _guard2140 ? idx_between_25_26_comb_out :
  'x;
assign idx_between_26_27_reg_write_en = _guard2145;
assign idx_between_26_27_reg_clk = clk;
assign idx_between_26_27_reg_reset = reset;
assign idx_between_26_27_reg_in =
  _guard2146 ? idx_between_26_27_comb_out :
  _guard2149 ? 1'd0 :
  'x;
assign index_ge_8_left = idx_add_out;
assign index_ge_8_right = 6'd8;
assign idx_between_18_34_comb_left = index_ge_18_out;
assign idx_between_18_34_comb_right = index_lt_34_out;
assign idx_between_6_10_reg_write_en = _guard2158;
assign idx_between_6_10_reg_clk = clk;
assign idx_between_6_10_reg_reset = reset;
assign idx_between_6_10_reg_in =
  _guard2159 ? idx_between_6_10_comb_out :
  _guard2162 ? 1'd0 :
  'x;
assign idx_between_16_32_reg_write_en = _guard2167;
assign idx_between_16_32_reg_clk = clk;
assign idx_between_16_32_reg_reset = reset;
assign idx_between_16_32_reg_in =
  _guard2168 ? idx_between_16_32_comb_out :
  _guard2171 ? 1'd0 :
  'x;
assign idx_between_16_32_comb_left = index_ge_16_out;
assign idx_between_16_32_comb_right = index_lt_32_out;
assign idx_between_22_38_comb_left = index_ge_22_out;
assign idx_between_22_38_comb_right = index_lt_38_out;
assign idx_between_17_33_reg_write_en = _guard2180;
assign idx_between_17_33_reg_clk = clk;
assign idx_between_17_33_reg_reset = reset;
assign idx_between_17_33_reg_in =
  _guard2181 ? idx_between_17_33_comb_out :
  _guard2184 ? 1'd0 :
  'x;
assign idx_between_13_29_comb_left = index_ge_13_out;
assign idx_between_13_29_comb_right = index_lt_29_out;
assign index_lt_13_left = idx_add_out;
assign index_lt_13_right = 6'd13;
assign idx_between_33_34_comb_left = index_ge_33_out;
assign idx_between_33_34_comb_right = index_lt_34_out;
assign idx_between_43_44_reg_write_en = _guard2195;
assign idx_between_43_44_reg_clk = clk;
assign idx_between_43_44_reg_reset = reset;
assign idx_between_43_44_reg_in =
  _guard2198 ? 1'd0 :
  _guard2199 ? idx_between_43_44_comb_out :
  'x;
assign done = _guard2200;
assign t2_addr0 =
  _guard2203 ? t2_idx_out :
  5'd0;
assign t3_reset = reset;
assign t10_reset = reset;
assign t12_reset = reset;
assign t13_addr0 =
  _guard2206 ? t13_idx_out :
  5'd0;
assign t13_reset = reset;
assign l15_addr0 =
  _guard2209 ? l15_idx_out :
  5'd0;
assign out_mem_4_write_data =
  _guard2212 ? pe_4_9_out :
  _guard2215 ? pe_4_0_out :
  _guard2218 ? pe_4_5_out :
  _guard2221 ? pe_4_12_out :
  _guard2224 ? pe_4_14_out :
  _guard2227 ? pe_4_15_out :
  _guard2230 ? pe_4_6_out :
  _guard2233 ? pe_4_11_out :
  _guard2236 ? pe_4_2_out :
  _guard2239 ? pe_4_8_out :
  _guard2242 ? pe_4_4_out :
  _guard2245 ? pe_4_7_out :
  _guard2248 ? pe_4_13_out :
  _guard2251 ? pe_4_3_out :
  _guard2254 ? pe_4_10_out :
  _guard2257 ? pe_4_1_out :
  32'd0;
assign out_mem_9_reset = reset;
assign out_mem_12_addr0 =
  _guard2260 ? 5'd1 :
  _guard2263 ? 5'd15 :
  _guard2266 ? 5'd0 :
  _guard2269 ? 5'd3 :
  _guard2272 ? 5'd13 :
  _guard2275 ? 5'd14 :
  _guard2278 ? 5'd5 :
  _guard2281 ? 5'd12 :
  _guard2284 ? 5'd2 :
  _guard2287 ? 5'd8 :
  _guard2290 ? 5'd10 :
  _guard2293 ? 5'd7 :
  _guard2296 ? 5'd11 :
  _guard2299 ? 5'd4 :
  _guard2302 ? 5'd6 :
  _guard2305 ? 5'd9 :
  5'd0;
assign out_mem_15_reset = reset;
assign t0_reset = reset;
assign t6_reset = reset;
assign t15_reset = reset;
assign l5_addr0 =
  _guard2308 ? l5_idx_out :
  5'd0;
assign l5_clk = clk;
assign l9_reset = reset;
assign out_mem_2_reset = reset;
assign out_mem_8_reset = reset;
assign out_mem_12_reset = reset;
assign out_mem_14_reset = reset;
assign out_mem_15_addr0 =
  _guard2311 ? 5'd1 :
  _guard2314 ? 5'd15 :
  _guard2317 ? 5'd0 :
  _guard2320 ? 5'd3 :
  _guard2323 ? 5'd13 :
  _guard2326 ? 5'd14 :
  _guard2329 ? 5'd5 :
  _guard2332 ? 5'd12 :
  _guard2335 ? 5'd2 :
  _guard2338 ? 5'd8 :
  _guard2341 ? 5'd10 :
  _guard2344 ? 5'd7 :
  _guard2347 ? 5'd11 :
  _guard2350 ? 5'd4 :
  _guard2353 ? 5'd6 :
  _guard2356 ? 5'd9 :
  5'd0;
assign t2_clk = clk;
assign t12_clk = clk;
assign l0_addr0 =
  _guard2359 ? l0_idx_out :
  5'd0;
assign l3_clk = clk;
assign out_mem_1_addr0 =
  _guard2362 ? 5'd1 :
  _guard2365 ? 5'd15 :
  _guard2368 ? 5'd0 :
  _guard2371 ? 5'd3 :
  _guard2374 ? 5'd13 :
  _guard2377 ? 5'd14 :
  _guard2380 ? 5'd5 :
  _guard2383 ? 5'd12 :
  _guard2386 ? 5'd2 :
  _guard2389 ? 5'd8 :
  _guard2392 ? 5'd10 :
  _guard2395 ? 5'd7 :
  _guard2398 ? 5'd11 :
  _guard2401 ? 5'd4 :
  _guard2404 ? 5'd6 :
  _guard2407 ? 5'd9 :
  5'd0;
assign out_mem_1_clk = clk;
assign out_mem_3_reset = reset;
assign out_mem_5_addr0 =
  _guard2410 ? 5'd1 :
  _guard2413 ? 5'd15 :
  _guard2416 ? 5'd0 :
  _guard2419 ? 5'd3 :
  _guard2422 ? 5'd13 :
  _guard2425 ? 5'd14 :
  _guard2428 ? 5'd5 :
  _guard2431 ? 5'd12 :
  _guard2434 ? 5'd2 :
  _guard2437 ? 5'd8 :
  _guard2440 ? 5'd10 :
  _guard2443 ? 5'd7 :
  _guard2446 ? 5'd11 :
  _guard2449 ? 5'd4 :
  _guard2452 ? 5'd6 :
  _guard2455 ? 5'd9 :
  5'd0;
assign out_mem_5_write_data =
  _guard2458 ? pe_5_2_out :
  _guard2461 ? pe_5_8_out :
  _guard2464 ? pe_5_13_out :
  _guard2467 ? pe_5_0_out :
  _guard2470 ? pe_5_4_out :
  _guard2473 ? pe_5_1_out :
  _guard2476 ? pe_5_7_out :
  _guard2479 ? pe_5_9_out :
  _guard2482 ? pe_5_10_out :
  _guard2485 ? pe_5_3_out :
  _guard2488 ? pe_5_5_out :
  _guard2491 ? pe_5_14_out :
  _guard2494 ? pe_5_6_out :
  _guard2497 ? pe_5_11_out :
  _guard2500 ? pe_5_15_out :
  _guard2503 ? pe_5_12_out :
  32'd0;
assign out_mem_11_addr0 =
  _guard2506 ? 5'd1 :
  _guard2509 ? 5'd15 :
  _guard2512 ? 5'd0 :
  _guard2515 ? 5'd3 :
  _guard2518 ? 5'd13 :
  _guard2521 ? 5'd14 :
  _guard2524 ? 5'd5 :
  _guard2527 ? 5'd12 :
  _guard2530 ? 5'd2 :
  _guard2533 ? 5'd8 :
  _guard2536 ? 5'd10 :
  _guard2539 ? 5'd7 :
  _guard2542 ? 5'd11 :
  _guard2545 ? 5'd4 :
  _guard2548 ? 5'd6 :
  _guard2551 ? 5'd9 :
  5'd0;
assign out_mem_13_reset = reset;
assign t15_clk = clk;
assign l6_addr0 =
  _guard2554 ? l6_idx_out :
  5'd0;
assign l13_reset = reset;
assign out_mem_0_write_data =
  _guard2557 ? pe_0_10_out :
  _guard2560 ? pe_0_1_out :
  _guard2563 ? pe_0_7_out :
  _guard2566 ? pe_0_3_out :
  _guard2569 ? pe_0_5_out :
  _guard2572 ? pe_0_8_out :
  _guard2575 ? pe_0_9_out :
  _guard2578 ? pe_0_2_out :
  _guard2581 ? pe_0_12_out :
  _guard2584 ? pe_0_15_out :
  _guard2587 ? pe_0_4_out :
  _guard2590 ? pe_0_14_out :
  _guard2593 ? pe_0_11_out :
  _guard2596 ? pe_0_0_out :
  _guard2599 ? pe_0_6_out :
  _guard2602 ? pe_0_13_out :
  32'd0;
assign out_mem_5_clk = clk;
assign out_mem_8_clk = clk;
assign out_mem_12_write_data =
  _guard2605 ? pe_12_10_out :
  _guard2608 ? pe_12_9_out :
  _guard2611 ? pe_12_12_out :
  _guard2614 ? pe_12_3_out :
  _guard2617 ? pe_12_4_out :
  _guard2620 ? pe_12_1_out :
  _guard2623 ? pe_12_7_out :
  _guard2626 ? pe_12_11_out :
  _guard2629 ? pe_12_6_out :
  _guard2632 ? pe_12_5_out :
  _guard2635 ? pe_12_13_out :
  _guard2638 ? pe_12_15_out :
  _guard2641 ? pe_12_0_out :
  _guard2644 ? pe_12_2_out :
  _guard2647 ? pe_12_8_out :
  _guard2650 ? pe_12_14_out :
  32'd0;
assign out_mem_14_clk = clk;
assign t5_reset = reset;
assign t14_clk = clk;
assign l7_reset = reset;
assign l8_reset = reset;
assign l10_reset = reset;
assign l11_reset = reset;
assign l13_addr0 =
  _guard2653 ? l13_idx_out :
  5'd0;
assign out_mem_6_addr0 =
  _guard2656 ? 5'd1 :
  _guard2659 ? 5'd15 :
  _guard2662 ? 5'd0 :
  _guard2665 ? 5'd3 :
  _guard2668 ? 5'd13 :
  _guard2671 ? 5'd14 :
  _guard2674 ? 5'd5 :
  _guard2677 ? 5'd12 :
  _guard2680 ? 5'd2 :
  _guard2683 ? 5'd8 :
  _guard2686 ? 5'd10 :
  _guard2689 ? 5'd7 :
  _guard2692 ? 5'd11 :
  _guard2695 ? 5'd4 :
  _guard2698 ? 5'd6 :
  _guard2701 ? 5'd9 :
  5'd0;
assign t0_clk = clk;
assign l5_reset = reset;
assign l11_addr0 =
  _guard2704 ? l11_idx_out :
  5'd0;
assign l14_addr0 =
  _guard2707 ? l14_idx_out :
  5'd0;
assign out_mem_1_reset = reset;
assign out_mem_3_write_data =
  _guard2710 ? pe_3_8_out :
  _guard2713 ? pe_3_4_out :
  _guard2716 ? pe_3_7_out :
  _guard2719 ? pe_3_15_out :
  _guard2722 ? pe_3_2_out :
  _guard2725 ? pe_3_5_out :
  _guard2728 ? pe_3_6_out :
  _guard2731 ? pe_3_0_out :
  _guard2734 ? pe_3_13_out :
  _guard2737 ? pe_3_14_out :
  _guard2740 ? pe_3_1_out :
  _guard2743 ? pe_3_10_out :
  _guard2746 ? pe_3_9_out :
  _guard2749 ? pe_3_11_out :
  _guard2752 ? pe_3_12_out :
  _guard2755 ? pe_3_3_out :
  32'd0;
assign out_mem_9_write_en = _guard2852;
assign out_mem_10_write_data =
  _guard2855 ? pe_10_5_out :
  _guard2858 ? pe_10_7_out :
  _guard2861 ? pe_10_9_out :
  _guard2864 ? pe_10_8_out :
  _guard2867 ? pe_10_13_out :
  _guard2870 ? pe_10_12_out :
  _guard2873 ? pe_10_0_out :
  _guard2876 ? pe_10_14_out :
  _guard2879 ? pe_10_10_out :
  _guard2882 ? pe_10_2_out :
  _guard2885 ? pe_10_3_out :
  _guard2888 ? pe_10_4_out :
  _guard2891 ? pe_10_15_out :
  _guard2894 ? pe_10_11_out :
  _guard2897 ? pe_10_1_out :
  _guard2900 ? pe_10_6_out :
  32'd0;
assign out_mem_12_write_en = _guard2997;
assign t4_reset = reset;
assign t5_addr0 =
  _guard3000 ? t5_idx_out :
  5'd0;
assign t5_clk = clk;
assign t6_clk = clk;
assign t15_addr0 =
  _guard3003 ? t15_idx_out :
  5'd0;
assign l0_reset = reset;
assign l1_addr0 =
  _guard3006 ? l1_idx_out :
  5'd0;
assign l7_clk = clk;
assign out_mem_5_write_en = _guard3103;
assign out_mem_5_reset = reset;
assign out_mem_7_addr0 =
  _guard3106 ? 5'd1 :
  _guard3109 ? 5'd15 :
  _guard3112 ? 5'd0 :
  _guard3115 ? 5'd3 :
  _guard3118 ? 5'd13 :
  _guard3121 ? 5'd14 :
  _guard3124 ? 5'd5 :
  _guard3127 ? 5'd12 :
  _guard3130 ? 5'd2 :
  _guard3133 ? 5'd8 :
  _guard3136 ? 5'd10 :
  _guard3139 ? 5'd7 :
  _guard3142 ? 5'd11 :
  _guard3145 ? 5'd4 :
  _guard3148 ? 5'd6 :
  _guard3151 ? 5'd9 :
  5'd0;
assign out_mem_9_addr0 =
  _guard3154 ? 5'd1 :
  _guard3157 ? 5'd15 :
  _guard3160 ? 5'd0 :
  _guard3163 ? 5'd3 :
  _guard3166 ? 5'd13 :
  _guard3169 ? 5'd14 :
  _guard3172 ? 5'd5 :
  _guard3175 ? 5'd12 :
  _guard3178 ? 5'd2 :
  _guard3181 ? 5'd8 :
  _guard3184 ? 5'd10 :
  _guard3187 ? 5'd7 :
  _guard3190 ? 5'd11 :
  _guard3193 ? 5'd4 :
  _guard3196 ? 5'd6 :
  _guard3199 ? 5'd9 :
  5'd0;
assign out_mem_13_write_en = _guard3296;
assign t4_clk = clk;
assign t10_clk = clk;
assign t14_addr0 =
  _guard3299 ? t14_idx_out :
  5'd0;
assign l14_clk = clk;
assign out_mem_10_addr0 =
  _guard3302 ? 5'd1 :
  _guard3305 ? 5'd15 :
  _guard3308 ? 5'd0 :
  _guard3311 ? 5'd3 :
  _guard3314 ? 5'd13 :
  _guard3317 ? 5'd14 :
  _guard3320 ? 5'd5 :
  _guard3323 ? 5'd12 :
  _guard3326 ? 5'd2 :
  _guard3329 ? 5'd8 :
  _guard3332 ? 5'd10 :
  _guard3335 ? 5'd7 :
  _guard3338 ? 5'd11 :
  _guard3341 ? 5'd4 :
  _guard3344 ? 5'd6 :
  _guard3347 ? 5'd9 :
  5'd0;
assign out_mem_11_clk = clk;
assign out_mem_13_clk = clk;
assign t4_addr0 =
  _guard3350 ? t4_idx_out :
  5'd0;
assign t6_addr0 =
  _guard3353 ? t6_idx_out :
  5'd0;
assign t8_reset = reset;
assign t12_addr0 =
  _guard3356 ? t12_idx_out :
  5'd0;
assign l15_clk = clk;
assign l15_reset = reset;
assign out_mem_0_clk = clk;
assign out_mem_7_write_en = _guard3453;
assign out_mem_7_clk = clk;
assign out_mem_7_reset = reset;
assign out_mem_10_reset = reset;
assign t1_reset = reset;
assign t8_addr0 =
  _guard3456 ? t8_idx_out :
  5'd0;
assign t13_clk = clk;
assign l6_clk = clk;
assign l9_clk = clk;
assign out_mem_3_clk = clk;
assign out_mem_4_addr0 =
  _guard3459 ? 5'd1 :
  _guard3462 ? 5'd15 :
  _guard3465 ? 5'd0 :
  _guard3468 ? 5'd3 :
  _guard3471 ? 5'd13 :
  _guard3474 ? 5'd14 :
  _guard3477 ? 5'd5 :
  _guard3480 ? 5'd12 :
  _guard3483 ? 5'd2 :
  _guard3486 ? 5'd8 :
  _guard3489 ? 5'd10 :
  _guard3492 ? 5'd7 :
  _guard3495 ? 5'd11 :
  _guard3498 ? 5'd4 :
  _guard3501 ? 5'd6 :
  _guard3504 ? 5'd9 :
  5'd0;
assign out_mem_4_clk = clk;
assign out_mem_4_reset = reset;
assign out_mem_6_reset = reset;
assign out_mem_9_clk = clk;
assign out_mem_11_write_en = _guard3601;
assign t7_clk = clk;
assign t8_clk = clk;
assign t9_addr0 =
  _guard3604 ? t9_idx_out :
  5'd0;
assign t9_reset = reset;
assign t14_reset = reset;
assign l3_addr0 =
  _guard3607 ? l3_idx_out :
  5'd0;
assign l4_reset = reset;
assign l10_addr0 =
  _guard3610 ? l10_idx_out :
  5'd0;
assign l12_clk = clk;
assign out_mem_2_write_data =
  _guard3613 ? pe_2_12_out :
  _guard3616 ? pe_2_11_out :
  _guard3619 ? pe_2_14_out :
  _guard3622 ? pe_2_7_out :
  _guard3625 ? pe_2_13_out :
  _guard3628 ? pe_2_4_out :
  _guard3631 ? pe_2_15_out :
  _guard3634 ? pe_2_1_out :
  _guard3637 ? pe_2_3_out :
  _guard3640 ? pe_2_5_out :
  _guard3643 ? pe_2_6_out :
  _guard3646 ? pe_2_8_out :
  _guard3649 ? pe_2_0_out :
  _guard3652 ? pe_2_2_out :
  _guard3655 ? pe_2_9_out :
  _guard3658 ? pe_2_10_out :
  32'd0;
assign out_mem_11_reset = reset;
assign out_mem_12_clk = clk;
assign out_mem_15_clk = clk;
assign t9_clk = clk;
assign t11_clk = clk;
assign l4_addr0 =
  _guard3661 ? l4_idx_out :
  5'd0;
assign l7_addr0 =
  _guard3664 ? l7_idx_out :
  5'd0;
assign out_mem_0_reset = reset;
assign out_mem_1_write_data =
  _guard3667 ? pe_1_4_out :
  _guard3670 ? pe_1_7_out :
  _guard3673 ? pe_1_2_out :
  _guard3676 ? pe_1_3_out :
  _guard3679 ? pe_1_8_out :
  _guard3682 ? pe_1_15_out :
  _guard3685 ? pe_1_0_out :
  _guard3688 ? pe_1_6_out :
  _guard3691 ? pe_1_12_out :
  _guard3694 ? pe_1_5_out :
  _guard3697 ? pe_1_9_out :
  _guard3700 ? pe_1_11_out :
  _guard3703 ? pe_1_1_out :
  _guard3706 ? pe_1_13_out :
  _guard3709 ? pe_1_10_out :
  _guard3712 ? pe_1_14_out :
  32'd0;
assign out_mem_1_write_en = _guard3809;
assign out_mem_4_write_en = _guard3906;
assign out_mem_6_clk = clk;
assign t0_addr0 =
  _guard3909 ? t0_idx_out :
  5'd0;
assign t1_addr0 =
  _guard3912 ? t1_idx_out :
  5'd0;
assign t1_clk = clk;
assign t11_addr0 =
  _guard3915 ? t11_idx_out :
  5'd0;
assign l1_reset = reset;
assign l2_clk = clk;
assign l2_reset = reset;
assign l11_clk = clk;
assign out_mem_0_write_en = _guard4012;
assign out_mem_2_write_en = _guard4109;
assign out_mem_2_clk = clk;
assign t3_clk = clk;
assign t7_reset = reset;
assign t11_reset = reset;
assign l8_addr0 =
  _guard4112 ? l8_idx_out :
  5'd0;
assign l10_clk = clk;
assign out_mem_3_write_en = _guard4209;
assign out_mem_6_write_data =
  _guard4212 ? pe_6_4_out :
  _guard4215 ? pe_6_11_out :
  _guard4218 ? pe_6_0_out :
  _guard4221 ? pe_6_1_out :
  _guard4224 ? pe_6_5_out :
  _guard4227 ? pe_6_12_out :
  _guard4230 ? pe_6_2_out :
  _guard4233 ? pe_6_3_out :
  _guard4236 ? pe_6_10_out :
  _guard4239 ? pe_6_7_out :
  _guard4242 ? pe_6_13_out :
  _guard4245 ? pe_6_14_out :
  _guard4248 ? pe_6_15_out :
  _guard4251 ? pe_6_6_out :
  _guard4254 ? pe_6_8_out :
  _guard4257 ? pe_6_9_out :
  32'd0;
assign out_mem_6_write_en = _guard4354;
assign out_mem_7_write_data =
  _guard4357 ? pe_7_9_out :
  _guard4360 ? pe_7_3_out :
  _guard4363 ? pe_7_15_out :
  _guard4366 ? pe_7_4_out :
  _guard4369 ? pe_7_0_out :
  _guard4372 ? pe_7_10_out :
  _guard4375 ? pe_7_5_out :
  _guard4378 ? pe_7_6_out :
  _guard4381 ? pe_7_14_out :
  _guard4384 ? pe_7_1_out :
  _guard4387 ? pe_7_12_out :
  _guard4390 ? pe_7_2_out :
  _guard4393 ? pe_7_7_out :
  _guard4396 ? pe_7_8_out :
  _guard4399 ? pe_7_11_out :
  _guard4402 ? pe_7_13_out :
  32'd0;
assign out_mem_10_write_en = _guard4499;
assign out_mem_14_write_en = _guard4596;
assign t10_addr0 =
  _guard4599 ? t10_idx_out :
  5'd0;
assign l0_clk = clk;
assign l1_clk = clk;
assign l2_addr0 =
  _guard4602 ? l2_idx_out :
  5'd0;
assign l3_reset = reset;
assign l4_clk = clk;
assign l6_reset = reset;
assign l9_addr0 =
  _guard4605 ? l9_idx_out :
  5'd0;
assign l12_addr0 =
  _guard4608 ? l12_idx_out :
  5'd0;
assign l14_reset = reset;
assign out_mem_0_addr0 =
  _guard4611 ? 5'd1 :
  _guard4614 ? 5'd15 :
  _guard4617 ? 5'd0 :
  _guard4620 ? 5'd3 :
  _guard4623 ? 5'd13 :
  _guard4626 ? 5'd14 :
  _guard4629 ? 5'd5 :
  _guard4632 ? 5'd12 :
  _guard4635 ? 5'd2 :
  _guard4638 ? 5'd8 :
  _guard4641 ? 5'd10 :
  _guard4644 ? 5'd7 :
  _guard4647 ? 5'd11 :
  _guard4650 ? 5'd4 :
  _guard4653 ? 5'd6 :
  _guard4656 ? 5'd9 :
  5'd0;
assign out_mem_3_addr0 =
  _guard4659 ? 5'd1 :
  _guard4662 ? 5'd15 :
  _guard4665 ? 5'd0 :
  _guard4668 ? 5'd3 :
  _guard4671 ? 5'd13 :
  _guard4674 ? 5'd14 :
  _guard4677 ? 5'd5 :
  _guard4680 ? 5'd12 :
  _guard4683 ? 5'd2 :
  _guard4686 ? 5'd8 :
  _guard4689 ? 5'd10 :
  _guard4692 ? 5'd7 :
  _guard4695 ? 5'd11 :
  _guard4698 ? 5'd4 :
  _guard4701 ? 5'd6 :
  _guard4704 ? 5'd9 :
  5'd0;
assign out_mem_8_addr0 =
  _guard4707 ? 5'd1 :
  _guard4710 ? 5'd15 :
  _guard4713 ? 5'd0 :
  _guard4716 ? 5'd3 :
  _guard4719 ? 5'd13 :
  _guard4722 ? 5'd14 :
  _guard4725 ? 5'd5 :
  _guard4728 ? 5'd12 :
  _guard4731 ? 5'd2 :
  _guard4734 ? 5'd8 :
  _guard4737 ? 5'd10 :
  _guard4740 ? 5'd7 :
  _guard4743 ? 5'd11 :
  _guard4746 ? 5'd4 :
  _guard4749 ? 5'd6 :
  _guard4752 ? 5'd9 :
  5'd0;
assign out_mem_10_clk = clk;
assign out_mem_11_write_data =
  _guard4755 ? pe_11_5_out :
  _guard4758 ? pe_11_12_out :
  _guard4761 ? pe_11_8_out :
  _guard4764 ? pe_11_15_out :
  _guard4767 ? pe_11_4_out :
  _guard4770 ? pe_11_0_out :
  _guard4773 ? pe_11_11_out :
  _guard4776 ? pe_11_6_out :
  _guard4779 ? pe_11_7_out :
  _guard4782 ? pe_11_9_out :
  _guard4785 ? pe_11_2_out :
  _guard4788 ? pe_11_3_out :
  _guard4791 ? pe_11_1_out :
  _guard4794 ? pe_11_13_out :
  _guard4797 ? pe_11_14_out :
  _guard4800 ? pe_11_10_out :
  32'd0;
assign t2_reset = reset;
assign t3_addr0 =
  _guard4803 ? t3_idx_out :
  5'd0;
assign t7_addr0 =
  _guard4806 ? t7_idx_out :
  5'd0;
assign l8_clk = clk;
assign l12_reset = reset;
assign l13_clk = clk;
assign out_mem_2_addr0 =
  _guard4809 ? 5'd1 :
  _guard4812 ? 5'd15 :
  _guard4815 ? 5'd0 :
  _guard4818 ? 5'd3 :
  _guard4821 ? 5'd13 :
  _guard4824 ? 5'd14 :
  _guard4827 ? 5'd5 :
  _guard4830 ? 5'd12 :
  _guard4833 ? 5'd2 :
  _guard4836 ? 5'd8 :
  _guard4839 ? 5'd10 :
  _guard4842 ? 5'd7 :
  _guard4845 ? 5'd11 :
  _guard4848 ? 5'd4 :
  _guard4851 ? 5'd6 :
  _guard4854 ? 5'd9 :
  5'd0;
assign out_mem_8_write_data =
  _guard4857 ? pe_8_6_out :
  _guard4860 ? pe_8_13_out :
  _guard4863 ? pe_8_1_out :
  _guard4866 ? pe_8_2_out :
  _guard4869 ? pe_8_4_out :
  _guard4872 ? pe_8_0_out :
  _guard4875 ? pe_8_5_out :
  _guard4878 ? pe_8_9_out :
  _guard4881 ? pe_8_15_out :
  _guard4884 ? pe_8_11_out :
  _guard4887 ? pe_8_3_out :
  _guard4890 ? pe_8_12_out :
  _guard4893 ? pe_8_10_out :
  _guard4896 ? pe_8_14_out :
  _guard4899 ? pe_8_7_out :
  _guard4902 ? pe_8_8_out :
  32'd0;
assign out_mem_8_write_en = _guard4999;
assign out_mem_9_write_data =
  _guard5002 ? pe_9_15_out :
  _guard5005 ? pe_9_3_out :
  _guard5008 ? pe_9_11_out :
  _guard5011 ? pe_9_7_out :
  _guard5014 ? pe_9_9_out :
  _guard5017 ? pe_9_13_out :
  _guard5020 ? pe_9_6_out :
  _guard5023 ? pe_9_10_out :
  _guard5026 ? pe_9_12_out :
  _guard5029 ? pe_9_0_out :
  _guard5032 ? pe_9_4_out :
  _guard5035 ? pe_9_5_out :
  _guard5038 ? pe_9_1_out :
  _guard5041 ? pe_9_8_out :
  _guard5044 ? pe_9_14_out :
  _guard5047 ? pe_9_2_out :
  32'd0;
assign out_mem_13_addr0 =
  _guard5050 ? 5'd1 :
  _guard5053 ? 5'd15 :
  _guard5056 ? 5'd0 :
  _guard5059 ? 5'd3 :
  _guard5062 ? 5'd13 :
  _guard5065 ? 5'd14 :
  _guard5068 ? 5'd5 :
  _guard5071 ? 5'd12 :
  _guard5074 ? 5'd2 :
  _guard5077 ? 5'd8 :
  _guard5080 ? 5'd10 :
  _guard5083 ? 5'd7 :
  _guard5086 ? 5'd11 :
  _guard5089 ? 5'd4 :
  _guard5092 ? 5'd6 :
  _guard5095 ? 5'd9 :
  5'd0;
assign out_mem_13_write_data =
  _guard5098 ? pe_13_14_out :
  _guard5101 ? pe_13_10_out :
  _guard5104 ? pe_13_7_out :
  _guard5107 ? pe_13_0_out :
  _guard5110 ? pe_13_3_out :
  _guard5113 ? pe_13_13_out :
  _guard5116 ? pe_13_5_out :
  _guard5119 ? pe_13_6_out :
  _guard5122 ? pe_13_8_out :
  _guard5125 ? pe_13_12_out :
  _guard5128 ? pe_13_1_out :
  _guard5131 ? pe_13_11_out :
  _guard5134 ? pe_13_4_out :
  _guard5137 ? pe_13_9_out :
  _guard5140 ? pe_13_15_out :
  _guard5143 ? pe_13_2_out :
  32'd0;
assign out_mem_14_addr0 =
  _guard5146 ? 5'd1 :
  _guard5149 ? 5'd15 :
  _guard5152 ? 5'd0 :
  _guard5155 ? 5'd3 :
  _guard5158 ? 5'd13 :
  _guard5161 ? 5'd14 :
  _guard5164 ? 5'd5 :
  _guard5167 ? 5'd12 :
  _guard5170 ? 5'd2 :
  _guard5173 ? 5'd8 :
  _guard5176 ? 5'd10 :
  _guard5179 ? 5'd7 :
  _guard5182 ? 5'd11 :
  _guard5185 ? 5'd4 :
  _guard5188 ? 5'd6 :
  _guard5191 ? 5'd9 :
  5'd0;
assign out_mem_14_write_data =
  _guard5194 ? pe_14_13_out :
  _guard5197 ? pe_14_1_out :
  _guard5200 ? pe_14_7_out :
  _guard5203 ? pe_14_8_out :
  _guard5206 ? pe_14_9_out :
  _guard5209 ? pe_14_14_out :
  _guard5212 ? pe_14_4_out :
  _guard5215 ? pe_14_12_out :
  _guard5218 ? pe_14_15_out :
  _guard5221 ? pe_14_0_out :
  _guard5224 ? pe_14_5_out :
  _guard5227 ? pe_14_6_out :
  _guard5230 ? pe_14_3_out :
  _guard5233 ? pe_14_10_out :
  _guard5236 ? pe_14_2_out :
  _guard5239 ? pe_14_11_out :
  32'd0;
assign out_mem_15_write_data =
  _guard5242 ? pe_15_2_out :
  _guard5245 ? pe_15_14_out :
  _guard5248 ? pe_15_9_out :
  _guard5251 ? pe_15_13_out :
  _guard5254 ? pe_15_0_out :
  _guard5257 ? pe_15_12_out :
  _guard5260 ? pe_15_11_out :
  _guard5263 ? pe_15_4_out :
  _guard5266 ? pe_15_3_out :
  _guard5269 ? pe_15_6_out :
  _guard5272 ? pe_15_15_out :
  _guard5275 ? pe_15_7_out :
  _guard5278 ? pe_15_1_out :
  _guard5281 ? pe_15_5_out :
  _guard5284 ? pe_15_10_out :
  _guard5287 ? pe_15_8_out :
  32'd0;
assign out_mem_15_write_en = _guard5384;
assign cond_wire0_in =
  _guard5385 ? idx_between_1_5_reg_out :
  _guard5388 ? cond0_out :
  1'd0;
assign cond_wire4_in =
  _guard5389 ? idx_between_1_17_reg_out :
  _guard5392 ? cond4_out :
  1'd0;
assign cond6_write_en = _guard5393;
assign cond6_clk = clk;
assign cond6_reset = reset;
assign cond6_in =
  _guard5394 ? idx_between_2_18_reg_out :
  1'd0;
assign cond_wire13_in =
  _guard5395 ? idx_between_23_24_reg_out :
  _guard5398 ? cond13_out :
  1'd0;
assign cond_wire16_in =
  _guard5401 ? cond16_out :
  _guard5402 ? idx_between_4_20_reg_out :
  1'd0;
assign cond30_write_en = _guard5403;
assign cond30_clk = clk;
assign cond30_reset = reset;
assign cond30_in =
  _guard5404 ? idx_between_7_11_reg_out :
  1'd0;
assign cond_wire32_in =
  _guard5405 ? idx_between_11_27_reg_out :
  _guard5408 ? cond32_out :
  1'd0;
assign cond_wire40_in =
  _guard5411 ? cond40_out :
  _guard5412 ? idx_between_9_13_reg_out :
  1'd0;
assign cond44_write_en = _guard5413;
assign cond44_clk = clk;
assign cond44_reset = reset;
assign cond44_in =
  _guard5414 ? idx_between_9_25_reg_out :
  1'd0;
assign cond45_write_en = _guard5415;
assign cond45_clk = clk;
assign cond45_reset = reset;
assign cond45_in =
  _guard5416 ? idx_between_10_14_reg_out :
  1'd0;
assign cond_wire73_in =
  _guard5419 ? cond73_out :
  _guard5420 ? idx_between_35_36_reg_out :
  1'd0;
assign cond81_write_en = _guard5421;
assign cond81_clk = clk;
assign cond81_reset = reset;
assign cond81_in =
  _guard5422 ? idx_between_2_18_reg_out :
  1'd0;
assign cond98_write_en = _guard5423;
assign cond98_clk = clk;
assign cond98_reset = reset;
assign cond98_in =
  _guard5424 ? idx_between_10_26_reg_out :
  1'd0;
assign cond100_write_en = _guard5425;
assign cond100_clk = clk;
assign cond100_reset = reset;
assign cond100_in =
  _guard5426 ? idx_between_7_11_reg_out :
  1'd0;
assign cond_wire101_in =
  _guard5427 ? idx_between_7_23_reg_out :
  _guard5430 ? cond101_out :
  1'd0;
assign cond107_write_en = _guard5431;
assign cond107_clk = clk;
assign cond107_reset = reset;
assign cond107_in =
  _guard5432 ? idx_between_28_29_reg_out :
  1'd0;
assign cond_wire107_in =
  _guard5435 ? cond107_out :
  _guard5436 ? idx_between_28_29_reg_out :
  1'd0;
assign cond115_write_en = _guard5437;
assign cond115_clk = clk;
assign cond115_reset = reset;
assign cond115_in =
  _guard5438 ? idx_between_30_31_reg_out :
  1'd0;
assign cond_wire121_in =
  _guard5441 ? cond121_out :
  _guard5442 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire127_in =
  _guard5445 ? cond127_out :
  _guard5446 ? idx_between_33_34_reg_out :
  1'd0;
assign cond_wire144_in =
  _guard5447 ? idx_between_2_18_reg_out :
  _guard5450 ? cond144_out :
  1'd0;
assign cond149_write_en = _guard5451;
assign cond149_clk = clk;
assign cond149_reset = reset;
assign cond149_in =
  _guard5452 ? idx_between_4_8_reg_out :
  1'd0;
assign cond150_write_en = _guard5453;
assign cond150_clk = clk;
assign cond150_reset = reset;
assign cond150_in =
  _guard5454 ? idx_between_4_20_reg_out :
  1'd0;
assign cond_wire160_in =
  _guard5455 ? idx_between_26_27_reg_out :
  _guard5458 ? cond160_out :
  1'd0;
assign cond169_write_en = _guard5459;
assign cond169_clk = clk;
assign cond169_reset = reset;
assign cond169_in =
  _guard5460 ? idx_between_9_13_reg_out :
  1'd0;
assign cond179_write_en = _guard5461;
assign cond179_clk = clk;
assign cond179_reset = reset;
assign cond179_in =
  _guard5462 ? idx_between_15_31_reg_out :
  1'd0;
assign cond193_write_en = _guard5463;
assign cond193_clk = clk;
assign cond193_reset = reset;
assign cond193_in =
  _guard5464 ? idx_between_15_19_reg_out :
  1'd0;
assign cond_wire208_in =
  _guard5467 ? cond208_out :
  _guard5468 ? idx_between_38_39_reg_out :
  1'd0;
assign cond214_write_en = _guard5469;
assign cond214_clk = clk;
assign cond214_reset = reset;
assign cond214_in =
  _guard5470 ? idx_between_5_9_reg_out :
  1'd0;
assign cond_wire230_in =
  _guard5473 ? cond230_out :
  _guard5474 ? idx_between_9_13_reg_out :
  1'd0;
assign cond236_write_en = _guard5475;
assign cond236_clk = clk;
assign cond236_reset = reset;
assign cond236_in =
  _guard5476 ? idx_between_14_30_reg_out :
  1'd0;
assign cond_wire239_in =
  _guard5477 ? idx_between_11_27_reg_out :
  _guard5480 ? cond239_out :
  1'd0;
assign cond245_write_en = _guard5481;
assign cond245_clk = clk;
assign cond245_reset = reset;
assign cond245_in =
  _guard5482 ? idx_between_32_33_reg_out :
  1'd0;
assign cond255_write_en = _guard5483;
assign cond255_clk = clk;
assign cond255_reset = reset;
assign cond255_in =
  _guard5484 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire261_in =
  _guard5485 ? idx_between_36_37_reg_out :
  _guard5488 ? cond261_out :
  1'd0;
assign cond276_write_en = _guard5489;
assign cond276_clk = clk;
assign cond276_reset = reset;
assign cond276_in =
  _guard5490 ? idx_between_5_21_reg_out :
  1'd0;
assign cond277_write_en = _guard5491;
assign cond277_clk = clk;
assign cond277_reset = reset;
assign cond277_in =
  _guard5492 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire285_in =
  _guard5493 ? idx_between_11_27_reg_out :
  _guard5496 ? cond285_out :
  1'd0;
assign cond290_write_en = _guard5497;
assign cond290_clk = clk;
assign cond290_reset = reset;
assign cond290_in =
  _guard5498 ? idx_between_28_29_reg_out :
  1'd0;
assign cond_wire321_in =
  _guard5499 ? idx_between_20_36_reg_out :
  _guard5502 ? cond321_out :
  1'd0;
assign cond_wire322_in =
  _guard5503 ? idx_between_36_37_reg_out :
  _guard5506 ? cond322_out :
  1'd0;
assign cond_wire328_in =
  _guard5507 ? idx_between_18_34_reg_out :
  _guard5510 ? cond328_out :
  1'd0;
assign cond329_write_en = _guard5511;
assign cond329_clk = clk;
assign cond329_reset = reset;
assign cond329_in =
  _guard5512 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire335_in =
  _guard5513 ? idx_between_20_24_reg_out :
  _guard5516 ? cond335_out :
  1'd0;
assign cond_wire341_in =
  _guard5517 ? idx_between_6_22_reg_out :
  _guard5520 ? cond341_out :
  1'd0;
assign cond346_write_en = _guard5521;
assign cond346_clk = clk;
assign cond346_reset = reset;
assign cond346_in =
  _guard5522 ? idx_between_11_27_reg_out :
  1'd0;
assign cond_wire346_in =
  _guard5523 ? idx_between_11_27_reg_out :
  _guard5526 ? cond346_out :
  1'd0;
assign cond_wire354_in =
  _guard5529 ? cond354_out :
  _guard5530 ? idx_between_13_29_reg_out :
  1'd0;
assign cond360_write_en = _guard5531;
assign cond360_clk = clk;
assign cond360_reset = reset;
assign cond360_in =
  _guard5532 ? idx_between_11_15_reg_out :
  1'd0;
assign cond_wire366_in =
  _guard5533 ? idx_between_16_32_reg_out :
  _guard5536 ? cond366_out :
  1'd0;
assign cond_wire371_in =
  _guard5539 ? cond371_out :
  _guard5540 ? idx_between_33_34_reg_out :
  1'd0;
assign cond382_write_en = _guard5541;
assign cond382_clk = clk;
assign cond382_reset = reset;
assign cond382_in =
  _guard5542 ? idx_between_20_36_reg_out :
  1'd0;
assign cond383_write_en = _guard5543;
assign cond383_clk = clk;
assign cond383_reset = reset;
assign cond383_in =
  _guard5544 ? idx_between_36_37_reg_out :
  1'd0;
assign cond397_write_en = _guard5545;
assign cond397_clk = clk;
assign cond397_reset = reset;
assign cond397_in =
  _guard5546 ? idx_between_20_36_reg_out :
  1'd0;
assign cond402_write_en = _guard5547;
assign cond402_clk = clk;
assign cond402_reset = reset;
assign cond402_in =
  _guard5548 ? idx_between_25_41_reg_out :
  1'd0;
assign cond407_write_en = _guard5549;
assign cond407_clk = clk;
assign cond407_reset = reset;
assign cond407_in =
  _guard5550 ? idx_between_11_27_reg_out :
  1'd0;
assign cond410_write_en = _guard5551;
assign cond410_clk = clk;
assign cond410_reset = reset;
assign cond410_in =
  _guard5552 ? idx_between_8_24_reg_out :
  1'd0;
assign cond_wire410_in =
  _guard5555 ? cond410_out :
  _guard5556 ? idx_between_8_24_reg_out :
  1'd0;
assign cond424_write_en = _guard5557;
assign cond424_clk = clk;
assign cond424_reset = reset;
assign cond424_in =
  _guard5558 ? idx_between_31_32_reg_out :
  1'd0;
assign cond432_write_en = _guard5559;
assign cond432_clk = clk;
assign cond432_reset = reset;
assign cond432_in =
  _guard5560 ? idx_between_33_34_reg_out :
  1'd0;
assign cond_wire441_in =
  _guard5561 ? idx_between_16_20_reg_out :
  _guard5564 ? cond441_out :
  1'd0;
assign cond_wire447_in =
  _guard5565 ? idx_between_21_37_reg_out :
  _guard5568 ? cond447_out :
  1'd0;
assign cond458_write_en = _guard5569;
assign cond458_clk = clk;
assign cond458_reset = reset;
assign cond458_in =
  _guard5570 ? idx_between_20_36_reg_out :
  1'd0;
assign cond460_write_en = _guard5571;
assign cond460_clk = clk;
assign cond460_reset = reset;
assign cond460_in =
  _guard5572 ? idx_between_40_41_reg_out :
  1'd0;
assign cond_wire464_in =
  _guard5575 ? cond464_out :
  _guard5576 ? idx_between_41_42_reg_out :
  1'd0;
assign cond_wire469_in =
  _guard5577 ? idx_between_7_23_reg_out :
  _guard5580 ? cond469_out :
  1'd0;
assign cond_wire481_in =
  _guard5583 ? cond481_out :
  _guard5584 ? idx_between_30_31_reg_out :
  1'd0;
assign cond489_write_en = _guard5585;
assign cond489_clk = clk;
assign cond489_reset = reset;
assign cond489_in =
  _guard5586 ? idx_between_32_33_reg_out :
  1'd0;
assign cond_wire489_in =
  _guard5589 ? cond489_out :
  _guard5590 ? idx_between_32_33_reg_out :
  1'd0;
assign cond_wire490_in =
  _guard5591 ? idx_between_13_17_reg_out :
  _guard5594 ? cond490_out :
  1'd0;
assign cond503_write_en = _guard5595;
assign cond503_clk = clk;
assign cond503_reset = reset;
assign cond503_in =
  _guard5596 ? idx_between_16_32_reg_out :
  1'd0;
assign cond504_write_en = _guard5597;
assign cond504_clk = clk;
assign cond504_reset = reset;
assign cond504_in =
  _guard5598 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire510_in =
  _guard5601 ? cond510_out :
  _guard5602 ? idx_between_18_22_reg_out :
  1'd0;
assign cond_wire511_in =
  _guard5603 ? idx_between_18_34_reg_out :
  _guard5606 ? cond511_out :
  1'd0;
assign cond_wire525_in =
  _guard5609 ? cond525_out :
  _guard5610 ? idx_between_41_42_reg_out :
  1'd0;
assign cond539_write_en = _guard5611;
assign cond539_clk = clk;
assign cond539_reset = reset;
assign cond539_in =
  _guard5612 ? idx_between_10_14_reg_out :
  1'd0;
assign cond_wire543_in =
  _guard5615 ? cond543_out :
  _guard5616 ? idx_between_11_15_reg_out :
  1'd0;
assign cond_wire568_in =
  _guard5617 ? idx_between_17_33_reg_out :
  _guard5620 ? cond568_out :
  1'd0;
assign cond576_write_en = _guard5621;
assign cond576_clk = clk;
assign cond576_reset = reset;
assign cond576_in =
  _guard5622 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire577_in =
  _guard5623 ? idx_between_23_39_reg_out :
  _guard5626 ? cond577_out :
  1'd0;
assign cond587_write_en = _guard5627;
assign cond587_clk = clk;
assign cond587_reset = reset;
assign cond587_in =
  _guard5628 ? idx_between_22_26_reg_out :
  1'd0;
assign cond_wire596_in =
  _guard5631 ? cond596_out :
  _guard5632 ? idx_between_24_40_reg_out :
  1'd0;
assign cond601_write_en = _guard5633;
assign cond601_clk = clk;
assign cond601_reset = reset;
assign cond601_in =
  _guard5634 ? idx_between_10_26_reg_out :
  1'd0;
assign cond615_write_en = _guard5635;
assign cond615_clk = clk;
assign cond615_reset = reset;
assign cond615_in =
  _guard5636 ? idx_between_33_34_reg_out :
  1'd0;
assign cond621_write_en = _guard5637;
assign cond621_clk = clk;
assign cond621_reset = reset;
assign cond621_in =
  _guard5638 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire622_in =
  _guard5641 ? cond622_out :
  _guard5642 ? idx_between_19_35_reg_out :
  1'd0;
assign cond637_write_en = _guard5643;
assign cond637_clk = clk;
assign cond637_reset = reset;
assign cond637_in =
  _guard5644 ? idx_between_19_35_reg_out :
  1'd0;
assign cond642_write_en = _guard5645;
assign cond642_clk = clk;
assign cond642_reset = reset;
assign cond642_in =
  _guard5646 ? idx_between_24_40_reg_out :
  1'd0;
assign cond_wire644_in =
  _guard5647 ? idx_between_21_25_reg_out :
  _guard5650 ? cond644_out :
  1'd0;
assign cond_wire653_in =
  _guard5651 ? idx_between_23_39_reg_out :
  _guard5654 ? cond653_out :
  1'd0;
assign cond656_write_en = _guard5655;
assign cond656_clk = clk;
assign cond656_reset = reset;
assign cond656_in =
  _guard5656 ? idx_between_24_28_reg_out :
  1'd0;
assign cond659_write_en = _guard5657;
assign cond659_clk = clk;
assign cond659_reset = reset;
assign cond659_in =
  _guard5658 ? idx_between_44_45_reg_out :
  1'd0;
assign cond679_write_en = _guard5659;
assign cond679_clk = clk;
assign cond679_reset = reset;
assign cond679_in =
  _guard5660 ? idx_between_18_34_reg_out :
  1'd0;
assign cond_wire688_in =
  _guard5661 ? idx_between_36_37_reg_out :
  _guard5664 ? cond688_out :
  1'd0;
assign cond_wire689_in =
  _guard5665 ? idx_between_17_21_reg_out :
  _guard5668 ? cond689_out :
  1'd0;
assign cond_wire711_in =
  _guard5669 ? idx_between_26_42_reg_out :
  _guard5672 ? cond711_out :
  1'd0;
assign cond_wire714_in =
  _guard5673 ? idx_between_23_39_reg_out :
  _guard5676 ? cond714_out :
  1'd0;
assign cond715_write_en = _guard5677;
assign cond715_clk = clk;
assign cond715_reset = reset;
assign cond715_in =
  _guard5678 ? idx_between_27_43_reg_out :
  1'd0;
assign cond718_write_en = _guard5679;
assign cond718_clk = clk;
assign cond718_reset = reset;
assign cond718_in =
  _guard5680 ? idx_between_24_40_reg_out :
  1'd0;
assign cond722_write_en = _guard5681;
assign cond722_clk = clk;
assign cond722_reset = reset;
assign cond722_in =
  _guard5682 ? idx_between_25_41_reg_out :
  1'd0;
assign cond725_write_en = _guard5683;
assign cond725_clk = clk;
assign cond725_reset = reset;
assign cond725_in =
  _guard5684 ? idx_between_26_30_reg_out :
  1'd0;
assign cond_wire743_in =
  _guard5687 ? cond743_out :
  _guard5688 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire745_in =
  _guard5691 ? cond745_out :
  _guard5692 ? idx_between_35_36_reg_out :
  1'd0;
assign cond_wire749_in =
  _guard5693 ? idx_between_36_37_reg_out :
  _guard5696 ? cond749_out :
  1'd0;
assign cond753_write_en = _guard5697;
assign cond753_clk = clk;
assign cond753_reset = reset;
assign cond753_in =
  _guard5698 ? idx_between_37_38_reg_out :
  1'd0;
assign cond765_write_en = _guard5699;
assign cond765_clk = clk;
assign cond765_reset = reset;
assign cond765_in =
  _guard5700 ? idx_between_40_41_reg_out :
  1'd0;
assign cond777_write_en = _guard5701;
assign cond777_clk = clk;
assign cond777_reset = reset;
assign cond777_in =
  _guard5702 ? idx_between_43_44_reg_out :
  1'd0;
assign cond780_write_en = _guard5703;
assign cond780_clk = clk;
assign cond780_reset = reset;
assign cond780_in =
  _guard5704 ? idx_between_28_44_reg_out :
  1'd0;
assign cond781_write_en = _guard5705;
assign cond781_clk = clk;
assign cond781_reset = reset;
assign cond781_in =
  _guard5706 ? idx_between_44_45_reg_out :
  1'd0;
assign cond782_write_en = _guard5707;
assign cond782_clk = clk;
assign cond782_reset = reset;
assign cond782_in =
  _guard5708 ? idx_between_25_29_reg_out :
  1'd0;
assign cond784_write_en = _guard5709;
assign cond784_clk = clk;
assign cond784_reset = reset;
assign cond784_in =
  _guard5710 ? idx_between_29_45_reg_out :
  1'd0;
assign cond_wire785_in =
  _guard5713 ? cond785_out :
  _guard5714 ? idx_between_45_46_reg_out :
  1'd0;
assign cond787_write_en = _guard5715;
assign cond787_clk = clk;
assign cond787_reset = reset;
assign cond787_in =
  _guard5716 ? idx_between_26_42_reg_out :
  1'd0;
assign cond_wire791_in =
  _guard5719 ? cond791_out :
  _guard5720 ? idx_between_27_43_reg_out :
  1'd0;
assign cond795_write_en = _guard5721;
assign cond795_clk = clk;
assign cond795_reset = reset;
assign cond795_in =
  _guard5722 ? idx_between_13_17_reg_out :
  1'd0;
assign cond_wire798_in =
  _guard5725 ? cond798_out :
  _guard5726 ? idx_between_33_34_reg_out :
  1'd0;
assign cond820_write_en = _guard5727;
assign cond820_clk = clk;
assign cond820_reset = reset;
assign cond820_in =
  _guard5728 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire821_in =
  _guard5729 ? idx_between_23_39_reg_out :
  _guard5732 ? cond821_out :
  1'd0;
assign cond834_write_en = _guard5733;
assign cond834_clk = clk;
assign cond834_reset = reset;
assign cond834_in =
  _guard5734 ? idx_between_42_43_reg_out :
  1'd0;
assign cond837_write_en = _guard5735;
assign cond837_clk = clk;
assign cond837_reset = reset;
assign cond837_in =
  _guard5736 ? idx_between_27_43_reg_out :
  1'd0;
assign cond_wire838_in =
  _guard5737 ? idx_between_43_44_reg_out :
  _guard5740 ? cond838_out :
  1'd0;
assign cond_wire852_in =
  _guard5743 ? cond852_out :
  _guard5744 ? idx_between_27_43_reg_out :
  1'd0;
assign cond_wire877_in =
  _guard5745 ? idx_between_18_34_reg_out :
  _guard5748 ? cond877_out :
  1'd0;
assign cond_wire883_in =
  _guard5749 ? idx_between_39_40_reg_out :
  _guard5752 ? cond883_out :
  1'd0;
assign cond888_write_en = _guard5753;
assign cond888_clk = clk;
assign cond888_reset = reset;
assign cond888_in =
  _guard5754 ? idx_between_21_25_reg_out :
  1'd0;
assign cond_wire891_in =
  _guard5757 ? cond891_out :
  _guard5758 ? idx_between_41_42_reg_out :
  1'd0;
assign cond_wire892_in =
  _guard5761 ? cond892_out :
  _guard5762 ? idx_between_22_26_reg_out :
  1'd0;
assign cond_wire893_in =
  _guard5765 ? cond893_out :
  _guard5766 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire900_in =
  _guard5767 ? idx_between_24_28_reg_out :
  _guard5770 ? cond900_out :
  1'd0;
assign cond921_write_en = _guard5771;
assign cond921_clk = clk;
assign cond921_reset = reset;
assign cond921_in =
  _guard5772 ? idx_between_29_45_reg_out :
  1'd0;
assign cond924_write_en = _guard5773;
assign cond924_clk = clk;
assign cond924_reset = reset;
assign cond924_in =
  _guard5774 ? idx_between_14_30_reg_out :
  1'd0;
assign cond927_write_en = _guard5775;
assign cond927_clk = clk;
assign cond927_reset = reset;
assign cond927_in =
  _guard5776 ? idx_between_19_35_reg_out :
  1'd0;
assign cond949_write_en = _guard5777;
assign cond949_clk = clk;
assign cond949_reset = reset;
assign cond949_in =
  _guard5778 ? idx_between_21_25_reg_out :
  1'd0;
assign cond_wire962_in =
  _guard5781 ? cond962_out :
  _guard5782 ? idx_between_24_40_reg_out :
  1'd0;
assign cond968_write_en = _guard5783;
assign cond968_clk = clk;
assign cond968_reset = reset;
assign cond968_in =
  _guard5784 ? idx_between_45_46_reg_out :
  1'd0;
assign cond_wire969_in =
  _guard5785 ? idx_between_26_30_reg_out :
  _guard5788 ? cond969_out :
  1'd0;
assign cond_wire970_in =
  _guard5791 ? cond970_out :
  _guard5792 ? idx_between_26_42_reg_out :
  1'd0;
assign cond979_write_en = _guard5793;
assign cond979_clk = clk;
assign cond979_reset = reset;
assign cond979_in =
  _guard5794 ? idx_between_32_48_reg_out :
  1'd0;
assign cond_wire980_in =
  _guard5795 ? idx_between_48_49_reg_out :
  _guard5798 ? cond980_out :
  1'd0;
assign cond1001_write_en = _guard5799;
assign cond1001_clk = clk;
assign cond1001_reset = reset;
assign cond1001_in =
  _guard5800 ? idx_between_38_39_reg_out :
  1'd0;
assign cond_wire1001_in =
  _guard5803 ? cond1001_out :
  _guard5804 ? idx_between_38_39_reg_out :
  1'd0;
assign cond1006_write_en = _guard5805;
assign cond1006_clk = clk;
assign cond1006_reset = reset;
assign cond1006_in =
  _guard5806 ? idx_between_20_24_reg_out :
  1'd0;
assign cond_wire1008_in =
  _guard5809 ? cond1008_out :
  _guard5810 ? idx_between_24_40_reg_out :
  1'd0;
assign cond_wire1021_in =
  _guard5811 ? idx_between_43_44_reg_out :
  _guard5814 ? cond1021_out :
  1'd0;
assign cond1022_write_en = _guard5815;
assign cond1022_clk = clk;
assign cond1022_reset = reset;
assign cond1022_in =
  _guard5816 ? idx_between_24_28_reg_out :
  1'd0;
assign cond1032_write_en = _guard5817;
assign cond1032_clk = clk;
assign cond1032_reset = reset;
assign cond1032_in =
  _guard5818 ? idx_between_30_46_reg_out :
  1'd0;
assign cond1047_write_en = _guard5819;
assign cond1047_clk = clk;
assign cond1047_reset = reset;
assign cond1047_in =
  _guard5820 ? idx_between_30_46_reg_out :
  1'd0;
assign cond1049_write_en = _guard5821;
assign cond1049_clk = clk;
assign cond1049_reset = reset;
assign cond1049_in =
  _guard5822 ? idx_between_50_51_reg_out :
  1'd0;
assign fsm_write_en = _guard5823;
assign fsm_clk = clk;
assign fsm_reset = reset;
assign fsm_in =
  _guard5826 ? 1'd0 :
  _guard5829 ? adder0_out :
  1'd0;
assign adder_left =
  _guard5830 ? fsm0_out :
  6'd0;
assign adder_right =
  _guard5831 ? 6'd1 :
  6'd0;
assign early_reset_static_par0_go_in = _guard5836;
assign top_0_6_write_en = _guard5839;
assign top_0_6_clk = clk;
assign top_0_6_reset = reset;
assign top_0_6_in = t6_read_data;
assign top_0_15_write_en = _guard5845;
assign top_0_15_clk = clk;
assign top_0_15_reset = reset;
assign top_0_15_in = t15_read_data;
assign left_1_4_write_en = _guard5851;
assign left_1_4_clk = clk;
assign left_1_4_reset = reset;
assign left_1_4_in = left_1_3_out;
assign top_1_5_write_en = _guard5857;
assign top_1_5_clk = clk;
assign top_1_5_reset = reset;
assign top_1_5_in = top_0_5_out;
assign left_1_5_write_en = _guard5863;
assign left_1_5_clk = clk;
assign left_1_5_reset = reset;
assign left_1_5_in = left_1_4_out;
assign left_1_9_write_en = _guard5869;
assign left_1_9_clk = clk;
assign left_1_9_reset = reset;
assign left_1_9_in = left_1_8_out;
assign pe_2_14_mul_ready =
  _guard5875 ? 1'd1 :
  _guard5878 ? 1'd0 :
  1'd0;
assign pe_2_14_clk = clk;
assign pe_2_14_top =
  _guard5891 ? top_2_14_out :
  32'd0;
assign pe_2_14_left =
  _guard5904 ? left_2_14_out :
  32'd0;
assign pe_2_14_reset = reset;
assign pe_2_14_go = _guard5917;
assign left_2_15_write_en = _guard5920;
assign left_2_15_clk = clk;
assign left_2_15_reset = reset;
assign left_2_15_in = left_2_14_out;
assign pe_3_4_mul_ready =
  _guard5926 ? 1'd1 :
  _guard5929 ? 1'd0 :
  1'd0;
assign pe_3_4_clk = clk;
assign pe_3_4_top =
  _guard5942 ? top_3_4_out :
  32'd0;
assign pe_3_4_left =
  _guard5955 ? left_3_4_out :
  32'd0;
assign pe_3_4_reset = reset;
assign pe_3_4_go = _guard5968;
assign pe_3_7_mul_ready =
  _guard5971 ? 1'd1 :
  _guard5974 ? 1'd0 :
  1'd0;
assign pe_3_7_clk = clk;
assign pe_3_7_top =
  _guard5987 ? top_3_7_out :
  32'd0;
assign pe_3_7_left =
  _guard6000 ? left_3_7_out :
  32'd0;
assign pe_3_7_reset = reset;
assign pe_3_7_go = _guard6013;
assign top_3_8_write_en = _guard6016;
assign top_3_8_clk = clk;
assign top_3_8_reset = reset;
assign top_3_8_in = top_2_8_out;
assign left_3_9_write_en = _guard6022;
assign left_3_9_clk = clk;
assign left_3_9_reset = reset;
assign left_3_9_in = left_3_8_out;
assign top_3_11_write_en = _guard6028;
assign top_3_11_clk = clk;
assign top_3_11_reset = reset;
assign top_3_11_in = top_2_11_out;
assign left_3_12_write_en = _guard6034;
assign left_3_12_clk = clk;
assign left_3_12_reset = reset;
assign left_3_12_in = left_3_11_out;
assign pe_4_0_mul_ready =
  _guard6040 ? 1'd1 :
  _guard6043 ? 1'd0 :
  1'd0;
assign pe_4_0_clk = clk;
assign pe_4_0_top =
  _guard6056 ? top_4_0_out :
  32'd0;
assign pe_4_0_left =
  _guard6069 ? left_4_0_out :
  32'd0;
assign pe_4_0_reset = reset;
assign pe_4_0_go = _guard6082;
assign left_4_2_write_en = _guard6085;
assign left_4_2_clk = clk;
assign left_4_2_reset = reset;
assign left_4_2_in = left_4_1_out;
assign pe_5_0_mul_ready =
  _guard6091 ? 1'd1 :
  _guard6094 ? 1'd0 :
  1'd0;
assign pe_5_0_clk = clk;
assign pe_5_0_top =
  _guard6107 ? top_5_0_out :
  32'd0;
assign pe_5_0_left =
  _guard6120 ? left_5_0_out :
  32'd0;
assign pe_5_0_reset = reset;
assign pe_5_0_go = _guard6133;
assign left_5_6_write_en = _guard6136;
assign left_5_6_clk = clk;
assign left_5_6_reset = reset;
assign left_5_6_in = left_5_5_out;
assign top_5_15_write_en = _guard6142;
assign top_5_15_clk = clk;
assign top_5_15_reset = reset;
assign top_5_15_in = top_4_15_out;
assign left_6_5_write_en = _guard6148;
assign left_6_5_clk = clk;
assign left_6_5_reset = reset;
assign left_6_5_in = left_6_4_out;
assign top_6_6_write_en = _guard6154;
assign top_6_6_clk = clk;
assign top_6_6_reset = reset;
assign top_6_6_in = top_5_6_out;
assign pe_6_11_mul_ready =
  _guard6160 ? 1'd1 :
  _guard6163 ? 1'd0 :
  1'd0;
assign pe_6_11_clk = clk;
assign pe_6_11_top =
  _guard6176 ? top_6_11_out :
  32'd0;
assign pe_6_11_left =
  _guard6189 ? left_6_11_out :
  32'd0;
assign pe_6_11_reset = reset;
assign pe_6_11_go = _guard6202;
assign left_7_12_write_en = _guard6205;
assign left_7_12_clk = clk;
assign left_7_12_reset = reset;
assign left_7_12_in = left_7_11_out;
assign pe_7_15_mul_ready =
  _guard6211 ? 1'd1 :
  _guard6214 ? 1'd0 :
  1'd0;
assign pe_7_15_clk = clk;
assign pe_7_15_top =
  _guard6227 ? top_7_15_out :
  32'd0;
assign pe_7_15_left =
  _guard6240 ? left_7_15_out :
  32'd0;
assign pe_7_15_reset = reset;
assign pe_7_15_go = _guard6253;
assign top_8_7_write_en = _guard6256;
assign top_8_7_clk = clk;
assign top_8_7_reset = reset;
assign top_8_7_in = top_7_7_out;
assign left_8_10_write_en = _guard6262;
assign left_8_10_clk = clk;
assign left_8_10_reset = reset;
assign left_8_10_in = left_8_9_out;
assign pe_9_7_mul_ready =
  _guard6268 ? 1'd1 :
  _guard6271 ? 1'd0 :
  1'd0;
assign pe_9_7_clk = clk;
assign pe_9_7_top =
  _guard6284 ? top_9_7_out :
  32'd0;
assign pe_9_7_left =
  _guard6297 ? left_9_7_out :
  32'd0;
assign pe_9_7_reset = reset;
assign pe_9_7_go = _guard6310;
assign left_10_6_write_en = _guard6313;
assign left_10_6_clk = clk;
assign left_10_6_reset = reset;
assign left_10_6_in = left_10_5_out;
assign pe_11_8_mul_ready =
  _guard6319 ? 1'd1 :
  _guard6322 ? 1'd0 :
  1'd0;
assign pe_11_8_clk = clk;
assign pe_11_8_top =
  _guard6335 ? top_11_8_out :
  32'd0;
assign pe_11_8_left =
  _guard6348 ? left_11_8_out :
  32'd0;
assign pe_11_8_reset = reset;
assign pe_11_8_go = _guard6361;
assign top_11_11_write_en = _guard6364;
assign top_11_11_clk = clk;
assign top_11_11_reset = reset;
assign top_11_11_in = top_10_11_out;
assign pe_11_15_mul_ready =
  _guard6370 ? 1'd1 :
  _guard6373 ? 1'd0 :
  1'd0;
assign pe_11_15_clk = clk;
assign pe_11_15_top =
  _guard6386 ? top_11_15_out :
  32'd0;
assign pe_11_15_left =
  _guard6399 ? left_11_15_out :
  32'd0;
assign pe_11_15_reset = reset;
assign pe_11_15_go = _guard6412;
assign left_12_5_write_en = _guard6415;
assign left_12_5_clk = clk;
assign left_12_5_reset = reset;
assign left_12_5_in = left_12_4_out;
assign pe_12_9_mul_ready =
  _guard6421 ? 1'd1 :
  _guard6424 ? 1'd0 :
  1'd0;
assign pe_12_9_clk = clk;
assign pe_12_9_top =
  _guard6437 ? top_12_9_out :
  32'd0;
assign pe_12_9_left =
  _guard6450 ? left_12_9_out :
  32'd0;
assign pe_12_9_reset = reset;
assign pe_12_9_go = _guard6463;
assign pe_12_12_mul_ready =
  _guard6466 ? 1'd1 :
  _guard6469 ? 1'd0 :
  1'd0;
assign pe_12_12_clk = clk;
assign pe_12_12_top =
  _guard6482 ? top_12_12_out :
  32'd0;
assign pe_12_12_left =
  _guard6495 ? left_12_12_out :
  32'd0;
assign pe_12_12_reset = reset;
assign pe_12_12_go = _guard6508;
assign top_12_14_write_en = _guard6511;
assign top_12_14_clk = clk;
assign top_12_14_reset = reset;
assign top_12_14_in = top_11_14_out;
assign top_13_0_write_en = _guard6517;
assign top_13_0_clk = clk;
assign top_13_0_reset = reset;
assign top_13_0_in = top_12_0_out;
assign top_13_10_write_en = _guard6523;
assign top_13_10_clk = clk;
assign top_13_10_reset = reset;
assign top_13_10_in = top_12_10_out;
assign left_14_8_write_en = _guard6529;
assign left_14_8_clk = clk;
assign left_14_8_reset = reset;
assign left_14_8_in = left_14_7_out;
assign top_14_12_write_en = _guard6535;
assign top_14_12_clk = clk;
assign top_14_12_reset = reset;
assign top_14_12_in = top_13_12_out;
assign pe_14_13_mul_ready =
  _guard6541 ? 1'd1 :
  _guard6544 ? 1'd0 :
  1'd0;
assign pe_14_13_clk = clk;
assign pe_14_13_top =
  _guard6557 ? top_14_13_out :
  32'd0;
assign pe_14_13_left =
  _guard6570 ? left_14_13_out :
  32'd0;
assign pe_14_13_reset = reset;
assign pe_14_13_go = _guard6583;
assign top_14_14_write_en = _guard6586;
assign top_14_14_clk = clk;
assign top_14_14_reset = reset;
assign top_14_14_in = top_13_14_out;
assign pe_15_2_mul_ready =
  _guard6592 ? 1'd1 :
  _guard6595 ? 1'd0 :
  1'd0;
assign pe_15_2_clk = clk;
assign pe_15_2_top =
  _guard6608 ? top_15_2_out :
  32'd0;
assign pe_15_2_left =
  _guard6621 ? left_15_2_out :
  32'd0;
assign pe_15_2_reset = reset;
assign pe_15_2_go = _guard6634;
assign top_15_12_write_en = _guard6637;
assign top_15_12_clk = clk;
assign top_15_12_reset = reset;
assign top_15_12_in = top_14_12_out;
assign l0_idx_write_en = _guard6647;
assign l0_idx_clk = clk;
assign l0_idx_reset = reset;
assign l0_idx_in =
  _guard6650 ? 5'd0 :
  _guard6653 ? l0_add_out :
  'x;
assign l11_idx_write_en = _guard6660;
assign l11_idx_clk = clk;
assign l11_idx_reset = reset;
assign l11_idx_in =
  _guard6663 ? 5'd0 :
  _guard6666 ? l11_add_out :
  'x;
assign idx_between_16_20_reg_write_en = _guard6671;
assign idx_between_16_20_reg_clk = clk;
assign idx_between_16_20_reg_reset = reset;
assign idx_between_16_20_reg_in =
  _guard6672 ? idx_between_16_20_comb_out :
  _guard6675 ? 1'd0 :
  'x;
assign idx_between_44_45_reg_write_en = _guard6680;
assign idx_between_44_45_reg_clk = clk;
assign idx_between_44_45_reg_reset = reset;
assign idx_between_44_45_reg_in =
  _guard6683 ? 1'd0 :
  _guard6684 ? idx_between_44_45_comb_out :
  'x;
assign idx_between_31_47_comb_left = index_ge_31_out;
assign idx_between_31_47_comb_right = index_lt_47_out;
assign index_ge_24_left = idx_add_out;
assign index_ge_24_right = 6'd24;
assign index_lt_50_left = idx_add_out;
assign index_lt_50_right = 6'd50;
assign index_ge_50_left = idx_add_out;
assign index_ge_50_right = 6'd50;
assign idx_between_46_47_comb_left = index_ge_46_out;
assign idx_between_46_47_comb_right = index_lt_47_out;
assign idx_between_23_24_reg_write_en = _guard6699;
assign idx_between_23_24_reg_clk = clk;
assign idx_between_23_24_reg_reset = reset;
assign idx_between_23_24_reg_in =
  _guard6700 ? idx_between_23_24_comb_out :
  _guard6703 ? 1'd0 :
  'x;
assign idx_between_28_32_reg_write_en = _guard6708;
assign idx_between_28_32_reg_clk = clk;
assign idx_between_28_32_reg_reset = reset;
assign idx_between_28_32_reg_in =
  _guard6709 ? idx_between_28_32_comb_out :
  _guard6712 ? 1'd0 :
  'x;
assign idx_between_10_26_comb_left = index_ge_10_out;
assign idx_between_10_26_comb_right = index_lt_26_out;
assign idx_between_29_33_comb_left = index_ge_29_out;
assign idx_between_29_33_comb_right = index_lt_33_out;
assign idx_between_7_11_reg_write_en = _guard6721;
assign idx_between_7_11_reg_clk = clk;
assign idx_between_7_11_reg_reset = reset;
assign idx_between_7_11_reg_in =
  _guard6724 ? 1'd0 :
  _guard6725 ? idx_between_7_11_comb_out :
  'x;
assign index_lt_11_left = idx_add_out;
assign index_lt_11_right = 6'd11;
assign idx_between_37_38_comb_left = index_ge_37_out;
assign idx_between_37_38_comb_right = index_lt_38_out;
assign index_ge_39_left = idx_add_out;
assign index_ge_39_right = 6'd39;
assign idx_between_2_18_reg_write_en = _guard6736;
assign idx_between_2_18_reg_clk = clk;
assign idx_between_2_18_reg_reset = reset;
assign idx_between_2_18_reg_in =
  _guard6737 ? idx_between_2_18_comb_out :
  _guard6740 ? 1'd0 :
  'x;
assign cond11_write_en = _guard6741;
assign cond11_clk = clk;
assign cond11_reset = reset;
assign cond11_in =
  _guard6742 ? idx_between_3_19_reg_out :
  1'd0;
assign cond15_write_en = _guard6743;
assign cond15_clk = clk;
assign cond15_reset = reset;
assign cond15_in =
  _guard6744 ? idx_between_4_8_reg_out :
  1'd0;
assign cond_wire27_in =
  _guard6747 ? cond27_out :
  _guard6748 ? idx_between_10_26_reg_out :
  1'd0;
assign cond43_write_en = _guard6749;
assign cond43_clk = clk;
assign cond43_reset = reset;
assign cond43_in =
  _guard6750 ? idx_between_29_30_reg_out :
  1'd0;
assign cond_wire43_in =
  _guard6753 ? cond43_out :
  _guard6754 ? idx_between_29_30_reg_out :
  1'd0;
assign cond_wire44_in =
  _guard6757 ? cond44_out :
  _guard6758 ? idx_between_9_25_reg_out :
  1'd0;
assign cond62_write_en = _guard6759;
assign cond62_clk = clk;
assign cond62_reset = reset;
assign cond62_in =
  _guard6760 ? idx_between_17_33_reg_out :
  1'd0;
assign cond_wire63_in =
  _guard6763 ? cond63_out :
  _guard6764 ? idx_between_33_34_reg_out :
  1'd0;
assign cond_wire67_in =
  _guard6765 ? idx_between_18_34_reg_out :
  _guard6768 ? cond67_out :
  1'd0;
assign cond73_write_en = _guard6769;
assign cond73_clk = clk;
assign cond73_reset = reset;
assign cond73_in =
  _guard6770 ? idx_between_35_36_reg_out :
  1'd0;
assign cond_wire77_in =
  _guard6771 ? idx_between_20_36_reg_out :
  _guard6774 ? cond77_out :
  1'd0;
assign cond103_write_en = _guard6775;
assign cond103_clk = clk;
assign cond103_reset = reset;
assign cond103_in =
  _guard6776 ? idx_between_27_28_reg_out :
  1'd0;
assign cond114_write_en = _guard6777;
assign cond114_clk = clk;
assign cond114_reset = reset;
assign cond114_in =
  _guard6778 ? idx_between_14_30_reg_out :
  1'd0;
assign cond118_write_en = _guard6779;
assign cond118_clk = clk;
assign cond118_reset = reset;
assign cond118_in =
  _guard6780 ? idx_between_15_31_reg_out :
  1'd0;
assign cond121_write_en = _guard6781;
assign cond121_clk = clk;
assign cond121_reset = reset;
assign cond121_in =
  _guard6782 ? idx_between_12_28_reg_out :
  1'd0;
assign cond123_write_en = _guard6783;
assign cond123_clk = clk;
assign cond123_reset = reset;
assign cond123_in =
  _guard6784 ? idx_between_32_33_reg_out :
  1'd0;
assign cond_wire126_in =
  _guard6785 ? idx_between_17_33_reg_out :
  _guard6788 ? cond126_out :
  1'd0;
assign cond_wire154_in =
  _guard6789 ? idx_between_5_21_reg_out :
  _guard6792 ? cond154_out :
  1'd0;
assign cond_wire195_in =
  _guard6795 ? cond195_out :
  _guard6796 ? idx_between_19_35_reg_out :
  1'd0;
assign cond206_write_en = _guard6797;
assign cond206_clk = clk;
assign cond206_reset = reset;
assign cond206_in =
  _guard6798 ? idx_between_18_34_reg_out :
  1'd0;
assign cond216_write_en = _guard6799;
assign cond216_clk = clk;
assign cond216_reset = reset;
assign cond216_in =
  _guard6800 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire218_in =
  _guard6801 ? idx_between_6_10_reg_out :
  _guard6804 ? cond218_out :
  1'd0;
assign cond_wire238_in =
  _guard6807 ? cond238_out :
  _guard6808 ? idx_between_11_15_reg_out :
  1'd0;
assign cond240_write_en = _guard6809;
assign cond240_clk = clk;
assign cond240_reset = reset;
assign cond240_in =
  _guard6810 ? idx_between_15_31_reg_out :
  1'd0;
assign cond251_write_en = _guard6811;
assign cond251_clk = clk;
assign cond251_reset = reset;
assign cond251_in =
  _guard6812 ? idx_between_14_30_reg_out :
  1'd0;
assign cond264_write_en = _guard6813;
assign cond264_clk = clk;
assign cond264_reset = reset;
assign cond264_in =
  _guard6814 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire265_in =
  _guard6817 ? cond265_out :
  _guard6818 ? idx_between_37_38_reg_out :
  1'd0;
assign cond271_write_en = _guard6819;
assign cond271_clk = clk;
assign cond271_reset = reset;
assign cond271_in =
  _guard6820 ? idx_between_19_35_reg_out :
  1'd0;
assign cond279_write_en = _guard6821;
assign cond279_clk = clk;
assign cond279_reset = reset;
assign cond279_in =
  _guard6822 ? idx_between_6_10_reg_out :
  1'd0;
assign cond_wire279_in =
  _guard6823 ? idx_between_6_10_reg_out :
  _guard6826 ? cond279_out :
  1'd0;
assign cond_wire290_in =
  _guard6829 ? cond290_out :
  _guard6830 ? idx_between_28_29_reg_out :
  1'd0;
assign cond_wire298_in =
  _guard6831 ? idx_between_30_31_reg_out :
  _guard6834 ? cond298_out :
  1'd0;
assign cond300_write_en = _guard6835;
assign cond300_clk = clk;
assign cond300_reset = reset;
assign cond300_in =
  _guard6836 ? idx_between_11_27_reg_out :
  1'd0;
assign cond_wire301_in =
  _guard6839 ? cond301_out :
  _guard6840 ? idx_between_15_31_reg_out :
  1'd0;
assign cond305_write_en = _guard6841;
assign cond305_clk = clk;
assign cond305_reset = reset;
assign cond305_in =
  _guard6842 ? idx_between_16_32_reg_out :
  1'd0;
assign cond313_write_en = _guard6843;
assign cond313_clk = clk;
assign cond313_reset = reset;
assign cond313_in =
  _guard6844 ? idx_between_18_34_reg_out :
  1'd0;
assign cond315_write_en = _guard6845;
assign cond315_clk = clk;
assign cond315_reset = reset;
assign cond315_in =
  _guard6846 ? idx_between_15_19_reg_out :
  1'd0;
assign cond324_write_en = _guard6847;
assign cond324_clk = clk;
assign cond324_reset = reset;
assign cond324_in =
  _guard6848 ? idx_between_17_33_reg_out :
  1'd0;
assign cond_wire339_in =
  _guard6849 ? idx_between_5_21_reg_out :
  _guard6852 ? cond339_out :
  1'd0;
assign cond_wire342_in =
  _guard6855 ? cond342_out :
  _guard6856 ? idx_between_10_26_reg_out :
  1'd0;
assign cond343_write_en = _guard6857;
assign cond343_clk = clk;
assign cond343_reset = reset;
assign cond343_in =
  _guard6858 ? idx_between_26_27_reg_out :
  1'd0;
assign cond_wire351_in =
  _guard6859 ? idx_between_28_29_reg_out :
  _guard6862 ? cond351_out :
  1'd0;
assign cond354_write_en = _guard6863;
assign cond354_clk = clk;
assign cond354_reset = reset;
assign cond354_in =
  _guard6864 ? idx_between_13_29_reg_out :
  1'd0;
assign cond_wire356_in =
  _guard6867 ? cond356_out :
  _guard6868 ? idx_between_10_14_reg_out :
  1'd0;
assign cond362_write_en = _guard6869;
assign cond362_clk = clk;
assign cond362_reset = reset;
assign cond362_in =
  _guard6870 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire362_in =
  _guard6873 ? cond362_out :
  _guard6874 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire364_in =
  _guard6875 ? idx_between_12_16_reg_out :
  _guard6878 ? cond364_out :
  1'd0;
assign cond_wire367_in =
  _guard6881 ? cond367_out :
  _guard6882 ? idx_between_32_33_reg_out :
  1'd0;
assign cond_wire386_in =
  _guard6885 ? cond386_out :
  _guard6886 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire388_in =
  _guard6889 ? cond388_out :
  _guard6890 ? idx_between_18_22_reg_out :
  1'd0;
assign cond390_write_en = _guard6891;
assign cond390_clk = clk;
assign cond390_reset = reset;
assign cond390_in =
  _guard6892 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire390_in =
  _guard6895 ? cond390_out :
  _guard6896 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire402_in =
  _guard6899 ? cond402_out :
  _guard6900 ? idx_between_25_41_reg_out :
  1'd0;
assign cond_wire404_in =
  _guard6901 ? idx_between_6_22_reg_out :
  _guard6904 ? cond404_out :
  1'd0;
assign cond_wire412_in =
  _guard6907 ? cond412_out :
  _guard6908 ? idx_between_28_29_reg_out :
  1'd0;
assign cond_wire419_in =
  _guard6909 ? idx_between_14_30_reg_out :
  _guard6912 ? cond419_out :
  1'd0;
assign cond433_write_en = _guard6913;
assign cond433_clk = clk;
assign cond433_reset = reset;
assign cond433_in =
  _guard6914 ? idx_between_14_18_reg_out :
  1'd0;
assign cond440_write_en = _guard6915;
assign cond440_clk = clk;
assign cond440_reset = reset;
assign cond440_in =
  _guard6916 ? idx_between_35_36_reg_out :
  1'd0;
assign cond445_write_en = _guard6917;
assign cond445_clk = clk;
assign cond445_reset = reset;
assign cond445_in =
  _guard6918 ? idx_between_17_21_reg_out :
  1'd0;
assign cond_wire445_in =
  _guard6921 ? cond445_out :
  _guard6922 ? idx_between_17_21_reg_out :
  1'd0;
assign cond449_write_en = _guard6923;
assign cond449_clk = clk;
assign cond449_reset = reset;
assign cond449_in =
  _guard6924 ? idx_between_18_22_reg_out :
  1'd0;
assign cond_wire456_in =
  _guard6927 ? cond456_out :
  _guard6928 ? idx_between_39_40_reg_out :
  1'd0;
assign cond457_write_en = _guard6929;
assign cond457_clk = clk;
assign cond457_reset = reset;
assign cond457_in =
  _guard6930 ? idx_between_20_24_reg_out :
  1'd0;
assign cond_wire467_in =
  _guard6933 ? cond467_out :
  _guard6934 ? idx_between_26_42_reg_out :
  1'd0;
assign cond473_write_en = _guard6935;
assign cond473_clk = clk;
assign cond473_reset = reset;
assign cond473_in =
  _guard6936 ? idx_between_28_29_reg_out :
  1'd0;
assign cond_wire473_in =
  _guard6939 ? cond473_out :
  _guard6940 ? idx_between_28_29_reg_out :
  1'd0;
assign cond_wire479_in =
  _guard6941 ? idx_between_10_26_reg_out :
  _guard6944 ? cond479_out :
  1'd0;
assign cond_wire491_in =
  _guard6945 ? idx_between_13_29_reg_out :
  _guard6948 ? cond491_out :
  1'd0;
assign cond_wire495_in =
  _guard6951 ? cond495_out :
  _guard6952 ? idx_between_14_30_reg_out :
  1'd0;
assign cond_wire496_in =
  _guard6953 ? idx_between_18_34_reg_out :
  _guard6956 ? cond496_out :
  1'd0;
assign cond498_write_en = _guard6957;
assign cond498_clk = clk;
assign cond498_reset = reset;
assign cond498_in =
  _guard6958 ? idx_between_15_19_reg_out :
  1'd0;
assign cond_wire516_in =
  _guard6959 ? idx_between_23_39_reg_out :
  _guard6962 ? cond516_out :
  1'd0;
assign cond_wire517_in =
  _guard6963 ? idx_between_39_40_reg_out :
  _guard6966 ? cond517_out :
  1'd0;
assign cond520_write_en = _guard6967;
assign cond520_clk = clk;
assign cond520_reset = reset;
assign cond520_in =
  _guard6968 ? idx_between_24_40_reg_out :
  1'd0;
assign cond547_write_en = _guard6969;
assign cond547_clk = clk;
assign cond547_reset = reset;
assign cond547_in =
  _guard6970 ? idx_between_12_16_reg_out :
  1'd0;
assign cond549_write_en = _guard6971;
assign cond549_clk = clk;
assign cond549_reset = reset;
assign cond549_in =
  _guard6972 ? idx_between_16_32_reg_out :
  1'd0;
assign cond572_write_en = _guard6973;
assign cond572_clk = clk;
assign cond572_reset = reset;
assign cond572_in =
  _guard6974 ? idx_between_18_34_reg_out :
  1'd0;
assign cond588_write_en = _guard6975;
assign cond588_clk = clk;
assign cond588_reset = reset;
assign cond588_in =
  _guard6976 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire594_in =
  _guard6977 ? idx_between_43_44_reg_out :
  _guard6980 ? cond594_out :
  1'd0;
assign cond_wire599_in =
  _guard6983 ? cond599_out :
  _guard6984 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire615_in =
  _guard6987 ? cond615_out :
  _guard6988 ? idx_between_33_34_reg_out :
  1'd0;
assign cond_wire641_in =
  _guard6989 ? idx_between_20_36_reg_out :
  _guard6992 ? cond641_out :
  1'd0;
assign cond661_write_en = _guard6993;
assign cond661_clk = clk;
assign cond661_reset = reset;
assign cond661_in =
  _guard6994 ? idx_between_25_41_reg_out :
  1'd0;
assign cond666_write_en = _guard6995;
assign cond666_clk = clk;
assign cond666_reset = reset;
assign cond666_in =
  _guard6996 ? idx_between_11_27_reg_out :
  1'd0;
assign cond670_write_en = _guard6997;
assign cond670_clk = clk;
assign cond670_reset = reset;
assign cond670_in =
  _guard6998 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire678_in =
  _guard6999 ? idx_between_14_30_reg_out :
  _guard7002 ? cond678_out :
  1'd0;
assign cond_wire695_in =
  _guard7005 ? cond695_out :
  _guard7006 ? idx_between_22_38_reg_out :
  1'd0;
assign cond697_write_en = _guard7007;
assign cond697_clk = clk;
assign cond697_reset = reset;
assign cond697_in =
  _guard7008 ? idx_between_19_23_reg_out :
  1'd0;
assign cond704_write_en = _guard7009;
assign cond704_clk = clk;
assign cond704_reset = reset;
assign cond704_in =
  _guard7010 ? idx_between_40_41_reg_out :
  1'd0;
assign cond_wire709_in =
  _guard7013 ? cond709_out :
  _guard7014 ? idx_between_22_26_reg_out :
  1'd0;
assign cond_wire742_in =
  _guard7015 ? idx_between_15_19_reg_out :
  _guard7018 ? cond742_out :
  1'd0;
assign cond_wire756_in =
  _guard7019 ? idx_between_22_38_reg_out :
  _guard7022 ? cond756_out :
  1'd0;
assign cond_wire760_in =
  _guard7025 ? cond760_out :
  _guard7026 ? idx_between_23_39_reg_out :
  1'd0;
assign cond770_write_en = _guard7027;
assign cond770_clk = clk;
assign cond770_reset = reset;
assign cond770_in =
  _guard7028 ? idx_between_22_26_reg_out :
  1'd0;
assign cond789_write_en = _guard7029;
assign cond789_clk = clk;
assign cond789_reset = reset;
assign cond789_in =
  _guard7030 ? idx_between_46_47_reg_out :
  1'd0;
assign cond_wire812_in =
  _guard7031 ? idx_between_17_33_reg_out :
  _guard7034 ? cond812_out :
  1'd0;
assign cond815_write_en = _guard7035;
assign cond815_clk = clk;
assign cond815_reset = reset;
assign cond815_in =
  _guard7036 ? idx_between_18_22_reg_out :
  1'd0;
assign cond819_write_en = _guard7037;
assign cond819_clk = clk;
assign cond819_reset = reset;
assign cond819_in =
  _guard7038 ? idx_between_19_23_reg_out :
  1'd0;
assign cond_wire820_in =
  _guard7041 ? cond820_out :
  _guard7042 ? idx_between_19_35_reg_out :
  1'd0;
assign cond838_write_en = _guard7043;
assign cond838_clk = clk;
assign cond838_reset = reset;
assign cond838_in =
  _guard7044 ? idx_between_43_44_reg_out :
  1'd0;
assign cond839_write_en = _guard7045;
assign cond839_clk = clk;
assign cond839_reset = reset;
assign cond839_in =
  _guard7046 ? idx_between_24_28_reg_out :
  1'd0;
assign cond_wire843_in =
  _guard7047 ? idx_between_25_29_reg_out :
  _guard7050 ? cond843_out :
  1'd0;
assign cond_wire844_in =
  _guard7053 ? cond844_out :
  _guard7054 ? idx_between_25_41_reg_out :
  1'd0;
assign cond_wire862_in =
  _guard7057 ? cond862_out :
  _guard7058 ? idx_between_18_34_reg_out :
  1'd0;
assign cond_wire903_in =
  _guard7059 ? idx_between_44_45_reg_out :
  _guard7062 ? cond903_out :
  1'd0;
assign cond908_write_en = _guard7063;
assign cond908_clk = clk;
assign cond908_reset = reset;
assign cond908_in =
  _guard7064 ? idx_between_26_30_reg_out :
  1'd0;
assign cond_wire922_in =
  _guard7067 ? cond922_out :
  _guard7068 ? idx_between_33_49_reg_out :
  1'd0;
assign cond_wire923_in =
  _guard7071 ? cond923_out :
  _guard7072 ? idx_between_49_50_reg_out :
  1'd0;
assign cond932_write_en = _guard7073;
assign cond932_clk = clk;
assign cond932_reset = reset;
assign cond932_in =
  _guard7074 ? idx_between_36_37_reg_out :
  1'd0;
assign cond950_write_en = _guard7075;
assign cond950_clk = clk;
assign cond950_reset = reset;
assign cond950_in =
  _guard7076 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire954_in =
  _guard7077 ? idx_between_22_38_reg_out :
  _guard7080 ? cond954_out :
  1'd0;
assign cond970_write_en = _guard7081;
assign cond970_clk = clk;
assign cond970_reset = reset;
assign cond970_in =
  _guard7082 ? idx_between_26_42_reg_out :
  1'd0;
assign cond973_write_en = _guard7083;
assign cond973_clk = clk;
assign cond973_reset = reset;
assign cond973_in =
  _guard7084 ? idx_between_27_31_reg_out :
  1'd0;
assign cond976_write_en = _guard7085;
assign cond976_clk = clk;
assign cond976_reset = reset;
assign cond976_in =
  _guard7086 ? idx_between_47_48_reg_out :
  1'd0;
assign cond981_write_en = _guard7087;
assign cond981_clk = clk;
assign cond981_reset = reset;
assign cond981_in =
  _guard7088 ? idx_between_29_33_reg_out :
  1'd0;
assign cond1003_write_en = _guard7089;
assign cond1003_clk = clk;
assign cond1003_reset = reset;
assign cond1003_in =
  _guard7090 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire1007_in =
  _guard7091 ? idx_between_20_36_reg_out :
  _guard7094 ? cond1007_out :
  1'd0;
assign cond_wire1017_in =
  _guard7095 ? idx_between_42_43_reg_out :
  _guard7098 ? cond1017_out :
  1'd0;
assign cond1023_write_en = _guard7099;
assign cond1023_clk = clk;
assign cond1023_reset = reset;
assign cond1023_in =
  _guard7100 ? idx_between_24_40_reg_out :
  1'd0;
assign cond1031_write_en = _guard7101;
assign cond1031_clk = clk;
assign cond1031_reset = reset;
assign cond1031_in =
  _guard7102 ? idx_between_26_42_reg_out :
  1'd0;
assign cond_wire1032_in =
  _guard7103 ? idx_between_30_46_reg_out :
  _guard7106 ? cond1032_out :
  1'd0;
assign cond_wire1035_in =
  _guard7107 ? idx_between_27_43_reg_out :
  _guard7110 ? cond1035_out :
  1'd0;
assign pe_0_1_mul_ready =
  _guard7113 ? 1'd1 :
  _guard7116 ? 1'd0 :
  1'd0;
assign pe_0_1_clk = clk;
assign pe_0_1_top =
  _guard7129 ? top_0_1_out :
  32'd0;
assign pe_0_1_left =
  _guard7142 ? left_0_1_out :
  32'd0;
assign pe_0_1_reset = reset;
assign pe_0_1_go = _guard7155;
assign left_0_6_write_en = _guard7158;
assign left_0_6_clk = clk;
assign left_0_6_reset = reset;
assign left_0_6_in = left_0_5_out;
assign pe_0_7_mul_ready =
  _guard7164 ? 1'd1 :
  _guard7167 ? 1'd0 :
  1'd0;
assign pe_0_7_clk = clk;
assign pe_0_7_top =
  _guard7180 ? top_0_7_out :
  32'd0;
assign pe_0_7_left =
  _guard7193 ? left_0_7_out :
  32'd0;
assign pe_0_7_reset = reset;
assign pe_0_7_go = _guard7206;
assign top_0_11_write_en = _guard7209;
assign top_0_11_clk = clk;
assign top_0_11_reset = reset;
assign top_0_11_in = t11_read_data;
assign left_1_2_write_en = _guard7215;
assign left_1_2_clk = clk;
assign left_1_2_reset = reset;
assign left_1_2_in = left_1_1_out;
assign pe_1_8_mul_ready =
  _guard7221 ? 1'd1 :
  _guard7224 ? 1'd0 :
  1'd0;
assign pe_1_8_clk = clk;
assign pe_1_8_top =
  _guard7237 ? top_1_8_out :
  32'd0;
assign pe_1_8_left =
  _guard7250 ? left_1_8_out :
  32'd0;
assign pe_1_8_reset = reset;
assign pe_1_8_go = _guard7263;
assign top_1_10_write_en = _guard7266;
assign top_1_10_clk = clk;
assign top_1_10_reset = reset;
assign top_1_10_in = top_0_10_out;
assign pe_1_15_mul_ready =
  _guard7272 ? 1'd1 :
  _guard7275 ? 1'd0 :
  1'd0;
assign pe_1_15_clk = clk;
assign pe_1_15_top =
  _guard7288 ? top_1_15_out :
  32'd0;
assign pe_1_15_left =
  _guard7301 ? left_1_15_out :
  32'd0;
assign pe_1_15_reset = reset;
assign pe_1_15_go = _guard7314;
assign left_2_2_write_en = _guard7317;
assign left_2_2_clk = clk;
assign left_2_2_reset = reset;
assign left_2_2_in = left_2_1_out;
assign top_2_5_write_en = _guard7323;
assign top_2_5_clk = clk;
assign top_2_5_reset = reset;
assign top_2_5_in = top_1_5_out;
assign pe_2_7_mul_ready =
  _guard7329 ? 1'd1 :
  _guard7332 ? 1'd0 :
  1'd0;
assign pe_2_7_clk = clk;
assign pe_2_7_top =
  _guard7345 ? top_2_7_out :
  32'd0;
assign pe_2_7_left =
  _guard7358 ? left_2_7_out :
  32'd0;
assign pe_2_7_reset = reset;
assign pe_2_7_go = _guard7371;
assign left_2_7_write_en = _guard7374;
assign left_2_7_clk = clk;
assign left_2_7_reset = reset;
assign left_2_7_in = left_2_6_out;
assign pe_2_13_mul_ready =
  _guard7380 ? 1'd1 :
  _guard7383 ? 1'd0 :
  1'd0;
assign pe_2_13_clk = clk;
assign pe_2_13_top =
  _guard7396 ? top_2_13_out :
  32'd0;
assign pe_2_13_left =
  _guard7409 ? left_2_13_out :
  32'd0;
assign pe_2_13_reset = reset;
assign pe_2_13_go = _guard7422;
assign top_2_15_write_en = _guard7425;
assign top_2_15_clk = clk;
assign top_2_15_reset = reset;
assign top_2_15_in = top_1_15_out;
assign pe_3_15_mul_ready =
  _guard7431 ? 1'd1 :
  _guard7434 ? 1'd0 :
  1'd0;
assign pe_3_15_clk = clk;
assign pe_3_15_top =
  _guard7447 ? top_3_15_out :
  32'd0;
assign pe_3_15_left =
  _guard7460 ? left_3_15_out :
  32'd0;
assign pe_3_15_reset = reset;
assign pe_3_15_go = _guard7473;
assign pe_4_5_mul_ready =
  _guard7476 ? 1'd1 :
  _guard7479 ? 1'd0 :
  1'd0;
assign pe_4_5_clk = clk;
assign pe_4_5_top =
  _guard7492 ? top_4_5_out :
  32'd0;
assign pe_4_5_left =
  _guard7505 ? left_4_5_out :
  32'd0;
assign pe_4_5_reset = reset;
assign pe_4_5_go = _guard7518;
assign left_4_5_write_en = _guard7521;
assign left_4_5_clk = clk;
assign left_4_5_reset = reset;
assign left_4_5_in = left_4_4_out;
assign top_4_9_write_en = _guard7527;
assign top_4_9_clk = clk;
assign top_4_9_reset = reset;
assign top_4_9_in = top_3_9_out;
assign left_4_9_write_en = _guard7533;
assign left_4_9_clk = clk;
assign left_4_9_reset = reset;
assign left_4_9_in = left_4_8_out;
assign left_4_14_write_en = _guard7539;
assign left_4_14_clk = clk;
assign left_4_14_reset = reset;
assign left_4_14_in = left_4_13_out;
assign top_5_0_write_en = _guard7545;
assign top_5_0_clk = clk;
assign top_5_0_reset = reset;
assign top_5_0_in = top_4_0_out;
assign top_5_3_write_en = _guard7551;
assign top_5_3_clk = clk;
assign top_5_3_reset = reset;
assign top_5_3_in = top_4_3_out;
assign left_6_8_write_en = _guard7557;
assign left_6_8_clk = clk;
assign left_6_8_reset = reset;
assign left_6_8_in = left_6_7_out;
assign top_7_10_write_en = _guard7563;
assign top_7_10_clk = clk;
assign top_7_10_reset = reset;
assign top_7_10_in = top_6_10_out;
assign top_8_0_write_en = _guard7569;
assign top_8_0_clk = clk;
assign top_8_0_reset = reset;
assign top_8_0_in = top_7_0_out;
assign left_8_5_write_en = _guard7575;
assign left_8_5_clk = clk;
assign left_8_5_reset = reset;
assign left_8_5_in = left_8_4_out;
assign top_8_11_write_en = _guard7581;
assign top_8_11_clk = clk;
assign top_8_11_reset = reset;
assign top_8_11_in = top_7_11_out;
assign pe_8_13_mul_ready =
  _guard7587 ? 1'd1 :
  _guard7590 ? 1'd0 :
  1'd0;
assign pe_8_13_clk = clk;
assign pe_8_13_top =
  _guard7603 ? top_8_13_out :
  32'd0;
assign pe_8_13_left =
  _guard7616 ? left_8_13_out :
  32'd0;
assign pe_8_13_reset = reset;
assign pe_8_13_go = _guard7629;
assign top_9_5_write_en = _guard7632;
assign top_9_5_clk = clk;
assign top_9_5_reset = reset;
assign top_9_5_in = top_8_5_out;
assign left_10_3_write_en = _guard7638;
assign left_10_3_clk = clk;
assign left_10_3_reset = reset;
assign left_10_3_in = left_10_2_out;
assign pe_10_7_mul_ready =
  _guard7644 ? 1'd1 :
  _guard7647 ? 1'd0 :
  1'd0;
assign pe_10_7_clk = clk;
assign pe_10_7_top =
  _guard7660 ? top_10_7_out :
  32'd0;
assign pe_10_7_left =
  _guard7673 ? left_10_7_out :
  32'd0;
assign pe_10_7_reset = reset;
assign pe_10_7_go = _guard7686;
assign pe_10_9_mul_ready =
  _guard7689 ? 1'd1 :
  _guard7692 ? 1'd0 :
  1'd0;
assign pe_10_9_clk = clk;
assign pe_10_9_top =
  _guard7705 ? top_10_9_out :
  32'd0;
assign pe_10_9_left =
  _guard7718 ? left_10_9_out :
  32'd0;
assign pe_10_9_reset = reset;
assign pe_10_9_go = _guard7731;
assign left_11_3_write_en = _guard7734;
assign left_11_3_clk = clk;
assign left_11_3_reset = reset;
assign left_11_3_in = left_11_2_out;
assign pe_11_4_mul_ready =
  _guard7740 ? 1'd1 :
  _guard7743 ? 1'd0 :
  1'd0;
assign pe_11_4_clk = clk;
assign pe_11_4_top =
  _guard7756 ? top_11_4_out :
  32'd0;
assign pe_11_4_left =
  _guard7769 ? left_11_4_out :
  32'd0;
assign pe_11_4_reset = reset;
assign pe_11_4_go = _guard7782;
assign left_12_0_write_en = _guard7785;
assign left_12_0_clk = clk;
assign left_12_0_reset = reset;
assign left_12_0_in = l12_read_data;
assign top_12_10_write_en = _guard7791;
assign top_12_10_clk = clk;
assign top_12_10_reset = reset;
assign top_12_10_in = top_11_10_out;
assign left_12_14_write_en = _guard7797;
assign left_12_14_clk = clk;
assign left_12_14_reset = reset;
assign left_12_14_in = left_12_13_out;
assign pe_13_7_mul_ready =
  _guard7803 ? 1'd1 :
  _guard7806 ? 1'd0 :
  1'd0;
assign pe_13_7_clk = clk;
assign pe_13_7_top =
  _guard7819 ? top_13_7_out :
  32'd0;
assign pe_13_7_left =
  _guard7832 ? left_13_7_out :
  32'd0;
assign pe_13_7_reset = reset;
assign pe_13_7_go = _guard7845;
assign left_13_10_write_en = _guard7848;
assign left_13_10_clk = clk;
assign left_13_10_reset = reset;
assign left_13_10_in = left_13_9_out;
assign left_13_11_write_en = _guard7854;
assign left_13_11_clk = clk;
assign left_13_11_reset = reset;
assign left_13_11_in = left_13_10_out;
assign left_13_15_write_en = _guard7860;
assign left_13_15_clk = clk;
assign left_13_15_reset = reset;
assign left_13_15_in = left_13_14_out;
assign left_14_1_write_en = _guard7866;
assign left_14_1_clk = clk;
assign left_14_1_reset = reset;
assign left_14_1_in = left_14_0_out;
assign top_14_4_write_en = _guard7872;
assign top_14_4_clk = clk;
assign top_14_4_reset = reset;
assign top_14_4_in = top_13_4_out;
assign left_14_7_write_en = _guard7878;
assign left_14_7_clk = clk;
assign left_14_7_reset = reset;
assign left_14_7_in = left_14_6_out;
assign left_14_11_write_en = _guard7884;
assign left_14_11_clk = clk;
assign left_14_11_reset = reset;
assign left_14_11_in = left_14_10_out;
assign left_15_9_write_en = _guard7890;
assign left_15_9_clk = clk;
assign left_15_9_reset = reset;
assign left_15_9_in = left_15_8_out;
assign left_15_11_write_en = _guard7896;
assign left_15_11_clk = clk;
assign left_15_11_reset = reset;
assign left_15_11_in = left_15_10_out;
assign pe_15_14_mul_ready =
  _guard7902 ? 1'd1 :
  _guard7905 ? 1'd0 :
  1'd0;
assign pe_15_14_clk = clk;
assign pe_15_14_top =
  _guard7918 ? top_15_14_out :
  32'd0;
assign pe_15_14_left =
  _guard7931 ? left_15_14_out :
  32'd0;
assign pe_15_14_reset = reset;
assign pe_15_14_go = _guard7944;
assign t10_idx_write_en = _guard7951;
assign t10_idx_clk = clk;
assign t10_idx_reset = reset;
assign t10_idx_in =
  _guard7954 ? 5'd0 :
  _guard7957 ? t10_add_out :
  'x;
assign l3_add_left = 5'd1;
assign l3_add_right = l3_idx_out;
assign l15_add_left = 5'd1;
assign l15_add_right = l15_idx_out;
assign idx_between_16_20_comb_left = index_ge_16_out;
assign idx_between_16_20_comb_right = index_lt_20_out;
assign index_ge_40_left = idx_add_out;
assign index_ge_40_right = 6'd40;
assign idx_between_27_43_comb_left = index_ge_27_out;
assign idx_between_27_43_comb_right = index_lt_43_out;
assign index_lt_19_left = idx_add_out;
assign index_lt_19_right = 6'd19;
assign index_ge_3_left = idx_add_out;
assign index_ge_3_right = 6'd3;
assign idx_between_31_35_reg_write_en = _guard7984;
assign idx_between_31_35_reg_clk = clk;
assign idx_between_31_35_reg_reset = reset;
assign idx_between_31_35_reg_in =
  _guard7987 ? 1'd0 :
  _guard7988 ? idx_between_31_35_comb_out :
  'x;
assign idx_between_5_9_comb_left = index_ge_5_out;
assign idx_between_5_9_comb_right = index_lt_9_out;
assign index_ge_46_left = idx_add_out;
assign index_ge_46_right = 6'd46;
assign idx_between_30_31_comb_left = index_ge_30_out;
assign idx_between_30_31_comb_right = index_lt_31_out;
assign index_ge_12_left = idx_add_out;
assign index_ge_12_right = 6'd12;
assign idx_between_4_8_reg_write_en = _guard8001;
assign idx_between_4_8_reg_clk = clk;
assign idx_between_4_8_reg_reset = reset;
assign idx_between_4_8_reg_in =
  _guard8004 ? 1'd0 :
  _guard8005 ? idx_between_4_8_comb_out :
  'x;
assign idx_between_10_14_comb_left = index_ge_10_out;
assign idx_between_10_14_comb_right = index_lt_14_out;
assign idx_between_6_10_comb_left = index_ge_6_out;
assign idx_between_6_10_comb_right = index_lt_10_out;
assign idx_between_13_29_reg_write_en = _guard8014;
assign idx_between_13_29_reg_clk = clk;
assign idx_between_13_29_reg_reset = reset;
assign idx_between_13_29_reg_in =
  _guard8015 ? idx_between_13_29_comb_out :
  _guard8018 ? 1'd0 :
  'x;
assign idx_between_9_13_comb_left = index_ge_9_out;
assign idx_between_9_13_comb_right = index_lt_13_out;
assign index_ge_37_left = idx_add_out;
assign index_ge_37_right = 6'd37;
assign index_lt_40_left = idx_add_out;
assign index_lt_40_right = 6'd40;
assign idx_between_34_35_comb_left = index_ge_34_out;
assign idx_between_34_35_comb_right = index_lt_35_out;
assign idx_between_2_18_comb_left = index_ge_2_out;
assign idx_between_2_18_comb_right = index_lt_18_out;
assign cond_write_en = _guard8029;
assign cond_clk = clk;
assign cond_reset = reset;
assign cond_in =
  _guard8030 ? idx_between_0_16_reg_out :
  1'd0;
assign cond_wire26_in =
  _guard8031 ? idx_between_6_22_reg_out :
  _guard8034 ? cond26_out :
  1'd0;
assign cond35_write_en = _guard8035;
assign cond35_clk = clk;
assign cond35_reset = reset;
assign cond35_in =
  _guard8036 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire35_in =
  _guard8039 ? cond35_out :
  _guard8040 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire50_in =
  _guard8043 ? cond50_out :
  _guard8044 ? idx_between_11_15_reg_out :
  1'd0;
assign cond_wire56_in =
  _guard8047 ? cond56_out :
  _guard8048 ? idx_between_12_28_reg_out :
  1'd0;
assign cond60_write_en = _guard8049;
assign cond60_clk = clk;
assign cond60_reset = reset;
assign cond60_in =
  _guard8050 ? idx_between_13_17_reg_out :
  1'd0;
assign cond69_write_en = _guard8051;
assign cond69_clk = clk;
assign cond69_reset = reset;
assign cond69_in =
  _guard8052 ? idx_between_14_30_reg_out :
  1'd0;
assign cond72_write_en = _guard8053;
assign cond72_clk = clk;
assign cond72_reset = reset;
assign cond72_in =
  _guard8054 ? idx_between_19_35_reg_out :
  1'd0;
assign cond76_write_en = _guard8055;
assign cond76_clk = clk;
assign cond76_reset = reset;
assign cond76_in =
  _guard8056 ? idx_between_16_32_reg_out :
  1'd0;
assign cond_wire85_in =
  _guard8057 ? idx_between_3_19_reg_out :
  _guard8060 ? cond85_out :
  1'd0;
assign cond92_write_en = _guard8061;
assign cond92_clk = clk;
assign cond92_reset = reset;
assign cond92_in =
  _guard8062 ? idx_between_5_9_reg_out :
  1'd0;
assign cond_wire116_in =
  _guard8065 ? cond116_out :
  _guard8066 ? idx_between_11_15_reg_out :
  1'd0;
assign cond_wire149_in =
  _guard8069 ? cond149_out :
  _guard8070 ? idx_between_4_8_reg_out :
  1'd0;
assign cond_wire163_in =
  _guard8071 ? idx_between_11_27_reg_out :
  _guard8074 ? cond163_out :
  1'd0;
assign cond_wire182_in =
  _guard8075 ? idx_between_12_28_reg_out :
  _guard8078 ? cond182_out :
  1'd0;
assign cond189_write_en = _guard8079;
assign cond189_clk = clk;
assign cond189_reset = reset;
assign cond189_in =
  _guard8080 ? idx_between_14_18_reg_out :
  1'd0;
assign cond_wire192_in =
  _guard8081 ? idx_between_34_35_reg_out :
  _guard8084 ? cond192_out :
  1'd0;
assign cond_wire200_in =
  _guard8085 ? idx_between_36_37_reg_out :
  _guard8088 ? cond200_out :
  1'd0;
assign cond_wire205_in =
  _guard8091 ? cond205_out :
  _guard8092 ? idx_between_18_22_reg_out :
  1'd0;
assign cond226_write_en = _guard8093;
assign cond226_clk = clk;
assign cond226_reset = reset;
assign cond226_in =
  _guard8094 ? idx_between_8_12_reg_out :
  1'd0;
assign cond233_write_en = _guard8095;
assign cond233_clk = clk;
assign cond233_reset = reset;
assign cond233_in =
  _guard8096 ? idx_between_29_30_reg_out :
  1'd0;
assign cond241_write_en = _guard8097;
assign cond241_clk = clk;
assign cond241_reset = reset;
assign cond241_in =
  _guard8098 ? idx_between_31_32_reg_out :
  1'd0;
assign cond_wire243_in =
  _guard8099 ? idx_between_12_28_reg_out :
  _guard8102 ? cond243_out :
  1'd0;
assign cond_wire245_in =
  _guard8105 ? cond245_out :
  _guard8106 ? idx_between_32_33_reg_out :
  1'd0;
assign cond248_write_en = _guard8107;
assign cond248_clk = clk;
assign cond248_reset = reset;
assign cond248_in =
  _guard8108 ? idx_between_17_33_reg_out :
  1'd0;
assign cond257_write_en = _guard8109;
assign cond257_clk = clk;
assign cond257_reset = reset;
assign cond257_in =
  _guard8110 ? idx_between_35_36_reg_out :
  1'd0;
assign cond_wire263_in =
  _guard8113 ? cond263_out :
  _guard8114 ? idx_between_17_33_reg_out :
  1'd0;
assign cond266_write_en = _guard8115;
assign cond266_clk = clk;
assign cond266_reset = reset;
assign cond266_in =
  _guard8116 ? idx_between_18_22_reg_out :
  1'd0;
assign cond_wire273_in =
  _guard8117 ? idx_between_39_40_reg_out :
  _guard8120 ? cond273_out :
  1'd0;
assign cond284_write_en = _guard8121;
assign cond284_clk = clk;
assign cond284_reset = reset;
assign cond284_in =
  _guard8122 ? idx_between_7_23_reg_out :
  1'd0;
assign cond309_write_en = _guard8123;
assign cond309_clk = clk;
assign cond309_reset = reset;
assign cond309_in =
  _guard8124 ? idx_between_17_33_reg_out :
  1'd0;
assign cond_wire310_in =
  _guard8125 ? idx_between_33_34_reg_out :
  _guard8128 ? cond310_out :
  1'd0;
assign cond319_write_en = _guard8129;
assign cond319_clk = clk;
assign cond319_reset = reset;
assign cond319_in =
  _guard8130 ? idx_between_16_20_reg_out :
  1'd0;
assign cond_wire325_in =
  _guard8133 ? cond325_out :
  _guard8134 ? idx_between_21_37_reg_out :
  1'd0;
assign cond333_write_en = _guard8135;
assign cond333_clk = clk;
assign cond333_reset = reset;
assign cond333_in =
  _guard8136 ? idx_between_23_39_reg_out :
  1'd0;
assign cond_wire334_in =
  _guard8137 ? idx_between_39_40_reg_out :
  _guard8140 ? cond334_out :
  1'd0;
assign cond357_write_en = _guard8141;
assign cond357_clk = clk;
assign cond357_reset = reset;
assign cond357_in =
  _guard8142 ? idx_between_10_26_reg_out :
  1'd0;
assign cond_wire374_in =
  _guard8143 ? idx_between_18_34_reg_out :
  _guard8146 ? cond374_out :
  1'd0;
assign cond_wire384_in =
  _guard8147 ? idx_between_17_21_reg_out :
  _guard8150 ? cond384_out :
  1'd0;
assign cond386_write_en = _guard8151;
assign cond386_clk = clk;
assign cond386_reset = reset;
assign cond386_in =
  _guard8152 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire395_in =
  _guard8155 ? cond395_out :
  _guard8156 ? idx_between_39_40_reg_out :
  1'd0;
assign cond416_write_en = _guard8157;
assign cond416_clk = clk;
assign cond416_reset = reset;
assign cond416_in =
  _guard8158 ? idx_between_29_30_reg_out :
  1'd0;
assign cond421_write_en = _guard8159;
assign cond421_clk = clk;
assign cond421_reset = reset;
assign cond421_in =
  _guard8160 ? idx_between_11_15_reg_out :
  1'd0;
assign cond443_write_en = _guard8161;
assign cond443_clk = clk;
assign cond443_reset = reset;
assign cond443_in =
  _guard8162 ? idx_between_20_36_reg_out :
  1'd0;
assign cond446_write_en = _guard8163;
assign cond446_clk = clk;
assign cond446_reset = reset;
assign cond446_in =
  _guard8164 ? idx_between_17_33_reg_out :
  1'd0;
assign cond455_write_en = _guard8165;
assign cond455_clk = clk;
assign cond455_reset = reset;
assign cond455_in =
  _guard8166 ? idx_between_23_39_reg_out :
  1'd0;
assign cond_wire458_in =
  _guard8169 ? cond458_out :
  _guard8170 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire459_in =
  _guard8173 ? cond459_out :
  _guard8174 ? idx_between_24_40_reg_out :
  1'd0;
assign cond474_write_en = _guard8175;
assign cond474_clk = clk;
assign cond474_reset = reset;
assign cond474_in =
  _guard8176 ? idx_between_9_13_reg_out :
  1'd0;
assign cond475_write_en = _guard8177;
assign cond475_clk = clk;
assign cond475_reset = reset;
assign cond475_in =
  _guard8178 ? idx_between_9_25_reg_out :
  1'd0;
assign cond485_write_en = _guard8179;
assign cond485_clk = clk;
assign cond485_reset = reset;
assign cond485_in =
  _guard8180 ? idx_between_31_32_reg_out :
  1'd0;
assign cond506_write_en = _guard8181;
assign cond506_clk = clk;
assign cond506_reset = reset;
assign cond506_in =
  _guard8182 ? idx_between_17_21_reg_out :
  1'd0;
assign cond_wire533_in =
  _guard8183 ? idx_between_43_44_reg_out :
  _guard8186 ? cond533_out :
  1'd0;
assign cond_wire541_in =
  _guard8187 ? idx_between_14_30_reg_out :
  _guard8190 ? cond541_out :
  1'd0;
assign cond_wire545_in =
  _guard8193 ? cond545_out :
  _guard8194 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire552_in =
  _guard8195 ? idx_between_13_29_reg_out :
  _guard8198 ? cond552_out :
  1'd0;
assign cond_wire560_in =
  _guard8201 ? cond560_out :
  _guard8202 ? idx_between_15_31_reg_out :
  1'd0;
assign cond561_write_en = _guard8203;
assign cond561_clk = clk;
assign cond561_reset = reset;
assign cond561_in =
  _guard8204 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire573_in =
  _guard8207 ? cond573_out :
  _guard8208 ? idx_between_22_38_reg_out :
  1'd0;
assign cond578_write_en = _guard8209;
assign cond578_clk = clk;
assign cond578_reset = reset;
assign cond578_in =
  _guard8210 ? idx_between_39_40_reg_out :
  1'd0;
assign cond584_write_en = _guard8211;
assign cond584_clk = clk;
assign cond584_reset = reset;
assign cond584_in =
  _guard8212 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire586_in =
  _guard8215 ? cond586_out :
  _guard8216 ? idx_between_41_42_reg_out :
  1'd0;
assign cond589_write_en = _guard8217;
assign cond589_clk = clk;
assign cond589_reset = reset;
assign cond589_in =
  _guard8218 ? idx_between_26_42_reg_out :
  1'd0;
assign cond592_write_en = _guard8219;
assign cond592_clk = clk;
assign cond592_reset = reset;
assign cond592_in =
  _guard8220 ? idx_between_23_39_reg_out :
  1'd0;
assign cond597_write_en = _guard8221;
assign cond597_clk = clk;
assign cond597_reset = reset;
assign cond597_in =
  _guard8222 ? idx_between_28_44_reg_out :
  1'd0;
assign cond_wire604_in =
  _guard8225 ? cond604_out :
  _guard8226 ? idx_between_11_15_reg_out :
  1'd0;
assign cond606_write_en = _guard8227;
assign cond606_clk = clk;
assign cond606_reset = reset;
assign cond606_in =
  _guard8228 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire610_in =
  _guard8229 ? idx_between_16_32_reg_out :
  _guard8232 ? cond610_out :
  1'd0;
assign cond614_write_en = _guard8233;
assign cond614_clk = clk;
assign cond614_reset = reset;
assign cond614_in =
  _guard8234 ? idx_between_17_33_reg_out :
  1'd0;
assign cond_wire617_in =
  _guard8235 ? idx_between_14_30_reg_out :
  _guard8238 ? cond617_out :
  1'd0;
assign cond_wire635_in =
  _guard8241 ? cond635_out :
  _guard8242 ? idx_between_38_39_reg_out :
  1'd0;
assign cond636_write_en = _guard8243;
assign cond636_clk = clk;
assign cond636_reset = reset;
assign cond636_in =
  _guard8244 ? idx_between_19_23_reg_out :
  1'd0;
assign cond_wire636_in =
  _guard8245 ? idx_between_19_23_reg_out :
  _guard8248 ? cond636_out :
  1'd0;
assign cond_wire637_in =
  _guard8251 ? cond637_out :
  _guard8252 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire645_in =
  _guard8253 ? idx_between_21_37_reg_out :
  _guard8256 ? cond645_out :
  1'd0;
assign cond655_write_en = _guard8257;
assign cond655_clk = clk;
assign cond655_reset = reset;
assign cond655_in =
  _guard8258 ? idx_between_43_44_reg_out :
  1'd0;
assign cond_wire656_in =
  _guard8261 ? cond656_out :
  _guard8262 ? idx_between_24_28_reg_out :
  1'd0;
assign cond_wire661_in =
  _guard8265 ? cond661_out :
  _guard8266 ? idx_between_25_41_reg_out :
  1'd0;
assign cond663_write_en = _guard8267;
assign cond663_clk = clk;
assign cond663_reset = reset;
assign cond663_in =
  _guard8268 ? idx_between_45_46_reg_out :
  1'd0;
assign cond665_write_en = _guard8269;
assign cond665_clk = clk;
assign cond665_reset = reset;
assign cond665_in =
  _guard8270 ? idx_between_11_15_reg_out :
  1'd0;
assign cond683_write_en = _guard8271;
assign cond683_clk = clk;
assign cond683_reset = reset;
assign cond683_in =
  _guard8272 ? idx_between_19_35_reg_out :
  1'd0;
assign cond684_write_en = _guard8273;
assign cond684_clk = clk;
assign cond684_reset = reset;
assign cond684_in =
  _guard8274 ? idx_between_35_36_reg_out :
  1'd0;
assign cond_wire691_in =
  _guard8275 ? idx_between_21_37_reg_out :
  _guard8278 ? cond691_out :
  1'd0;
assign cond710_write_en = _guard8279;
assign cond710_clk = clk;
assign cond710_reset = reset;
assign cond710_in =
  _guard8280 ? idx_between_22_38_reg_out :
  1'd0;
assign cond723_write_en = _guard8281;
assign cond723_clk = clk;
assign cond723_reset = reset;
assign cond723_in =
  _guard8282 ? idx_between_29_45_reg_out :
  1'd0;
assign cond742_write_en = _guard8283;
assign cond742_clk = clk;
assign cond742_reset = reset;
assign cond742_in =
  _guard8284 ? idx_between_15_19_reg_out :
  1'd0;
assign cond745_write_en = _guard8285;
assign cond745_clk = clk;
assign cond745_reset = reset;
assign cond745_in =
  _guard8286 ? idx_between_35_36_reg_out :
  1'd0;
assign cond747_write_en = _guard8287;
assign cond747_clk = clk;
assign cond747_reset = reset;
assign cond747_in =
  _guard8288 ? idx_between_16_32_reg_out :
  1'd0;
assign cond751_write_en = _guard8289;
assign cond751_clk = clk;
assign cond751_reset = reset;
assign cond751_in =
  _guard8290 ? idx_between_17_33_reg_out :
  1'd0;
assign cond755_write_en = _guard8291;
assign cond755_clk = clk;
assign cond755_reset = reset;
assign cond755_in =
  _guard8292 ? idx_between_18_34_reg_out :
  1'd0;
assign cond786_write_en = _guard8293;
assign cond786_clk = clk;
assign cond786_reset = reset;
assign cond786_in =
  _guard8294 ? idx_between_26_30_reg_out :
  1'd0;
assign cond791_write_en = _guard8295;
assign cond791_clk = clk;
assign cond791_reset = reset;
assign cond791_in =
  _guard8296 ? idx_between_27_43_reg_out :
  1'd0;
assign cond_wire797_in =
  _guard8297 ? idx_between_17_33_reg_out :
  _guard8300 ? cond797_out :
  1'd0;
assign cond800_write_en = _guard8301;
assign cond800_clk = clk;
assign cond800_reset = reset;
assign cond800_in =
  _guard8302 ? idx_between_14_30_reg_out :
  1'd0;
assign cond_wire822_in =
  _guard8305 ? cond822_out :
  _guard8306 ? idx_between_39_40_reg_out :
  1'd0;
assign cond_wire826_in =
  _guard8309 ? cond826_out :
  _guard8310 ? idx_between_40_41_reg_out :
  1'd0;
assign cond827_write_en = _guard8311;
assign cond827_clk = clk;
assign cond827_reset = reset;
assign cond827_in =
  _guard8312 ? idx_between_21_25_reg_out :
  1'd0;
assign cond_wire831_in =
  _guard8313 ? idx_between_22_26_reg_out :
  _guard8316 ? cond831_out :
  1'd0;
assign cond835_write_en = _guard8317;
assign cond835_clk = clk;
assign cond835_reset = reset;
assign cond835_in =
  _guard8318 ? idx_between_23_27_reg_out :
  1'd0;
assign cond_wire842_in =
  _guard8319 ? idx_between_44_45_reg_out :
  _guard8322 ? cond842_out :
  1'd0;
assign cond852_write_en = _guard8323;
assign cond852_clk = clk;
assign cond852_reset = reset;
assign cond852_in =
  _guard8324 ? idx_between_27_43_reg_out :
  1'd0;
assign cond853_write_en = _guard8325;
assign cond853_clk = clk;
assign cond853_reset = reset;
assign cond853_in =
  _guard8326 ? idx_between_31_47_reg_out :
  1'd0;
assign cond864_write_en = _guard8327;
assign cond864_clk = clk;
assign cond864_reset = reset;
assign cond864_in =
  _guard8328 ? idx_between_15_19_reg_out :
  1'd0;
assign cond867_write_en = _guard8329;
assign cond867_clk = clk;
assign cond867_reset = reset;
assign cond867_in =
  _guard8330 ? idx_between_35_36_reg_out :
  1'd0;
assign cond868_write_en = _guard8331;
assign cond868_clk = clk;
assign cond868_reset = reset;
assign cond868_in =
  _guard8332 ? idx_between_16_20_reg_out :
  1'd0;
assign cond880_write_en = _guard8333;
assign cond880_clk = clk;
assign cond880_reset = reset;
assign cond880_in =
  _guard8334 ? idx_between_19_23_reg_out :
  1'd0;
assign cond894_write_en = _guard8335;
assign cond894_clk = clk;
assign cond894_reset = reset;
assign cond894_in =
  _guard8336 ? idx_between_26_42_reg_out :
  1'd0;
assign cond901_write_en = _guard8337;
assign cond901_clk = clk;
assign cond901_reset = reset;
assign cond901_in =
  _guard8338 ? idx_between_24_40_reg_out :
  1'd0;
assign cond_wire901_in =
  _guard8341 ? cond901_out :
  _guard8342 ? idx_between_24_40_reg_out :
  1'd0;
assign cond_wire920_in =
  _guard8343 ? idx_between_29_33_reg_out :
  _guard8346 ? cond920_out :
  1'd0;
assign cond_wire925_in =
  _guard8347 ? idx_between_15_19_reg_out :
  _guard8350 ? cond925_out :
  1'd0;
assign cond943_write_en = _guard8351;
assign cond943_clk = clk;
assign cond943_reset = reset;
assign cond943_in =
  _guard8352 ? idx_between_23_39_reg_out :
  1'd0;
assign cond945_write_en = _guard8353;
assign cond945_clk = clk;
assign cond945_reset = reset;
assign cond945_in =
  _guard8354 ? idx_between_20_24_reg_out :
  1'd0;
assign cond_wire946_in =
  _guard8355 ? idx_between_20_36_reg_out :
  _guard8358 ? cond946_out :
  1'd0;
assign cond_wire955_in =
  _guard8361 ? cond955_out :
  _guard8362 ? idx_between_26_42_reg_out :
  1'd0;
assign cond_wire977_in =
  _guard8365 ? cond977_out :
  _guard8366 ? idx_between_28_32_reg_out :
  1'd0;
assign cond_wire984_in =
  _guard8369 ? cond984_out :
  _guard8370 ? idx_between_49_50_reg_out :
  1'd0;
assign cond993_write_en = _guard8371;
assign cond993_clk = clk;
assign cond993_reset = reset;
assign cond993_in =
  _guard8372 ? idx_between_36_37_reg_out :
  1'd0;
assign cond1000_write_en = _guard8373;
assign cond1000_clk = clk;
assign cond1000_reset = reset;
assign cond1000_in =
  _guard8374 ? idx_between_22_38_reg_out :
  1'd0;
assign cond1012_write_en = _guard8375;
assign cond1012_clk = clk;
assign cond1012_reset = reset;
assign cond1012_in =
  _guard8376 ? idx_between_25_41_reg_out :
  1'd0;
assign cond1024_write_en = _guard8377;
assign cond1024_clk = clk;
assign cond1024_reset = reset;
assign cond1024_in =
  _guard8378 ? idx_between_28_44_reg_out :
  1'd0;
assign cond_wire1028_in =
  _guard8379 ? idx_between_29_45_reg_out :
  _guard8382 ? cond1028_out :
  1'd0;
assign cond_wire1029_in =
  _guard8385 ? cond1029_out :
  _guard8386 ? idx_between_45_46_reg_out :
  1'd0;
assign cond1041_write_en = _guard8387;
assign cond1041_clk = clk;
assign cond1041_reset = reset;
assign cond1041_in =
  _guard8388 ? idx_between_48_49_reg_out :
  1'd0;
assign cond1044_write_en = _guard8389;
assign cond1044_clk = clk;
assign cond1044_reset = reset;
assign cond1044_in =
  _guard8390 ? idx_between_33_49_reg_out :
  1'd0;
assign cond_wire1051_in =
  _guard8391 ? idx_between_35_51_reg_out :
  _guard8394 ? cond1051_out :
  1'd0;
assign left_0_12_write_en = _guard8397;
assign left_0_12_clk = clk;
assign left_0_12_reset = reset;
assign left_0_12_in = left_0_11_out;
assign pe_1_0_mul_ready =
  _guard8403 ? 1'd1 :
  _guard8406 ? 1'd0 :
  1'd0;
assign pe_1_0_clk = clk;
assign pe_1_0_top =
  _guard8419 ? top_1_0_out :
  32'd0;
assign pe_1_0_left =
  _guard8432 ? left_1_0_out :
  32'd0;
assign pe_1_0_reset = reset;
assign pe_1_0_go = _guard8445;
assign left_1_0_write_en = _guard8448;
assign left_1_0_clk = clk;
assign left_1_0_reset = reset;
assign left_1_0_in = l1_read_data;
assign left_1_1_write_en = _guard8454;
assign left_1_1_clk = clk;
assign left_1_1_reset = reset;
assign left_1_1_in = left_1_0_out;
assign top_1_2_write_en = _guard8460;
assign top_1_2_clk = clk;
assign top_1_2_reset = reset;
assign top_1_2_in = top_0_2_out;
assign left_1_11_write_en = _guard8466;
assign left_1_11_clk = clk;
assign left_1_11_reset = reset;
assign left_1_11_in = left_1_10_out;
assign top_1_15_write_en = _guard8472;
assign top_1_15_clk = clk;
assign top_1_15_reset = reset;
assign top_1_15_in = top_0_15_out;
assign left_2_0_write_en = _guard8478;
assign left_2_0_clk = clk;
assign left_2_0_reset = reset;
assign left_2_0_in = l2_read_data;
assign left_2_9_write_en = _guard8484;
assign left_2_9_clk = clk;
assign left_2_9_reset = reset;
assign left_2_9_in = left_2_8_out;
assign top_2_12_write_en = _guard8490;
assign top_2_12_clk = clk;
assign top_2_12_reset = reset;
assign top_2_12_in = top_1_12_out;
assign left_3_1_write_en = _guard8496;
assign left_3_1_clk = clk;
assign left_3_1_reset = reset;
assign left_3_1_in = left_3_0_out;
assign pe_3_2_mul_ready =
  _guard8502 ? 1'd1 :
  _guard8505 ? 1'd0 :
  1'd0;
assign pe_3_2_clk = clk;
assign pe_3_2_top =
  _guard8518 ? top_3_2_out :
  32'd0;
assign pe_3_2_left =
  _guard8531 ? left_3_2_out :
  32'd0;
assign pe_3_2_reset = reset;
assign pe_3_2_go = _guard8544;
assign pe_3_5_mul_ready =
  _guard8547 ? 1'd1 :
  _guard8550 ? 1'd0 :
  1'd0;
assign pe_3_5_clk = clk;
assign pe_3_5_top =
  _guard8563 ? top_3_5_out :
  32'd0;
assign pe_3_5_left =
  _guard8576 ? left_3_5_out :
  32'd0;
assign pe_3_5_reset = reset;
assign pe_3_5_go = _guard8589;
assign pe_3_6_mul_ready =
  _guard8592 ? 1'd1 :
  _guard8595 ? 1'd0 :
  1'd0;
assign pe_3_6_clk = clk;
assign pe_3_6_top =
  _guard8608 ? top_3_6_out :
  32'd0;
assign pe_3_6_left =
  _guard8621 ? left_3_6_out :
  32'd0;
assign pe_3_6_reset = reset;
assign pe_3_6_go = _guard8634;
assign left_3_7_write_en = _guard8637;
assign left_3_7_clk = clk;
assign left_3_7_reset = reset;
assign left_3_7_in = left_3_6_out;
assign left_3_11_write_en = _guard8643;
assign left_3_11_clk = clk;
assign left_3_11_reset = reset;
assign left_3_11_in = left_3_10_out;
assign left_3_13_write_en = _guard8649;
assign left_3_13_clk = clk;
assign left_3_13_reset = reset;
assign left_3_13_in = left_3_12_out;
assign top_4_5_write_en = _guard8655;
assign top_4_5_clk = clk;
assign top_4_5_reset = reset;
assign top_4_5_in = top_3_5_out;
assign pe_5_4_mul_ready =
  _guard8661 ? 1'd1 :
  _guard8664 ? 1'd0 :
  1'd0;
assign pe_5_4_clk = clk;
assign pe_5_4_top =
  _guard8677 ? top_5_4_out :
  32'd0;
assign pe_5_4_left =
  _guard8690 ? left_5_4_out :
  32'd0;
assign pe_5_4_reset = reset;
assign pe_5_4_go = _guard8703;
assign top_7_2_write_en = _guard8706;
assign top_7_2_clk = clk;
assign top_7_2_reset = reset;
assign top_7_2_in = top_6_2_out;
assign pe_7_4_mul_ready =
  _guard8712 ? 1'd1 :
  _guard8715 ? 1'd0 :
  1'd0;
assign pe_7_4_clk = clk;
assign pe_7_4_top =
  _guard8728 ? top_7_4_out :
  32'd0;
assign pe_7_4_left =
  _guard8741 ? left_7_4_out :
  32'd0;
assign pe_7_4_reset = reset;
assign pe_7_4_go = _guard8754;
assign left_7_8_write_en = _guard8757;
assign left_7_8_clk = clk;
assign left_7_8_reset = reset;
assign left_7_8_in = left_7_7_out;
assign top_7_11_write_en = _guard8763;
assign top_7_11_clk = clk;
assign top_7_11_reset = reset;
assign top_7_11_in = top_6_11_out;
assign pe_8_1_mul_ready =
  _guard8769 ? 1'd1 :
  _guard8772 ? 1'd0 :
  1'd0;
assign pe_8_1_clk = clk;
assign pe_8_1_top =
  _guard8785 ? top_8_1_out :
  32'd0;
assign pe_8_1_left =
  _guard8798 ? left_8_1_out :
  32'd0;
assign pe_8_1_reset = reset;
assign pe_8_1_go = _guard8811;
assign left_8_2_write_en = _guard8814;
assign left_8_2_clk = clk;
assign left_8_2_reset = reset;
assign left_8_2_in = left_8_1_out;
assign left_8_7_write_en = _guard8820;
assign left_8_7_clk = clk;
assign left_8_7_reset = reset;
assign left_8_7_in = left_8_6_out;
assign top_9_4_write_en = _guard8826;
assign top_9_4_clk = clk;
assign top_9_4_reset = reset;
assign top_9_4_in = top_8_4_out;
assign left_9_4_write_en = _guard8832;
assign left_9_4_clk = clk;
assign left_9_4_reset = reset;
assign left_9_4_in = left_9_3_out;
assign pe_9_9_mul_ready =
  _guard8838 ? 1'd1 :
  _guard8841 ? 1'd0 :
  1'd0;
assign pe_9_9_clk = clk;
assign pe_9_9_top =
  _guard8854 ? top_9_9_out :
  32'd0;
assign pe_9_9_left =
  _guard8867 ? left_9_9_out :
  32'd0;
assign pe_9_9_reset = reset;
assign pe_9_9_go = _guard8880;
assign top_9_12_write_en = _guard8883;
assign top_9_12_clk = clk;
assign top_9_12_reset = reset;
assign top_9_12_in = top_8_12_out;
assign pe_9_13_mul_ready =
  _guard8889 ? 1'd1 :
  _guard8892 ? 1'd0 :
  1'd0;
assign pe_9_13_clk = clk;
assign pe_9_13_top =
  _guard8905 ? top_9_13_out :
  32'd0;
assign pe_9_13_left =
  _guard8918 ? left_9_13_out :
  32'd0;
assign pe_9_13_reset = reset;
assign pe_9_13_go = _guard8931;
assign top_10_2_write_en = _guard8934;
assign top_10_2_clk = clk;
assign top_10_2_reset = reset;
assign top_10_2_in = top_9_2_out;
assign pe_10_8_mul_ready =
  _guard8940 ? 1'd1 :
  _guard8943 ? 1'd0 :
  1'd0;
assign pe_10_8_clk = clk;
assign pe_10_8_top =
  _guard8956 ? top_10_8_out :
  32'd0;
assign pe_10_8_left =
  _guard8969 ? left_10_8_out :
  32'd0;
assign pe_10_8_reset = reset;
assign pe_10_8_go = _guard8982;
assign pe_10_13_mul_ready =
  _guard8985 ? 1'd1 :
  _guard8988 ? 1'd0 :
  1'd0;
assign pe_10_13_clk = clk;
assign pe_10_13_top =
  _guard9001 ? top_10_13_out :
  32'd0;
assign pe_10_13_left =
  _guard9014 ? left_10_13_out :
  32'd0;
assign pe_10_13_reset = reset;
assign pe_10_13_go = _guard9027;
assign top_11_8_write_en = _guard9030;
assign top_11_8_clk = clk;
assign top_11_8_reset = reset;
assign top_11_8_in = top_10_8_out;
assign left_11_8_write_en = _guard9036;
assign left_11_8_clk = clk;
assign left_11_8_reset = reset;
assign left_11_8_in = left_11_7_out;
assign left_12_13_write_en = _guard9042;
assign left_12_13_clk = clk;
assign left_12_13_reset = reset;
assign left_12_13_in = left_12_12_out;
assign top_13_5_write_en = _guard9048;
assign top_13_5_clk = clk;
assign top_13_5_reset = reset;
assign top_13_5_in = top_12_5_out;
assign pe_14_1_mul_ready =
  _guard9054 ? 1'd1 :
  _guard9057 ? 1'd0 :
  1'd0;
assign pe_14_1_clk = clk;
assign pe_14_1_top =
  _guard9070 ? top_14_1_out :
  32'd0;
assign pe_14_1_left =
  _guard9083 ? left_14_1_out :
  32'd0;
assign pe_14_1_reset = reset;
assign pe_14_1_go = _guard9096;
assign pe_14_7_mul_ready =
  _guard9099 ? 1'd1 :
  _guard9102 ? 1'd0 :
  1'd0;
assign pe_14_7_clk = clk;
assign pe_14_7_top =
  _guard9115 ? top_14_7_out :
  32'd0;
assign pe_14_7_left =
  _guard9128 ? left_14_7_out :
  32'd0;
assign pe_14_7_reset = reset;
assign pe_14_7_go = _guard9141;
assign pe_14_8_mul_ready =
  _guard9144 ? 1'd1 :
  _guard9147 ? 1'd0 :
  1'd0;
assign pe_14_8_clk = clk;
assign pe_14_8_top =
  _guard9160 ? top_14_8_out :
  32'd0;
assign pe_14_8_left =
  _guard9173 ? left_14_8_out :
  32'd0;
assign pe_14_8_reset = reset;
assign pe_14_8_go = _guard9186;
assign pe_14_9_mul_ready =
  _guard9189 ? 1'd1 :
  _guard9192 ? 1'd0 :
  1'd0;
assign pe_14_9_clk = clk;
assign pe_14_9_top =
  _guard9205 ? top_14_9_out :
  32'd0;
assign pe_14_9_left =
  _guard9218 ? left_14_9_out :
  32'd0;
assign pe_14_9_reset = reset;
assign pe_14_9_go = _guard9231;
assign top_14_9_write_en = _guard9234;
assign top_14_9_clk = clk;
assign top_14_9_reset = reset;
assign top_14_9_in = top_13_9_out;
assign top_14_11_write_en = _guard9240;
assign top_14_11_clk = clk;
assign top_14_11_reset = reset;
assign top_14_11_in = top_13_11_out;
assign pe_14_14_mul_ready =
  _guard9246 ? 1'd1 :
  _guard9249 ? 1'd0 :
  1'd0;
assign pe_14_14_clk = clk;
assign pe_14_14_top =
  _guard9262 ? top_14_14_out :
  32'd0;
assign pe_14_14_left =
  _guard9275 ? left_14_14_out :
  32'd0;
assign pe_14_14_reset = reset;
assign pe_14_14_go = _guard9288;
assign left_14_15_write_en = _guard9291;
assign left_14_15_clk = clk;
assign left_14_15_reset = reset;
assign left_14_15_in = left_14_14_out;
assign pe_15_9_mul_ready =
  _guard9297 ? 1'd1 :
  _guard9300 ? 1'd0 :
  1'd0;
assign pe_15_9_clk = clk;
assign pe_15_9_top =
  _guard9313 ? top_15_9_out :
  32'd0;
assign pe_15_9_left =
  _guard9326 ? left_15_9_out :
  32'd0;
assign pe_15_9_reset = reset;
assign pe_15_9_go = _guard9339;
assign top_15_9_write_en = _guard9342;
assign top_15_9_clk = clk;
assign top_15_9_reset = reset;
assign top_15_9_in = top_14_9_out;
assign top_15_11_write_en = _guard9348;
assign top_15_11_clk = clk;
assign top_15_11_reset = reset;
assign top_15_11_in = top_14_11_out;
assign left_15_14_write_en = _guard9354;
assign left_15_14_clk = clk;
assign left_15_14_reset = reset;
assign left_15_14_in = left_15_13_out;
assign t1_idx_write_en = _guard9364;
assign t1_idx_clk = clk;
assign t1_idx_reset = reset;
assign t1_idx_in =
  _guard9367 ? 5'd0 :
  _guard9370 ? t1_add_out :
  'x;
assign t7_idx_write_en = _guard9377;
assign t7_idx_clk = clk;
assign t7_idx_reset = reset;
assign t7_idx_in =
  _guard9380 ? 5'd0 :
  _guard9383 ? t7_add_out :
  'x;
assign t9_idx_write_en = _guard9390;
assign t9_idx_clk = clk;
assign t9_idx_reset = reset;
assign t9_idx_in =
  _guard9393 ? 5'd0 :
  _guard9396 ? t9_add_out :
  'x;
assign l9_idx_write_en = _guard9403;
assign l9_idx_clk = clk;
assign l9_idx_reset = reset;
assign l9_idx_in =
  _guard9406 ? 5'd0 :
  _guard9409 ? l9_add_out :
  'x;
assign l13_add_left = 5'd1;
assign l13_add_right = l13_idx_out;
assign idx_between_25_41_comb_left = index_ge_25_out;
assign idx_between_25_41_comb_right = index_lt_41_out;
assign idx_between_22_26_comb_left = index_ge_22_out;
assign idx_between_22_26_comb_right = index_lt_26_out;
assign idx_between_21_37_comb_left = index_ge_21_out;
assign idx_between_21_37_comb_right = index_lt_37_out;
assign idx_between_3_19_reg_write_en = _guard9426;
assign idx_between_3_19_reg_clk = clk;
assign idx_between_3_19_reg_reset = reset;
assign idx_between_3_19_reg_in =
  _guard9429 ? 1'd0 :
  _guard9430 ? idx_between_3_19_comb_out :
  'x;
assign idx_between_23_24_comb_left = index_ge_23_out;
assign idx_between_23_24_comb_right = index_lt_24_out;
assign idx_between_14_30_reg_write_en = _guard9437;
assign idx_between_14_30_reg_clk = clk;
assign idx_between_14_30_reg_reset = reset;
assign idx_between_14_30_reg_in =
  _guard9440 ? 1'd0 :
  _guard9441 ? idx_between_14_30_comb_out :
  'x;
assign idx_between_26_27_comb_left = index_ge_26_out;
assign idx_between_26_27_comb_right = index_lt_27_out;
assign index_ge_18_left = idx_add_out;
assign index_ge_18_right = 6'd18;
assign idx_between_18_22_comb_left = index_ge_18_out;
assign idx_between_18_22_comb_right = index_lt_22_out;
assign idx_between_23_39_reg_write_en = _guard9452;
assign idx_between_23_39_reg_clk = clk;
assign idx_between_23_39_reg_reset = reset;
assign idx_between_23_39_reg_in =
  _guard9453 ? idx_between_23_39_comb_out :
  _guard9456 ? 1'd0 :
  'x;
assign cond18_write_en = _guard9457;
assign cond18_clk = clk;
assign cond18_reset = reset;
assign cond18_in =
  _guard9458 ? idx_between_24_25_reg_out :
  1'd0;
assign cond_wire24_in =
  _guard9459 ? idx_between_5_21_reg_out :
  _guard9462 ? cond24_out :
  1'd0;
assign cond_wire31_in =
  _guard9463 ? idx_between_7_23_reg_out :
  _guard9466 ? cond31_out :
  1'd0;
assign cond_wire46_in =
  _guard9469 ? cond46_out :
  _guard9470 ? idx_between_10_26_reg_out :
  1'd0;
assign cond_wire48_in =
  _guard9473 ? cond48_out :
  _guard9474 ? idx_between_30_31_reg_out :
  1'd0;
assign cond_wire72_in =
  _guard9477 ? cond72_out :
  _guard9478 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire76_in =
  _guard9479 ? idx_between_16_32_reg_out :
  _guard9482 ? cond76_out :
  1'd0;
assign cond_wire100_in =
  _guard9485 ? cond100_out :
  _guard9486 ? idx_between_7_11_reg_out :
  1'd0;
assign cond105_write_en = _guard9487;
assign cond105_clk = clk;
assign cond105_reset = reset;
assign cond105_in =
  _guard9488 ? idx_between_8_24_reg_out :
  1'd0;
assign cond_wire134_in =
  _guard9491 ? cond134_out :
  _guard9492 ? idx_between_19_35_reg_out :
  1'd0;
assign cond146_write_en = _guard9493;
assign cond146_clk = clk;
assign cond146_reset = reset;
assign cond146_in =
  _guard9494 ? idx_between_3_19_reg_out :
  1'd0;
assign cond_wire146_in =
  _guard9495 ? idx_between_3_19_reg_out :
  _guard9498 ? cond146_out :
  1'd0;
assign cond151_write_en = _guard9499;
assign cond151_clk = clk;
assign cond151_reset = reset;
assign cond151_in =
  _guard9500 ? idx_between_8_24_reg_out :
  1'd0;
assign cond_wire157_in =
  _guard9501 ? idx_between_6_10_reg_out :
  _guard9504 ? cond157_out :
  1'd0;
assign cond_wire167_in =
  _guard9507 ? cond167_out :
  _guard9508 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire174_in =
  _guard9511 ? cond174_out :
  _guard9512 ? idx_between_10_26_reg_out :
  1'd0;
assign cond177_write_en = _guard9513;
assign cond177_clk = clk;
assign cond177_reset = reset;
assign cond177_in =
  _guard9514 ? idx_between_11_15_reg_out :
  1'd0;
assign cond178_write_en = _guard9515;
assign cond178_clk = clk;
assign cond178_reset = reset;
assign cond178_in =
  _guard9516 ? idx_between_11_27_reg_out :
  1'd0;
assign cond_wire191_in =
  _guard9517 ? idx_between_18_34_reg_out :
  _guard9520 ? cond191_out :
  1'd0;
assign cond_wire198_in =
  _guard9521 ? idx_between_16_32_reg_out :
  _guard9524 ? cond198_out :
  1'd0;
assign cond204_write_en = _guard9525;
assign cond204_clk = clk;
assign cond204_reset = reset;
assign cond204_in =
  _guard9526 ? idx_between_37_38_reg_out :
  1'd0;
assign cond215_write_en = _guard9527;
assign cond215_clk = clk;
assign cond215_reset = reset;
assign cond215_in =
  _guard9528 ? idx_between_5_21_reg_out :
  1'd0;
assign cond_wire216_in =
  _guard9531 ? cond216_out :
  _guard9532 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire228_in =
  _guard9535 ? cond228_out :
  _guard9536 ? idx_between_12_28_reg_out :
  1'd0;
assign cond231_write_en = _guard9537;
assign cond231_clk = clk;
assign cond231_reset = reset;
assign cond231_in =
  _guard9538 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire231_in =
  _guard9541 ? cond231_out :
  _guard9542 ? idx_between_9_25_reg_out :
  1'd0;
assign cond237_write_en = _guard9543;
assign cond237_clk = clk;
assign cond237_reset = reset;
assign cond237_in =
  _guard9544 ? idx_between_30_31_reg_out :
  1'd0;
assign cond270_write_en = _guard9545;
assign cond270_clk = clk;
assign cond270_reset = reset;
assign cond270_in =
  _guard9546 ? idx_between_19_23_reg_out :
  1'd0;
assign cond288_write_en = _guard9547;
assign cond288_clk = clk;
assign cond288_reset = reset;
assign cond288_in =
  _guard9548 ? idx_between_8_24_reg_out :
  1'd0;
assign cond302_write_en = _guard9549;
assign cond302_clk = clk;
assign cond302_reset = reset;
assign cond302_in =
  _guard9550 ? idx_between_31_32_reg_out :
  1'd0;
assign cond_wire308_in =
  _guard9551 ? idx_between_13_29_reg_out :
  _guard9554 ? cond308_out :
  1'd0;
assign cond325_write_en = _guard9555;
assign cond325_clk = clk;
assign cond325_reset = reset;
assign cond325_in =
  _guard9556 ? idx_between_21_37_reg_out :
  1'd0;
assign cond349_write_en = _guard9557;
assign cond349_clk = clk;
assign cond349_reset = reset;
assign cond349_in =
  _guard9558 ? idx_between_8_24_reg_out :
  1'd0;
assign cond352_write_en = _guard9559;
assign cond352_clk = clk;
assign cond352_reset = reset;
assign cond352_in =
  _guard9560 ? idx_between_9_13_reg_out :
  1'd0;
assign cond372_write_en = _guard9561;
assign cond372_clk = clk;
assign cond372_reset = reset;
assign cond372_in =
  _guard9562 ? idx_between_14_18_reg_out :
  1'd0;
assign cond_wire372_in =
  _guard9565 ? cond372_out :
  _guard9566 ? idx_between_14_18_reg_out :
  1'd0;
assign cond_wire375_in =
  _guard9567 ? idx_between_34_35_reg_out :
  _guard9570 ? cond375_out :
  1'd0;
assign cond376_write_en = _guard9571;
assign cond376_clk = clk;
assign cond376_reset = reset;
assign cond376_in =
  _guard9572 ? idx_between_15_19_reg_out :
  1'd0;
assign cond_wire376_in =
  _guard9573 ? idx_between_15_19_reg_out :
  _guard9576 ? cond376_out :
  1'd0;
assign cond394_write_en = _guard9577;
assign cond394_clk = clk;
assign cond394_reset = reset;
assign cond394_in =
  _guard9578 ? idx_between_23_39_reg_out :
  1'd0;
assign cond395_write_en = _guard9579;
assign cond395_clk = clk;
assign cond395_reset = reset;
assign cond395_in =
  _guard9580 ? idx_between_39_40_reg_out :
  1'd0;
assign cond_wire405_in =
  _guard9581 ? idx_between_7_11_reg_out :
  _guard9584 ? cond405_out :
  1'd0;
assign cond406_write_en = _guard9585;
assign cond406_clk = clk;
assign cond406_reset = reset;
assign cond406_in =
  _guard9586 ? idx_between_7_23_reg_out :
  1'd0;
assign cond_wire408_in =
  _guard9589 ? cond408_out :
  _guard9590 ? idx_between_27_28_reg_out :
  1'd0;
assign cond_wire457_in =
  _guard9593 ? cond457_out :
  _guard9594 ? idx_between_20_24_reg_out :
  1'd0;
assign cond_wire460_in =
  _guard9597 ? cond460_out :
  _guard9598 ? idx_between_40_41_reg_out :
  1'd0;
assign cond_wire463_in =
  _guard9601 ? cond463_out :
  _guard9602 ? idx_between_25_41_reg_out :
  1'd0;
assign cond465_write_en = _guard9603;
assign cond465_clk = clk;
assign cond465_reset = reset;
assign cond465_in =
  _guard9604 ? idx_between_22_26_reg_out :
  1'd0;
assign cond_wire477_in =
  _guard9605 ? idx_between_29_30_reg_out :
  _guard9608 ? cond477_out :
  1'd0;
assign cond_wire535_in =
  _guard9609 ? idx_between_9_13_reg_out :
  _guard9612 ? cond535_out :
  1'd0;
assign cond542_write_en = _guard9613;
assign cond542_clk = clk;
assign cond542_reset = reset;
assign cond542_in =
  _guard9614 ? idx_between_30_31_reg_out :
  1'd0;
assign cond_wire547_in =
  _guard9617 ? cond547_out :
  _guard9618 ? idx_between_12_16_reg_out :
  1'd0;
assign cond_wire550_in =
  _guard9619 ? idx_between_32_33_reg_out :
  _guard9622 ? cond550_out :
  1'd0;
assign cond_wire553_in =
  _guard9623 ? idx_between_17_33_reg_out :
  _guard9626 ? cond553_out :
  1'd0;
assign cond_wire563_in =
  _guard9627 ? idx_between_16_20_reg_out :
  _guard9630 ? cond563_out :
  1'd0;
assign cond_wire565_in =
  _guard9631 ? idx_between_20_36_reg_out :
  _guard9634 ? cond565_out :
  1'd0;
assign cond_wire587_in =
  _guard9637 ? cond587_out :
  _guard9638 ? idx_between_22_26_reg_out :
  1'd0;
assign cond600_write_en = _guard9639;
assign cond600_clk = clk;
assign cond600_reset = reset;
assign cond600_in =
  _guard9640 ? idx_between_10_14_reg_out :
  1'd0;
assign cond602_write_en = _guard9641;
assign cond602_clk = clk;
assign cond602_reset = reset;
assign cond602_in =
  _guard9642 ? idx_between_14_30_reg_out :
  1'd0;
assign cond_wire607_in =
  _guard9643 ? idx_between_31_32_reg_out :
  _guard9646 ? cond607_out :
  1'd0;
assign cond_wire609_in =
  _guard9647 ? idx_between_12_28_reg_out :
  _guard9650 ? cond609_out :
  1'd0;
assign cond_wire621_in =
  _guard9653 ? cond621_out :
  _guard9654 ? idx_between_15_31_reg_out :
  1'd0;
assign cond628_write_en = _guard9655;
assign cond628_clk = clk;
assign cond628_reset = reset;
assign cond628_in =
  _guard9656 ? idx_between_17_21_reg_out :
  1'd0;
assign cond631_write_en = _guard9657;
assign cond631_clk = clk;
assign cond631_reset = reset;
assign cond631_in =
  _guard9658 ? idx_between_37_38_reg_out :
  1'd0;
assign cond_wire638_in =
  _guard9659 ? idx_between_23_39_reg_out :
  _guard9662 ? cond638_out :
  1'd0;
assign cond647_write_en = _guard9663;
assign cond647_clk = clk;
assign cond647_reset = reset;
assign cond647_in =
  _guard9664 ? idx_between_41_42_reg_out :
  1'd0;
assign cond_wire648_in =
  _guard9667 ? cond648_out :
  _guard9668 ? idx_between_22_26_reg_out :
  1'd0;
assign cond_wire652_in =
  _guard9671 ? cond652_out :
  _guard9672 ? idx_between_23_27_reg_out :
  1'd0;
assign cond_wire655_in =
  _guard9673 ? idx_between_43_44_reg_out :
  _guard9676 ? cond655_out :
  1'd0;
assign cond_wire671_in =
  _guard9677 ? idx_between_16_32_reg_out :
  _guard9680 ? cond671_out :
  1'd0;
assign cond_wire674_in =
  _guard9681 ? idx_between_13_29_reg_out :
  _guard9684 ? cond674_out :
  1'd0;
assign cond675_write_en = _guard9685;
assign cond675_clk = clk;
assign cond675_reset = reset;
assign cond675_in =
  _guard9686 ? idx_between_17_33_reg_out :
  1'd0;
assign cond_wire677_in =
  _guard9687 ? idx_between_14_18_reg_out :
  _guard9690 ? cond677_out :
  1'd0;
assign cond_wire685_in =
  _guard9691 ? idx_between_16_20_reg_out :
  _guard9694 ? cond685_out :
  1'd0;
assign cond693_write_en = _guard9695;
assign cond693_clk = clk;
assign cond693_reset = reset;
assign cond693_in =
  _guard9696 ? idx_between_18_22_reg_out :
  1'd0;
assign cond_wire697_in =
  _guard9697 ? idx_between_19_23_reg_out :
  _guard9700 ? cond697_out :
  1'd0;
assign cond_wire710_in =
  _guard9703 ? cond710_out :
  _guard9704 ? idx_between_22_38_reg_out :
  1'd0;
assign cond716_write_en = _guard9705;
assign cond716_clk = clk;
assign cond716_reset = reset;
assign cond716_in =
  _guard9706 ? idx_between_43_44_reg_out :
  1'd0;
assign cond_wire717_in =
  _guard9707 ? idx_between_24_28_reg_out :
  _guard9710 ? cond717_out :
  1'd0;
assign cond728_write_en = _guard9711;
assign cond728_clk = clk;
assign cond728_reset = reset;
assign cond728_in =
  _guard9712 ? idx_between_46_47_reg_out :
  1'd0;
assign cond729_write_en = _guard9713;
assign cond729_clk = clk;
assign cond729_reset = reset;
assign cond729_in =
  _guard9714 ? idx_between_11_27_reg_out :
  1'd0;
assign cond_wire734_in =
  _guard9717 ? cond734_out :
  _guard9718 ? idx_between_13_17_reg_out :
  1'd0;
assign cond_wire738_in =
  _guard9719 ? idx_between_14_18_reg_out :
  _guard9722 ? cond738_out :
  1'd0;
assign cond_wire761_in =
  _guard9723 ? idx_between_39_40_reg_out :
  _guard9726 ? cond761_out :
  1'd0;
assign cond_wire762_in =
  _guard9729 ? cond762_out :
  _guard9730 ? idx_between_20_24_reg_out :
  1'd0;
assign cond764_write_en = _guard9731;
assign cond764_clk = clk;
assign cond764_reset = reset;
assign cond764_in =
  _guard9732 ? idx_between_24_40_reg_out :
  1'd0;
assign cond766_write_en = _guard9733;
assign cond766_clk = clk;
assign cond766_reset = reset;
assign cond766_in =
  _guard9734 ? idx_between_21_25_reg_out :
  1'd0;
assign cond_wire767_in =
  _guard9737 ? cond767_out :
  _guard9738 ? idx_between_21_37_reg_out :
  1'd0;
assign cond769_write_en = _guard9739;
assign cond769_clk = clk;
assign cond769_reset = reset;
assign cond769_in =
  _guard9740 ? idx_between_41_42_reg_out :
  1'd0;
assign cond_wire774_in =
  _guard9743 ? cond774_out :
  _guard9744 ? idx_between_23_27_reg_out :
  1'd0;
assign cond775_write_en = _guard9745;
assign cond775_clk = clk;
assign cond775_reset = reset;
assign cond775_in =
  _guard9746 ? idx_between_23_39_reg_out :
  1'd0;
assign cond778_write_en = _guard9747;
assign cond778_clk = clk;
assign cond778_reset = reset;
assign cond778_in =
  _guard9748 ? idx_between_24_28_reg_out :
  1'd0;
assign cond_wire780_in =
  _guard9751 ? cond780_out :
  _guard9752 ? idx_between_28_44_reg_out :
  1'd0;
assign cond_wire792_in =
  _guard9755 ? cond792_out :
  _guard9756 ? idx_between_31_47_reg_out :
  1'd0;
assign cond797_write_en = _guard9757;
assign cond797_clk = clk;
assign cond797_reset = reset;
assign cond797_in =
  _guard9758 ? idx_between_17_33_reg_out :
  1'd0;
assign cond_wire801_in =
  _guard9759 ? idx_between_18_34_reg_out :
  _guard9762 ? cond801_out :
  1'd0;
assign cond_wire802_in =
  _guard9763 ? idx_between_34_35_reg_out :
  _guard9766 ? cond802_out :
  1'd0;
assign cond_wire806_in =
  _guard9769 ? cond806_out :
  _guard9770 ? idx_between_35_36_reg_out :
  1'd0;
assign cond_wire807_in =
  _guard9771 ? idx_between_16_20_reg_out :
  _guard9774 ? cond807_out :
  1'd0;
assign cond808_write_en = _guard9775;
assign cond808_clk = clk;
assign cond808_reset = reset;
assign cond808_in =
  _guard9776 ? idx_between_16_32_reg_out :
  1'd0;
assign cond811_write_en = _guard9777;
assign cond811_clk = clk;
assign cond811_reset = reset;
assign cond811_in =
  _guard9778 ? idx_between_17_21_reg_out :
  1'd0;
assign cond_wire814_in =
  _guard9781 ? cond814_out :
  _guard9782 ? idx_between_37_38_reg_out :
  1'd0;
assign cond_wire818_in =
  _guard9785 ? cond818_out :
  _guard9786 ? idx_between_38_39_reg_out :
  1'd0;
assign cond_wire829_in =
  _guard9789 ? cond829_out :
  _guard9790 ? idx_between_25_41_reg_out :
  1'd0;
assign cond836_write_en = _guard9791;
assign cond836_clk = clk;
assign cond836_reset = reset;
assign cond836_in =
  _guard9792 ? idx_between_23_39_reg_out :
  1'd0;
assign cond_wire845_in =
  _guard9793 ? idx_between_29_45_reg_out :
  _guard9796 ? cond845_out :
  1'd0;
assign cond_wire859_in =
  _guard9797 ? idx_between_13_29_reg_out :
  _guard9800 ? cond859_out :
  1'd0;
assign cond_wire871_in =
  _guard9801 ? idx_between_36_37_reg_out :
  _guard9804 ? cond871_out :
  1'd0;
assign cond_wire878_in =
  _guard9807 ? cond878_out :
  _guard9808 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire889_in =
  _guard9811 ? cond889_out :
  _guard9812 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire904_in =
  _guard9813 ? idx_between_25_29_reg_out :
  _guard9816 ? cond904_out :
  1'd0;
assign cond_wire906_in =
  _guard9817 ? idx_between_29_45_reg_out :
  _guard9820 ? cond906_out :
  1'd0;
assign cond916_write_en = _guard9821;
assign cond916_clk = clk;
assign cond916_reset = reset;
assign cond916_in =
  _guard9822 ? idx_between_28_32_reg_out :
  1'd0;
assign cond917_write_en = _guard9823;
assign cond917_clk = clk;
assign cond917_reset = reset;
assign cond917_in =
  _guard9824 ? idx_between_28_44_reg_out :
  1'd0;
assign cond919_write_en = _guard9825;
assign cond919_clk = clk;
assign cond919_reset = reset;
assign cond919_in =
  _guard9826 ? idx_between_48_49_reg_out :
  1'd0;
assign cond_wire919_in =
  _guard9829 ? cond919_out :
  _guard9830 ? idx_between_48_49_reg_out :
  1'd0;
assign cond931_write_en = _guard9831;
assign cond931_clk = clk;
assign cond931_reset = reset;
assign cond931_in =
  _guard9832 ? idx_between_20_36_reg_out :
  1'd0;
assign cond947_write_en = _guard9833;
assign cond947_clk = clk;
assign cond947_reset = reset;
assign cond947_in =
  _guard9834 ? idx_between_24_40_reg_out :
  1'd0;
assign cond953_write_en = _guard9835;
assign cond953_clk = clk;
assign cond953_reset = reset;
assign cond953_in =
  _guard9836 ? idx_between_22_26_reg_out :
  1'd0;
assign cond967_write_en = _guard9837;
assign cond967_clk = clk;
assign cond967_reset = reset;
assign cond967_in =
  _guard9838 ? idx_between_29_45_reg_out :
  1'd0;
assign cond_wire968_in =
  _guard9841 ? cond968_out :
  _guard9842 ? idx_between_45_46_reg_out :
  1'd0;
assign cond985_write_en = _guard9843;
assign cond985_clk = clk;
assign cond985_reset = reset;
assign cond985_in =
  _guard9844 ? idx_between_30_34_reg_out :
  1'd0;
assign cond1017_write_en = _guard9845;
assign cond1017_clk = clk;
assign cond1017_reset = reset;
assign cond1017_in =
  _guard9846 ? idx_between_42_43_reg_out :
  1'd0;
assign cond_wire1018_in =
  _guard9849 ? cond1018_out :
  _guard9850 ? idx_between_23_27_reg_out :
  1'd0;
assign cond_wire1023_in =
  _guard9853 ? cond1023_out :
  _guard9854 ? idx_between_24_40_reg_out :
  1'd0;
assign cond1034_write_en = _guard9855;
assign cond1034_clk = clk;
assign cond1034_reset = reset;
assign cond1034_in =
  _guard9856 ? idx_between_27_31_reg_out :
  1'd0;
assign cond1038_write_en = _guard9857;
assign cond1038_clk = clk;
assign cond1038_reset = reset;
assign cond1038_in =
  _guard9858 ? idx_between_28_32_reg_out :
  1'd0;
assign cond1039_write_en = _guard9859;
assign cond1039_clk = clk;
assign cond1039_reset = reset;
assign cond1039_in =
  _guard9860 ? idx_between_28_44_reg_out :
  1'd0;
assign cond_wire1043_in =
  _guard9861 ? idx_between_29_45_reg_out :
  _guard9864 ? cond1043_out :
  1'd0;
assign left_0_0_write_en = _guard9867;
assign left_0_0_clk = clk;
assign left_0_0_reset = reset;
assign left_0_0_in = l0_read_data;
assign pe_0_3_mul_ready =
  _guard9873 ? 1'd1 :
  _guard9876 ? 1'd0 :
  1'd0;
assign pe_0_3_clk = clk;
assign pe_0_3_top =
  _guard9889 ? top_0_3_out :
  32'd0;
assign pe_0_3_left =
  _guard9902 ? left_0_3_out :
  32'd0;
assign pe_0_3_reset = reset;
assign pe_0_3_go = _guard9915;
assign pe_0_5_mul_ready =
  _guard9918 ? 1'd1 :
  _guard9921 ? 1'd0 :
  1'd0;
assign pe_0_5_clk = clk;
assign pe_0_5_top =
  _guard9934 ? top_0_5_out :
  32'd0;
assign pe_0_5_left =
  _guard9947 ? left_0_5_out :
  32'd0;
assign pe_0_5_reset = reset;
assign pe_0_5_go = _guard9960;
assign pe_0_8_mul_ready =
  _guard9963 ? 1'd1 :
  _guard9966 ? 1'd0 :
  1'd0;
assign pe_0_8_clk = clk;
assign pe_0_8_top =
  _guard9979 ? top_0_8_out :
  32'd0;
assign pe_0_8_left =
  _guard9992 ? left_0_8_out :
  32'd0;
assign pe_0_8_reset = reset;
assign pe_0_8_go = _guard10005;
assign pe_0_9_mul_ready =
  _guard10008 ? 1'd1 :
  _guard10011 ? 1'd0 :
  1'd0;
assign pe_0_9_clk = clk;
assign pe_0_9_top =
  _guard10024 ? top_0_9_out :
  32'd0;
assign pe_0_9_left =
  _guard10037 ? left_0_9_out :
  32'd0;
assign pe_0_9_reset = reset;
assign pe_0_9_go = _guard10050;
assign top_0_12_write_en = _guard10053;
assign top_0_12_clk = clk;
assign top_0_12_reset = reset;
assign top_0_12_in = t12_read_data;
assign top_1_3_write_en = _guard10059;
assign top_1_3_clk = clk;
assign top_1_3_reset = reset;
assign top_1_3_in = top_0_3_out;
assign top_1_4_write_en = _guard10065;
assign top_1_4_clk = clk;
assign top_1_4_reset = reset;
assign top_1_4_in = top_0_4_out;
assign top_1_8_write_en = _guard10071;
assign top_1_8_clk = clk;
assign top_1_8_reset = reset;
assign top_1_8_in = top_0_8_out;
assign left_2_3_write_en = _guard10077;
assign left_2_3_clk = clk;
assign left_2_3_reset = reset;
assign left_2_3_in = left_2_2_out;
assign pe_2_4_mul_ready =
  _guard10083 ? 1'd1 :
  _guard10086 ? 1'd0 :
  1'd0;
assign pe_2_4_clk = clk;
assign pe_2_4_top =
  _guard10099 ? top_2_4_out :
  32'd0;
assign pe_2_4_left =
  _guard10112 ? left_2_4_out :
  32'd0;
assign pe_2_4_reset = reset;
assign pe_2_4_go = _guard10125;
assign top_2_6_write_en = _guard10128;
assign top_2_6_clk = clk;
assign top_2_6_reset = reset;
assign top_2_6_in = top_1_6_out;
assign top_2_11_write_en = _guard10134;
assign top_2_11_clk = clk;
assign top_2_11_reset = reset;
assign top_2_11_in = top_1_11_out;
assign pe_2_15_mul_ready =
  _guard10140 ? 1'd1 :
  _guard10143 ? 1'd0 :
  1'd0;
assign pe_2_15_clk = clk;
assign pe_2_15_top =
  _guard10156 ? top_2_15_out :
  32'd0;
assign pe_2_15_left =
  _guard10169 ? left_2_15_out :
  32'd0;
assign pe_2_15_reset = reset;
assign pe_2_15_go = _guard10182;
assign pe_3_0_mul_ready =
  _guard10185 ? 1'd1 :
  _guard10188 ? 1'd0 :
  1'd0;
assign pe_3_0_clk = clk;
assign pe_3_0_top =
  _guard10201 ? top_3_0_out :
  32'd0;
assign pe_3_0_left =
  _guard10214 ? left_3_0_out :
  32'd0;
assign pe_3_0_reset = reset;
assign pe_3_0_go = _guard10227;
assign top_3_2_write_en = _guard10230;
assign top_3_2_clk = clk;
assign top_3_2_reset = reset;
assign top_3_2_in = top_2_2_out;
assign top_3_14_write_en = _guard10236;
assign top_3_14_clk = clk;
assign top_3_14_reset = reset;
assign top_3_14_in = top_2_14_out;
assign top_4_0_write_en = _guard10242;
assign top_4_0_clk = clk;
assign top_4_0_reset = reset;
assign top_4_0_in = top_3_0_out;
assign left_4_6_write_en = _guard10248;
assign left_4_6_clk = clk;
assign left_4_6_reset = reset;
assign left_4_6_in = left_4_5_out;
assign left_4_7_write_en = _guard10254;
assign left_4_7_clk = clk;
assign left_4_7_reset = reset;
assign left_4_7_in = left_4_6_out;
assign pe_5_1_mul_ready =
  _guard10260 ? 1'd1 :
  _guard10263 ? 1'd0 :
  1'd0;
assign pe_5_1_clk = clk;
assign pe_5_1_top =
  _guard10276 ? top_5_1_out :
  32'd0;
assign pe_5_1_left =
  _guard10289 ? left_5_1_out :
  32'd0;
assign pe_5_1_reset = reset;
assign pe_5_1_go = _guard10302;
assign pe_5_7_mul_ready =
  _guard10305 ? 1'd1 :
  _guard10308 ? 1'd0 :
  1'd0;
assign pe_5_7_clk = clk;
assign pe_5_7_top =
  _guard10321 ? top_5_7_out :
  32'd0;
assign pe_5_7_left =
  _guard10334 ? left_5_7_out :
  32'd0;
assign pe_5_7_reset = reset;
assign pe_5_7_go = _guard10347;
assign pe_6_0_mul_ready =
  _guard10350 ? 1'd1 :
  _guard10353 ? 1'd0 :
  1'd0;
assign pe_6_0_clk = clk;
assign pe_6_0_top =
  _guard10366 ? top_6_0_out :
  32'd0;
assign pe_6_0_left =
  _guard10379 ? left_6_0_out :
  32'd0;
assign pe_6_0_reset = reset;
assign pe_6_0_go = _guard10392;
assign top_6_0_write_en = _guard10395;
assign top_6_0_clk = clk;
assign top_6_0_reset = reset;
assign top_6_0_in = top_5_0_out;
assign pe_6_1_mul_ready =
  _guard10401 ? 1'd1 :
  _guard10404 ? 1'd0 :
  1'd0;
assign pe_6_1_clk = clk;
assign pe_6_1_top =
  _guard10417 ? top_6_1_out :
  32'd0;
assign pe_6_1_left =
  _guard10430 ? left_6_1_out :
  32'd0;
assign pe_6_1_reset = reset;
assign pe_6_1_go = _guard10443;
assign left_6_11_write_en = _guard10446;
assign left_6_11_clk = clk;
assign left_6_11_reset = reset;
assign left_6_11_in = left_6_10_out;
assign left_7_5_write_en = _guard10452;
assign left_7_5_clk = clk;
assign left_7_5_reset = reset;
assign left_7_5_in = left_7_4_out;
assign pe_8_2_mul_ready =
  _guard10458 ? 1'd1 :
  _guard10461 ? 1'd0 :
  1'd0;
assign pe_8_2_clk = clk;
assign pe_8_2_top =
  _guard10474 ? top_8_2_out :
  32'd0;
assign pe_8_2_left =
  _guard10487 ? left_8_2_out :
  32'd0;
assign pe_8_2_reset = reset;
assign pe_8_2_go = _guard10500;
assign top_8_3_write_en = _guard10503;
assign top_8_3_clk = clk;
assign top_8_3_reset = reset;
assign top_8_3_in = top_7_3_out;
assign pe_8_4_mul_ready =
  _guard10509 ? 1'd1 :
  _guard10512 ? 1'd0 :
  1'd0;
assign pe_8_4_clk = clk;
assign pe_8_4_top =
  _guard10525 ? top_8_4_out :
  32'd0;
assign pe_8_4_left =
  _guard10538 ? left_8_4_out :
  32'd0;
assign pe_8_4_reset = reset;
assign pe_8_4_go = _guard10551;
assign top_10_6_write_en = _guard10554;
assign top_10_6_clk = clk;
assign top_10_6_reset = reset;
assign top_10_6_in = top_9_6_out;
assign left_10_9_write_en = _guard10560;
assign left_10_9_clk = clk;
assign left_10_9_reset = reset;
assign left_10_9_in = left_10_8_out;
assign pe_11_0_mul_ready =
  _guard10566 ? 1'd1 :
  _guard10569 ? 1'd0 :
  1'd0;
assign pe_11_0_clk = clk;
assign pe_11_0_top =
  _guard10582 ? top_11_0_out :
  32'd0;
assign pe_11_0_left =
  _guard10595 ? left_11_0_out :
  32'd0;
assign pe_11_0_reset = reset;
assign pe_11_0_go = _guard10608;
assign top_11_3_write_en = _guard10611;
assign top_11_3_clk = clk;
assign top_11_3_reset = reset;
assign top_11_3_in = top_10_3_out;
assign top_11_5_write_en = _guard10617;
assign top_11_5_clk = clk;
assign top_11_5_reset = reset;
assign top_11_5_in = top_10_5_out;
assign pe_11_11_mul_ready =
  _guard10623 ? 1'd1 :
  _guard10626 ? 1'd0 :
  1'd0;
assign pe_11_11_clk = clk;
assign pe_11_11_top =
  _guard10639 ? top_11_11_out :
  32'd0;
assign pe_11_11_left =
  _guard10652 ? left_11_11_out :
  32'd0;
assign pe_11_11_reset = reset;
assign pe_11_11_go = _guard10665;
assign left_11_15_write_en = _guard10668;
assign left_11_15_clk = clk;
assign left_11_15_reset = reset;
assign left_11_15_in = left_11_14_out;
assign top_12_0_write_en = _guard10674;
assign top_12_0_clk = clk;
assign top_12_0_reset = reset;
assign top_12_0_in = top_11_0_out;
assign top_12_2_write_en = _guard10680;
assign top_12_2_clk = clk;
assign top_12_2_reset = reset;
assign top_12_2_in = top_11_2_out;
assign top_12_7_write_en = _guard10686;
assign top_12_7_clk = clk;
assign top_12_7_reset = reset;
assign top_12_7_in = top_11_7_out;
assign left_12_8_write_en = _guard10692;
assign left_12_8_clk = clk;
assign left_12_8_reset = reset;
assign left_12_8_in = left_12_7_out;
assign top_13_4_write_en = _guard10698;
assign top_13_4_clk = clk;
assign top_13_4_reset = reset;
assign top_13_4_in = top_12_4_out;
assign top_13_9_write_en = _guard10704;
assign top_13_9_clk = clk;
assign top_13_9_reset = reset;
assign top_13_9_in = top_12_9_out;
assign top_13_15_write_en = _guard10710;
assign top_13_15_clk = clk;
assign top_13_15_reset = reset;
assign top_13_15_in = top_12_15_out;
assign top_14_8_write_en = _guard10716;
assign top_14_8_clk = clk;
assign top_14_8_reset = reset;
assign top_14_8_in = top_13_8_out;
assign top_15_4_write_en = _guard10722;
assign top_15_4_clk = clk;
assign top_15_4_reset = reset;
assign top_15_4_in = top_14_4_out;
assign left_15_10_write_en = _guard10728;
assign left_15_10_clk = clk;
assign left_15_10_reset = reset;
assign left_15_10_in = left_15_9_out;
assign l11_add_left = 5'd1;
assign l11_add_right = l11_idx_out;
assign index_lt_30_left = idx_add_out;
assign index_lt_30_right = 6'd30;
assign index_ge_25_left = idx_add_out;
assign index_ge_25_right = 6'd25;
assign idx_between_17_21_reg_write_en = _guard10746;
assign idx_between_17_21_reg_clk = clk;
assign idx_between_17_21_reg_reset = reset;
assign idx_between_17_21_reg_in =
  _guard10747 ? idx_between_17_21_comb_out :
  _guard10750 ? 1'd0 :
  'x;
assign index_lt_27_left = idx_add_out;
assign index_lt_27_right = 6'd27;
assign index_ge_20_left = idx_add_out;
assign index_ge_20_right = 6'd20;
assign idx_between_29_45_reg_write_en = _guard10759;
assign idx_between_29_45_reg_clk = clk;
assign idx_between_29_45_reg_reset = reset;
assign idx_between_29_45_reg_in =
  _guard10760 ? idx_between_29_45_comb_out :
  _guard10763 ? 1'd0 :
  'x;
assign idx_between_22_23_reg_write_en = _guard10768;
assign idx_between_22_23_reg_clk = clk;
assign idx_between_22_23_reg_reset = reset;
assign idx_between_22_23_reg_in =
  _guard10771 ? 1'd0 :
  _guard10772 ? idx_between_22_23_comb_out :
  'x;
assign idx_between_21_25_reg_write_en = _guard10777;
assign idx_between_21_25_reg_clk = clk;
assign idx_between_21_25_reg_reset = reset;
assign idx_between_21_25_reg_in =
  _guard10778 ? idx_between_21_25_comb_out :
  _guard10781 ? 1'd0 :
  'x;
assign idx_between_49_50_comb_left = index_ge_49_out;
assign idx_between_49_50_comb_right = index_lt_50_out;
assign idx_between_6_22_comb_left = index_ge_6_out;
assign idx_between_6_22_comb_right = index_lt_22_out;
assign idx_between_11_27_comb_left = index_ge_11_out;
assign idx_between_11_27_comb_right = index_lt_27_out;
assign idx_between_21_22_reg_write_en = _guard10792;
assign idx_between_21_22_reg_clk = clk;
assign idx_between_21_22_reg_reset = reset;
assign idx_between_21_22_reg_in =
  _guard10793 ? idx_between_21_22_comb_out :
  _guard10796 ? 1'd0 :
  'x;
assign idx_between_31_32_comb_left = index_ge_31_out;
assign idx_between_31_32_comb_right = index_lt_32_out;
assign idx_between_14_18_comb_left = index_ge_14_out;
assign idx_between_14_18_comb_right = index_lt_18_out;
assign idx_between_36_37_reg_write_en = _guard10805;
assign idx_between_36_37_reg_clk = clk;
assign idx_between_36_37_reg_reset = reset;
assign idx_between_36_37_reg_in =
  _guard10808 ? 1'd0 :
  _guard10809 ? idx_between_36_37_comb_out :
  'x;
assign idx_between_28_44_comb_left = index_ge_28_out;
assign idx_between_28_44_comb_right = index_lt_44_out;
assign idx_between_15_19_comb_left = index_ge_15_out;
assign idx_between_15_19_comb_right = index_lt_19_out;
assign idx_between_20_36_reg_write_en = _guard10818;
assign idx_between_20_36_reg_clk = clk;
assign idx_between_20_36_reg_reset = reset;
assign idx_between_20_36_reg_in =
  _guard10819 ? idx_between_20_36_comb_out :
  _guard10822 ? 1'd0 :
  'x;
assign idx_between_20_36_comb_left = index_ge_20_out;
assign idx_between_20_36_comb_right = index_lt_36_out;
assign cond_wire18_in =
  _guard10827 ? cond18_out :
  _guard10828 ? idx_between_24_25_reg_out :
  1'd0;
assign cond19_write_en = _guard10829;
assign cond19_clk = clk;
assign cond19_reset = reset;
assign cond19_in =
  _guard10830 ? idx_between_4_20_reg_out :
  1'd0;
assign cond_wire29_in =
  _guard10831 ? idx_between_6_22_reg_out :
  _guard10834 ? cond29_out :
  1'd0;
assign cond34_write_en = _guard10835;
assign cond34_clk = clk;
assign cond34_reset = reset;
assign cond34_in =
  _guard10836 ? idx_between_7_23_reg_out :
  1'd0;
assign cond40_write_en = _guard10837;
assign cond40_clk = clk;
assign cond40_reset = reset;
assign cond40_in =
  _guard10838 ? idx_between_9_13_reg_out :
  1'd0;
assign cond57_write_en = _guard10839;
assign cond57_clk = clk;
assign cond57_reset = reset;
assign cond57_in =
  _guard10840 ? idx_between_16_32_reg_out :
  1'd0;
assign cond_wire59_in =
  _guard10841 ? idx_between_12_28_reg_out :
  _guard10844 ? cond59_out :
  1'd0;
assign cond_wire61_in =
  _guard10845 ? idx_between_13_29_reg_out :
  _guard10848 ? cond61_out :
  1'd0;
assign cond74_write_en = _guard10849;
assign cond74_clk = clk;
assign cond74_reset = reset;
assign cond74_in =
  _guard10850 ? idx_between_15_31_reg_out :
  1'd0;
assign cond95_write_en = _guard10851;
assign cond95_clk = clk;
assign cond95_reset = reset;
assign cond95_in =
  _guard10852 ? idx_between_25_26_reg_out :
  1'd0;
assign cond109_write_en = _guard10853;
assign cond109_clk = clk;
assign cond109_reset = reset;
assign cond109_in =
  _guard10854 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire111_in =
  _guard10855 ? idx_between_29_30_reg_out :
  _guard10858 ? cond111_out :
  1'd0;
assign cond_wire112_in =
  _guard10861 ? cond112_out :
  _guard10862 ? idx_between_10_14_reg_out :
  1'd0;
assign cond_wire118_in =
  _guard10865 ? cond118_out :
  _guard10866 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire137_in =
  _guard10867 ? idx_between_16_32_reg_out :
  _guard10870 ? cond137_out :
  1'd0;
assign cond158_write_en = _guard10871;
assign cond158_clk = clk;
assign cond158_reset = reset;
assign cond158_in =
  _guard10872 ? idx_between_6_22_reg_out :
  1'd0;
assign cond159_write_en = _guard10873;
assign cond159_clk = clk;
assign cond159_reset = reset;
assign cond159_in =
  _guard10874 ? idx_between_10_26_reg_out :
  1'd0;
assign cond162_write_en = _guard10875;
assign cond162_clk = clk;
assign cond162_reset = reset;
assign cond162_in =
  _guard10876 ? idx_between_7_23_reg_out :
  1'd0;
assign cond164_write_en = _guard10877;
assign cond164_clk = clk;
assign cond164_reset = reset;
assign cond164_in =
  _guard10878 ? idx_between_27_28_reg_out :
  1'd0;
assign cond166_write_en = _guard10879;
assign cond166_clk = clk;
assign cond166_reset = reset;
assign cond166_in =
  _guard10880 ? idx_between_8_24_reg_out :
  1'd0;
assign cond_wire170_in =
  _guard10883 ? cond170_out :
  _guard10884 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire175_in =
  _guard10885 ? idx_between_14_30_reg_out :
  _guard10888 ? cond175_out :
  1'd0;
assign cond180_write_en = _guard10889;
assign cond180_clk = clk;
assign cond180_reset = reset;
assign cond180_in =
  _guard10890 ? idx_between_31_32_reg_out :
  1'd0;
assign cond_wire197_in =
  _guard10891 ? idx_between_16_20_reg_out :
  _guard10894 ? cond197_out :
  1'd0;
assign cond198_write_en = _guard10895;
assign cond198_clk = clk;
assign cond198_reset = reset;
assign cond198_in =
  _guard10896 ? idx_between_16_32_reg_out :
  1'd0;
assign cond217_write_en = _guard10897;
assign cond217_clk = clk;
assign cond217_reset = reset;
assign cond217_in =
  _guard10898 ? idx_between_25_26_reg_out :
  1'd0;
assign cond222_write_en = _guard10899;
assign cond222_clk = clk;
assign cond222_reset = reset;
assign cond222_in =
  _guard10900 ? idx_between_7_11_reg_out :
  1'd0;
assign cond_wire222_in =
  _guard10901 ? idx_between_7_11_reg_out :
  _guard10904 ? cond222_out :
  1'd0;
assign cond_wire223_in =
  _guard10905 ? idx_between_7_23_reg_out :
  _guard10908 ? cond223_out :
  1'd0;
assign cond_wire225_in =
  _guard10909 ? idx_between_27_28_reg_out :
  _guard10912 ? cond225_out :
  1'd0;
assign cond_wire237_in =
  _guard10915 ? cond237_out :
  _guard10916 ? idx_between_30_31_reg_out :
  1'd0;
assign cond247_write_en = _guard10917;
assign cond247_clk = clk;
assign cond247_reset = reset;
assign cond247_in =
  _guard10918 ? idx_between_13_29_reg_out :
  1'd0;
assign cond_wire260_in =
  _guard10919 ? idx_between_20_36_reg_out :
  _guard10922 ? cond260_out :
  1'd0;
assign cond_wire284_in =
  _guard10923 ? idx_between_7_23_reg_out :
  _guard10926 ? cond284_out :
  1'd0;
assign cond289_write_en = _guard10927;
assign cond289_clk = clk;
assign cond289_reset = reset;
assign cond289_in =
  _guard10928 ? idx_between_12_28_reg_out :
  1'd0;
assign cond293_write_en = _guard10929;
assign cond293_clk = clk;
assign cond293_reset = reset;
assign cond293_in =
  _guard10930 ? idx_between_13_29_reg_out :
  1'd0;
assign cond_wire296_in =
  _guard10933 ? cond296_out :
  _guard10934 ? idx_between_10_26_reg_out :
  1'd0;
assign cond297_write_en = _guard10935;
assign cond297_clk = clk;
assign cond297_reset = reset;
assign cond297_in =
  _guard10936 ? idx_between_14_30_reg_out :
  1'd0;
assign cond_wire317_in =
  _guard10939 ? cond317_out :
  _guard10940 ? idx_between_19_35_reg_out :
  1'd0;
assign cond322_write_en = _guard10941;
assign cond322_clk = clk;
assign cond322_reset = reset;
assign cond322_in =
  _guard10942 ? idx_between_36_37_reg_out :
  1'd0;
assign cond_wire327_in =
  _guard10943 ? idx_between_18_22_reg_out :
  _guard10946 ? cond327_out :
  1'd0;
assign cond_wire329_in =
  _guard10949 ? cond329_out :
  _guard10950 ? idx_between_22_38_reg_out :
  1'd0;
assign cond336_write_en = _guard10951;
assign cond336_clk = clk;
assign cond336_reset = reset;
assign cond336_in =
  _guard10952 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire344_in =
  _guard10953 ? idx_between_7_11_reg_out :
  _guard10956 ? cond344_out :
  1'd0;
assign cond_wire348_in =
  _guard10957 ? idx_between_8_12_reg_out :
  _guard10960 ? cond348_out :
  1'd0;
assign cond355_write_en = _guard10961;
assign cond355_clk = clk;
assign cond355_reset = reset;
assign cond355_in =
  _guard10962 ? idx_between_29_30_reg_out :
  1'd0;
assign cond373_write_en = _guard10963;
assign cond373_clk = clk;
assign cond373_reset = reset;
assign cond373_in =
  _guard10964 ? idx_between_14_30_reg_out :
  1'd0;
assign cond_wire383_in =
  _guard10967 ? cond383_out :
  _guard10968 ? idx_between_36_37_reg_out :
  1'd0;
assign cond388_write_en = _guard10969;
assign cond388_clk = clk;
assign cond388_reset = reset;
assign cond388_in =
  _guard10970 ? idx_between_18_22_reg_out :
  1'd0;
assign cond404_write_en = _guard10971;
assign cond404_clk = clk;
assign cond404_reset = reset;
assign cond404_in =
  _guard10972 ? idx_between_6_22_reg_out :
  1'd0;
assign cond408_write_en = _guard10973;
assign cond408_clk = clk;
assign cond408_reset = reset;
assign cond408_in =
  _guard10974 ? idx_between_27_28_reg_out :
  1'd0;
assign cond412_write_en = _guard10975;
assign cond412_clk = clk;
assign cond412_reset = reset;
assign cond412_in =
  _guard10976 ? idx_between_28_29_reg_out :
  1'd0;
assign cond_wire424_in =
  _guard10979 ? cond424_out :
  _guard10980 ? idx_between_31_32_reg_out :
  1'd0;
assign cond_wire427_in =
  _guard10981 ? idx_between_16_32_reg_out :
  _guard10984 ? cond427_out :
  1'd0;
assign cond438_write_en = _guard10985;
assign cond438_clk = clk;
assign cond438_reset = reset;
assign cond438_in =
  _guard10986 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire438_in =
  _guard10989 ? cond438_out :
  _guard10990 ? idx_between_15_31_reg_out :
  1'd0;
assign cond439_write_en = _guard10991;
assign cond439_clk = clk;
assign cond439_reset = reset;
assign cond439_in =
  _guard10992 ? idx_between_19_35_reg_out :
  1'd0;
assign cond464_write_en = _guard10993;
assign cond464_clk = clk;
assign cond464_reset = reset;
assign cond464_in =
  _guard10994 ? idx_between_41_42_reg_out :
  1'd0;
assign cond478_write_en = _guard10995;
assign cond478_clk = clk;
assign cond478_reset = reset;
assign cond478_in =
  _guard10996 ? idx_between_10_14_reg_out :
  1'd0;
assign cond494_write_en = _guard10997;
assign cond494_clk = clk;
assign cond494_reset = reset;
assign cond494_in =
  _guard10998 ? idx_between_14_18_reg_out :
  1'd0;
assign cond_wire498_in =
  _guard10999 ? idx_between_15_19_reg_out :
  _guard11002 ? cond498_out :
  1'd0;
assign cond508_write_en = _guard11003;
assign cond508_clk = clk;
assign cond508_reset = reset;
assign cond508_in =
  _guard11004 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire509_in =
  _guard11005 ? idx_between_37_38_reg_out :
  _guard11008 ? cond509_out :
  1'd0;
assign cond523_write_en = _guard11009;
assign cond523_clk = clk;
assign cond523_reset = reset;
assign cond523_in =
  _guard11010 ? idx_between_21_37_reg_out :
  1'd0;
assign cond527_write_en = _guard11011;
assign cond527_clk = clk;
assign cond527_reset = reset;
assign cond527_in =
  _guard11012 ? idx_between_22_38_reg_out :
  1'd0;
assign cond544_write_en = _guard11013;
assign cond544_clk = clk;
assign cond544_reset = reset;
assign cond544_in =
  _guard11014 ? idx_between_11_27_reg_out :
  1'd0;
assign cond_wire544_in =
  _guard11015 ? idx_between_11_27_reg_out :
  _guard11018 ? cond544_out :
  1'd0;
assign cond_wire554_in =
  _guard11021 ? cond554_out :
  _guard11022 ? idx_between_33_34_reg_out :
  1'd0;
assign cond563_write_en = _guard11023;
assign cond563_clk = clk;
assign cond563_reset = reset;
assign cond563_in =
  _guard11024 ? idx_between_16_20_reg_out :
  1'd0;
assign cond565_write_en = _guard11025;
assign cond565_clk = clk;
assign cond565_reset = reset;
assign cond565_in =
  _guard11026 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire569_in =
  _guard11029 ? cond569_out :
  _guard11030 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire580_in =
  _guard11031 ? idx_between_20_36_reg_out :
  _guard11034 ? cond580_out :
  1'd0;
assign cond583_write_en = _guard11035;
assign cond583_clk = clk;
assign cond583_reset = reset;
assign cond583_in =
  _guard11036 ? idx_between_21_25_reg_out :
  1'd0;
assign cond_wire598_in =
  _guard11037 ? idx_between_44_45_reg_out :
  _guard11040 ? cond598_out :
  1'd0;
assign cond_wire600_in =
  _guard11043 ? cond600_out :
  _guard11044 ? idx_between_10_14_reg_out :
  1'd0;
assign cond_wire612_in =
  _guard11045 ? idx_between_13_17_reg_out :
  _guard11048 ? cond612_out :
  1'd0;
assign cond_wire614_in =
  _guard11049 ? idx_between_17_33_reg_out :
  _guard11052 ? cond614_out :
  1'd0;
assign cond_wire623_in =
  _guard11053 ? idx_between_35_36_reg_out :
  _guard11056 ? cond623_out :
  1'd0;
assign cond629_write_en = _guard11057;
assign cond629_clk = clk;
assign cond629_reset = reset;
assign cond629_in =
  _guard11058 ? idx_between_17_33_reg_out :
  1'd0;
assign cond_wire642_in =
  _guard11061 ? cond642_out :
  _guard11062 ? idx_between_24_40_reg_out :
  1'd0;
assign cond652_write_en = _guard11063;
assign cond652_clk = clk;
assign cond652_reset = reset;
assign cond652_in =
  _guard11064 ? idx_between_23_27_reg_out :
  1'd0;
assign cond660_write_en = _guard11065;
assign cond660_clk = clk;
assign cond660_reset = reset;
assign cond660_in =
  _guard11066 ? idx_between_25_29_reg_out :
  1'd0;
assign cond687_write_en = _guard11067;
assign cond687_clk = clk;
assign cond687_reset = reset;
assign cond687_in =
  _guard11068 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire690_in =
  _guard11069 ? idx_between_17_33_reg_out :
  _guard11072 ? cond690_out :
  1'd0;
assign cond701_write_en = _guard11073;
assign cond701_clk = clk;
assign cond701_reset = reset;
assign cond701_in =
  _guard11074 ? idx_between_20_24_reg_out :
  1'd0;
assign cond736_write_en = _guard11075;
assign cond736_clk = clk;
assign cond736_reset = reset;
assign cond736_in =
  _guard11076 ? idx_between_17_33_reg_out :
  1'd0;
assign cond746_write_en = _guard11077;
assign cond746_clk = clk;
assign cond746_reset = reset;
assign cond746_in =
  _guard11078 ? idx_between_16_20_reg_out :
  1'd0;
assign cond_wire747_in =
  _guard11079 ? idx_between_16_32_reg_out :
  _guard11082 ? cond747_out :
  1'd0;
assign cond771_write_en = _guard11083;
assign cond771_clk = clk;
assign cond771_reset = reset;
assign cond771_in =
  _guard11084 ? idx_between_22_38_reg_out :
  1'd0;
assign cond776_write_en = _guard11085;
assign cond776_clk = clk;
assign cond776_reset = reset;
assign cond776_in =
  _guard11086 ? idx_between_27_43_reg_out :
  1'd0;
assign cond779_write_en = _guard11087;
assign cond779_clk = clk;
assign cond779_reset = reset;
assign cond779_in =
  _guard11088 ? idx_between_24_40_reg_out :
  1'd0;
assign cond_wire781_in =
  _guard11091 ? cond781_out :
  _guard11092 ? idx_between_44_45_reg_out :
  1'd0;
assign cond799_write_en = _guard11093;
assign cond799_clk = clk;
assign cond799_reset = reset;
assign cond799_in =
  _guard11094 ? idx_between_14_18_reg_out :
  1'd0;
assign cond_wire800_in =
  _guard11097 ? cond800_out :
  _guard11098 ? idx_between_14_30_reg_out :
  1'd0;
assign cond814_write_en = _guard11099;
assign cond814_clk = clk;
assign cond814_reset = reset;
assign cond814_in =
  _guard11100 ? idx_between_37_38_reg_out :
  1'd0;
assign cond_wire823_in =
  _guard11103 ? cond823_out :
  _guard11104 ? idx_between_20_24_reg_out :
  1'd0;
assign cond828_write_en = _guard11105;
assign cond828_clk = clk;
assign cond828_reset = reset;
assign cond828_in =
  _guard11106 ? idx_between_21_37_reg_out :
  1'd0;
assign cond840_write_en = _guard11107;
assign cond840_clk = clk;
assign cond840_reset = reset;
assign cond840_in =
  _guard11108 ? idx_between_24_40_reg_out :
  1'd0;
assign cond844_write_en = _guard11109;
assign cond844_clk = clk;
assign cond844_reset = reset;
assign cond844_in =
  _guard11110 ? idx_between_25_41_reg_out :
  1'd0;
assign cond858_write_en = _guard11111;
assign cond858_clk = clk;
assign cond858_reset = reset;
assign cond858_in =
  _guard11112 ? idx_between_48_49_reg_out :
  1'd0;
assign cond859_write_en = _guard11113;
assign cond859_clk = clk;
assign cond859_reset = reset;
assign cond859_in =
  _guard11114 ? idx_between_13_29_reg_out :
  1'd0;
assign cond862_write_en = _guard11115;
assign cond862_clk = clk;
assign cond862_reset = reset;
assign cond862_in =
  _guard11116 ? idx_between_18_34_reg_out :
  1'd0;
assign cond_wire868_in =
  _guard11117 ? idx_between_16_20_reg_out :
  _guard11120 ? cond868_out :
  1'd0;
assign cond_wire870_in =
  _guard11121 ? idx_between_20_36_reg_out :
  _guard11124 ? cond870_out :
  1'd0;
assign cond874_write_en = _guard11125;
assign cond874_clk = clk;
assign cond874_reset = reset;
assign cond874_in =
  _guard11126 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire875_in =
  _guard11129 ? cond875_out :
  _guard11130 ? idx_between_37_38_reg_out :
  1'd0;
assign cond_wire880_in =
  _guard11131 ? idx_between_19_23_reg_out :
  _guard11134 ? cond880_out :
  1'd0;
assign cond882_write_en = _guard11135;
assign cond882_clk = clk;
assign cond882_reset = reset;
assign cond882_in =
  _guard11136 ? idx_between_23_39_reg_out :
  1'd0;
assign cond890_write_en = _guard11137;
assign cond890_clk = clk;
assign cond890_reset = reset;
assign cond890_in =
  _guard11138 ? idx_between_25_41_reg_out :
  1'd0;
assign cond897_write_en = _guard11139;
assign cond897_clk = clk;
assign cond897_reset = reset;
assign cond897_in =
  _guard11140 ? idx_between_23_39_reg_out :
  1'd0;
assign cond903_write_en = _guard11141;
assign cond903_clk = clk;
assign cond903_reset = reset;
assign cond903_in =
  _guard11142 ? idx_between_44_45_reg_out :
  1'd0;
assign cond906_write_en = _guard11143;
assign cond906_clk = clk;
assign cond906_reset = reset;
assign cond906_in =
  _guard11144 ? idx_between_29_45_reg_out :
  1'd0;
assign cond918_write_en = _guard11145;
assign cond918_clk = clk;
assign cond918_reset = reset;
assign cond918_in =
  _guard11146 ? idx_between_32_48_reg_out :
  1'd0;
assign cond_wire937_in =
  _guard11147 ? idx_between_18_22_reg_out :
  _guard11150 ? cond937_out :
  1'd0;
assign cond_wire951_in =
  _guard11153 ? cond951_out :
  _guard11154 ? idx_between_25_41_reg_out :
  1'd0;
assign cond962_write_en = _guard11155;
assign cond962_clk = clk;
assign cond962_reset = reset;
assign cond962_in =
  _guard11156 ? idx_between_24_40_reg_out :
  1'd0;
assign cond974_write_en = _guard11157;
assign cond974_clk = clk;
assign cond974_reset = reset;
assign cond974_in =
  _guard11158 ? idx_between_27_43_reg_out :
  1'd0;
assign cond_wire987_in =
  _guard11161 ? cond987_out :
  _guard11162 ? idx_between_34_50_reg_out :
  1'd0;
assign cond992_write_en = _guard11163;
assign cond992_clk = clk;
assign cond992_reset = reset;
assign cond992_in =
  _guard11164 ? idx_between_20_36_reg_out :
  1'd0;
assign cond994_write_en = _guard11165;
assign cond994_clk = clk;
assign cond994_reset = reset;
assign cond994_in =
  _guard11166 ? idx_between_17_21_reg_out :
  1'd0;
assign cond1010_write_en = _guard11167;
assign cond1010_clk = clk;
assign cond1010_reset = reset;
assign cond1010_in =
  _guard11168 ? idx_between_21_25_reg_out :
  1'd0;
assign cond_wire1015_in =
  _guard11169 ? idx_between_22_38_reg_out :
  _guard11172 ? cond1015_out :
  1'd0;
assign cond1025_write_en = _guard11173;
assign cond1025_clk = clk;
assign cond1025_reset = reset;
assign cond1025_in =
  _guard11174 ? idx_between_44_45_reg_out :
  1'd0;
assign cond_wire1041_in =
  _guard11177 ? cond1041_out :
  _guard11178 ? idx_between_48_49_reg_out :
  1'd0;
assign cond_wire1042_in =
  _guard11179 ? idx_between_29_33_reg_out :
  _guard11182 ? cond1042_out :
  1'd0;
assign cond_wire1052_in =
  _guard11183 ? idx_between_51_52_reg_out :
  _guard11186 ? cond1052_out :
  1'd0;
assign pe_0_2_mul_ready =
  _guard11189 ? 1'd1 :
  _guard11192 ? 1'd0 :
  1'd0;
assign pe_0_2_clk = clk;
assign pe_0_2_top =
  _guard11205 ? top_0_2_out :
  32'd0;
assign pe_0_2_left =
  _guard11218 ? left_0_2_out :
  32'd0;
assign pe_0_2_reset = reset;
assign pe_0_2_go = _guard11231;
assign pe_0_12_mul_ready =
  _guard11234 ? 1'd1 :
  _guard11237 ? 1'd0 :
  1'd0;
assign pe_0_12_clk = clk;
assign pe_0_12_top =
  _guard11250 ? top_0_12_out :
  32'd0;
assign pe_0_12_left =
  _guard11263 ? left_0_12_out :
  32'd0;
assign pe_0_12_reset = reset;
assign pe_0_12_go = _guard11276;
assign pe_0_15_mul_ready =
  _guard11279 ? 1'd1 :
  _guard11282 ? 1'd0 :
  1'd0;
assign pe_0_15_clk = clk;
assign pe_0_15_top =
  _guard11295 ? top_0_15_out :
  32'd0;
assign pe_0_15_left =
  _guard11308 ? left_0_15_out :
  32'd0;
assign pe_0_15_reset = reset;
assign pe_0_15_go = _guard11321;
assign pe_1_6_mul_ready =
  _guard11324 ? 1'd1 :
  _guard11327 ? 1'd0 :
  1'd0;
assign pe_1_6_clk = clk;
assign pe_1_6_top =
  _guard11340 ? top_1_6_out :
  32'd0;
assign pe_1_6_left =
  _guard11353 ? left_1_6_out :
  32'd0;
assign pe_1_6_reset = reset;
assign pe_1_6_go = _guard11366;
assign left_3_5_write_en = _guard11369;
assign left_3_5_clk = clk;
assign left_3_5_reset = reset;
assign left_3_5_in = left_3_4_out;
assign pe_3_13_mul_ready =
  _guard11375 ? 1'd1 :
  _guard11378 ? 1'd0 :
  1'd0;
assign pe_3_13_clk = clk;
assign pe_3_13_top =
  _guard11391 ? top_3_13_out :
  32'd0;
assign pe_3_13_left =
  _guard11404 ? left_3_13_out :
  32'd0;
assign pe_3_13_reset = reset;
assign pe_3_13_go = _guard11417;
assign pe_3_14_mul_ready =
  _guard11420 ? 1'd1 :
  _guard11423 ? 1'd0 :
  1'd0;
assign pe_3_14_clk = clk;
assign pe_3_14_top =
  _guard11436 ? top_3_14_out :
  32'd0;
assign pe_3_14_left =
  _guard11449 ? left_3_14_out :
  32'd0;
assign pe_3_14_reset = reset;
assign pe_3_14_go = _guard11462;
assign left_4_8_write_en = _guard11465;
assign left_4_8_clk = clk;
assign left_4_8_reset = reset;
assign left_4_8_in = left_4_7_out;
assign pe_4_12_mul_ready =
  _guard11471 ? 1'd1 :
  _guard11474 ? 1'd0 :
  1'd0;
assign pe_4_12_clk = clk;
assign pe_4_12_top =
  _guard11487 ? top_4_12_out :
  32'd0;
assign pe_4_12_left =
  _guard11500 ? left_4_12_out :
  32'd0;
assign pe_4_12_reset = reset;
assign pe_4_12_go = _guard11513;
assign top_5_5_write_en = _guard11516;
assign top_5_5_clk = clk;
assign top_5_5_reset = reset;
assign top_5_5_in = top_4_5_out;
assign pe_5_9_mul_ready =
  _guard11522 ? 1'd1 :
  _guard11525 ? 1'd0 :
  1'd0;
assign pe_5_9_clk = clk;
assign pe_5_9_top =
  _guard11538 ? top_5_9_out :
  32'd0;
assign pe_5_9_left =
  _guard11551 ? left_5_9_out :
  32'd0;
assign pe_5_9_reset = reset;
assign pe_5_9_go = _guard11564;
assign pe_5_10_mul_ready =
  _guard11567 ? 1'd1 :
  _guard11570 ? 1'd0 :
  1'd0;
assign pe_5_10_clk = clk;
assign pe_5_10_top =
  _guard11583 ? top_5_10_out :
  32'd0;
assign pe_5_10_left =
  _guard11596 ? left_5_10_out :
  32'd0;
assign pe_5_10_reset = reset;
assign pe_5_10_go = _guard11609;
assign left_5_11_write_en = _guard11612;
assign left_5_11_clk = clk;
assign left_5_11_reset = reset;
assign left_5_11_in = left_5_10_out;
assign left_6_1_write_en = _guard11618;
assign left_6_1_clk = clk;
assign left_6_1_reset = reset;
assign left_6_1_in = left_6_0_out;
assign pe_6_5_mul_ready =
  _guard11624 ? 1'd1 :
  _guard11627 ? 1'd0 :
  1'd0;
assign pe_6_5_clk = clk;
assign pe_6_5_top =
  _guard11640 ? top_6_5_out :
  32'd0;
assign pe_6_5_left =
  _guard11653 ? left_6_5_out :
  32'd0;
assign pe_6_5_reset = reset;
assign pe_6_5_go = _guard11666;
assign left_6_7_write_en = _guard11669;
assign left_6_7_clk = clk;
assign left_6_7_reset = reset;
assign left_6_7_in = left_6_6_out;
assign pe_6_12_mul_ready =
  _guard11675 ? 1'd1 :
  _guard11678 ? 1'd0 :
  1'd0;
assign pe_6_12_clk = clk;
assign pe_6_12_top =
  _guard11691 ? top_6_12_out :
  32'd0;
assign pe_6_12_left =
  _guard11704 ? left_6_12_out :
  32'd0;
assign pe_6_12_reset = reset;
assign pe_6_12_go = _guard11717;
assign top_6_12_write_en = _guard11720;
assign top_6_12_clk = clk;
assign top_6_12_reset = reset;
assign top_6_12_in = top_5_12_out;
assign pe_7_0_mul_ready =
  _guard11726 ? 1'd1 :
  _guard11729 ? 1'd0 :
  1'd0;
assign pe_7_0_clk = clk;
assign pe_7_0_top =
  _guard11742 ? top_7_0_out :
  32'd0;
assign pe_7_0_left =
  _guard11755 ? left_7_0_out :
  32'd0;
assign pe_7_0_reset = reset;
assign pe_7_0_go = _guard11768;
assign top_7_4_write_en = _guard11771;
assign top_7_4_clk = clk;
assign top_7_4_reset = reset;
assign top_7_4_in = top_6_4_out;
assign pe_7_10_mul_ready =
  _guard11777 ? 1'd1 :
  _guard11780 ? 1'd0 :
  1'd0;
assign pe_7_10_clk = clk;
assign pe_7_10_top =
  _guard11793 ? top_7_10_out :
  32'd0;
assign pe_7_10_left =
  _guard11806 ? left_7_10_out :
  32'd0;
assign pe_7_10_reset = reset;
assign pe_7_10_go = _guard11819;
assign pe_8_0_mul_ready =
  _guard11822 ? 1'd1 :
  _guard11825 ? 1'd0 :
  1'd0;
assign pe_8_0_clk = clk;
assign pe_8_0_top =
  _guard11838 ? top_8_0_out :
  32'd0;
assign pe_8_0_left =
  _guard11851 ? left_8_0_out :
  32'd0;
assign pe_8_0_reset = reset;
assign pe_8_0_go = _guard11864;
assign left_8_4_write_en = _guard11867;
assign left_8_4_clk = clk;
assign left_8_4_reset = reset;
assign left_8_4_in = left_8_3_out;
assign pe_8_5_mul_ready =
  _guard11873 ? 1'd1 :
  _guard11876 ? 1'd0 :
  1'd0;
assign pe_8_5_clk = clk;
assign pe_8_5_top =
  _guard11889 ? top_8_5_out :
  32'd0;
assign pe_8_5_left =
  _guard11902 ? left_8_5_out :
  32'd0;
assign pe_8_5_reset = reset;
assign pe_8_5_go = _guard11915;
assign top_8_8_write_en = _guard11918;
assign top_8_8_clk = clk;
assign top_8_8_reset = reset;
assign top_8_8_in = top_7_8_out;
assign left_8_8_write_en = _guard11924;
assign left_8_8_clk = clk;
assign left_8_8_reset = reset;
assign left_8_8_in = left_8_7_out;
assign top_8_14_write_en = _guard11930;
assign top_8_14_clk = clk;
assign top_8_14_reset = reset;
assign top_8_14_in = top_7_14_out;
assign top_9_1_write_en = _guard11936;
assign top_9_1_clk = clk;
assign top_9_1_reset = reset;
assign top_9_1_in = top_8_1_out;
assign pe_9_6_mul_ready =
  _guard11942 ? 1'd1 :
  _guard11945 ? 1'd0 :
  1'd0;
assign pe_9_6_clk = clk;
assign pe_9_6_top =
  _guard11958 ? top_9_6_out :
  32'd0;
assign pe_9_6_left =
  _guard11971 ? left_9_6_out :
  32'd0;
assign pe_9_6_reset = reset;
assign pe_9_6_go = _guard11984;
assign left_9_9_write_en = _guard11987;
assign left_9_9_clk = clk;
assign left_9_9_reset = reset;
assign left_9_9_in = left_9_8_out;
assign left_9_10_write_en = _guard11993;
assign left_9_10_clk = clk;
assign left_9_10_reset = reset;
assign left_9_10_in = left_9_9_out;
assign top_9_15_write_en = _guard11999;
assign top_9_15_clk = clk;
assign top_9_15_reset = reset;
assign top_9_15_in = top_8_15_out;
assign top_10_0_write_en = _guard12005;
assign top_10_0_clk = clk;
assign top_10_0_reset = reset;
assign top_10_0_in = top_9_0_out;
assign top_10_5_write_en = _guard12011;
assign top_10_5_clk = clk;
assign top_10_5_reset = reset;
assign top_10_5_in = top_9_5_out;
assign left_10_10_write_en = _guard12017;
assign left_10_10_clk = clk;
assign left_10_10_reset = reset;
assign left_10_10_in = left_10_9_out;
assign pe_10_12_mul_ready =
  _guard12023 ? 1'd1 :
  _guard12026 ? 1'd0 :
  1'd0;
assign pe_10_12_clk = clk;
assign pe_10_12_top =
  _guard12039 ? top_10_12_out :
  32'd0;
assign pe_10_12_left =
  _guard12052 ? left_10_12_out :
  32'd0;
assign pe_10_12_reset = reset;
assign pe_10_12_go = _guard12065;
assign top_11_1_write_en = _guard12068;
assign top_11_1_clk = clk;
assign top_11_1_reset = reset;
assign top_11_1_in = top_10_1_out;
assign pe_11_6_mul_ready =
  _guard12074 ? 1'd1 :
  _guard12077 ? 1'd0 :
  1'd0;
assign pe_11_6_clk = clk;
assign pe_11_6_top =
  _guard12090 ? top_11_6_out :
  32'd0;
assign pe_11_6_left =
  _guard12103 ? left_11_6_out :
  32'd0;
assign pe_11_6_reset = reset;
assign pe_11_6_go = _guard12116;
assign pe_11_7_mul_ready =
  _guard12119 ? 1'd1 :
  _guard12122 ? 1'd0 :
  1'd0;
assign pe_11_7_clk = clk;
assign pe_11_7_top =
  _guard12135 ? top_11_7_out :
  32'd0;
assign pe_11_7_left =
  _guard12148 ? left_11_7_out :
  32'd0;
assign pe_11_7_reset = reset;
assign pe_11_7_go = _guard12161;
assign top_12_1_write_en = _guard12164;
assign top_12_1_clk = clk;
assign top_12_1_reset = reset;
assign top_12_1_in = top_11_1_out;
assign pe_12_3_mul_ready =
  _guard12170 ? 1'd1 :
  _guard12173 ? 1'd0 :
  1'd0;
assign pe_12_3_clk = clk;
assign pe_12_3_top =
  _guard12186 ? top_12_3_out :
  32'd0;
assign pe_12_3_left =
  _guard12199 ? left_12_3_out :
  32'd0;
assign pe_12_3_reset = reset;
assign pe_12_3_go = _guard12212;
assign pe_12_4_mul_ready =
  _guard12215 ? 1'd1 :
  _guard12218 ? 1'd0 :
  1'd0;
assign pe_12_4_clk = clk;
assign pe_12_4_top =
  _guard12231 ? top_12_4_out :
  32'd0;
assign pe_12_4_left =
  _guard12244 ? left_12_4_out :
  32'd0;
assign pe_12_4_reset = reset;
assign pe_12_4_go = _guard12257;
assign left_12_9_write_en = _guard12260;
assign left_12_9_clk = clk;
assign left_12_9_reset = reset;
assign left_12_9_in = left_12_8_out;
assign top_12_11_write_en = _guard12266;
assign top_12_11_clk = clk;
assign top_12_11_reset = reset;
assign top_12_11_in = top_11_11_out;
assign top_12_12_write_en = _guard12272;
assign top_12_12_clk = clk;
assign top_12_12_reset = reset;
assign top_12_12_in = top_11_12_out;
assign pe_13_0_mul_ready =
  _guard12278 ? 1'd1 :
  _guard12281 ? 1'd0 :
  1'd0;
assign pe_13_0_clk = clk;
assign pe_13_0_top =
  _guard12294 ? top_13_0_out :
  32'd0;
assign pe_13_0_left =
  _guard12307 ? left_13_0_out :
  32'd0;
assign pe_13_0_reset = reset;
assign pe_13_0_go = _guard12320;
assign pe_13_3_mul_ready =
  _guard12323 ? 1'd1 :
  _guard12326 ? 1'd0 :
  1'd0;
assign pe_13_3_clk = clk;
assign pe_13_3_top =
  _guard12339 ? top_13_3_out :
  32'd0;
assign pe_13_3_left =
  _guard12352 ? left_13_3_out :
  32'd0;
assign pe_13_3_reset = reset;
assign pe_13_3_go = _guard12365;
assign left_13_7_write_en = _guard12368;
assign left_13_7_clk = clk;
assign left_13_7_reset = reset;
assign left_13_7_in = left_13_6_out;
assign left_13_8_write_en = _guard12374;
assign left_13_8_clk = clk;
assign left_13_8_reset = reset;
assign left_13_8_in = left_13_7_out;
assign pe_13_13_mul_ready =
  _guard12380 ? 1'd1 :
  _guard12383 ? 1'd0 :
  1'd0;
assign pe_13_13_clk = clk;
assign pe_13_13_top =
  _guard12396 ? top_13_13_out :
  32'd0;
assign pe_13_13_left =
  _guard12409 ? left_13_13_out :
  32'd0;
assign pe_13_13_reset = reset;
assign pe_13_13_go = _guard12422;
assign left_13_13_write_en = _guard12425;
assign left_13_13_clk = clk;
assign left_13_13_reset = reset;
assign left_13_13_in = left_13_12_out;
assign left_14_3_write_en = _guard12431;
assign left_14_3_clk = clk;
assign left_14_3_reset = reset;
assign left_14_3_in = left_14_2_out;
assign top_15_5_write_en = _guard12437;
assign top_15_5_clk = clk;
assign top_15_5_reset = reset;
assign top_15_5_in = top_14_5_out;
assign left_15_7_write_en = _guard12443;
assign left_15_7_clk = clk;
assign left_15_7_reset = reset;
assign left_15_7_in = left_15_6_out;
assign pe_15_13_mul_ready =
  _guard12449 ? 1'd1 :
  _guard12452 ? 1'd0 :
  1'd0;
assign pe_15_13_clk = clk;
assign pe_15_13_top =
  _guard12465 ? top_15_13_out :
  32'd0;
assign pe_15_13_left =
  _guard12478 ? left_15_13_out :
  32'd0;
assign pe_15_13_reset = reset;
assign pe_15_13_go = _guard12491;
assign t0_idx_write_en = _guard12498;
assign t0_idx_clk = clk;
assign t0_idx_reset = reset;
assign t0_idx_in =
  _guard12501 ? 5'd0 :
  _guard12504 ? t0_add_out :
  'x;
assign t4_idx_write_en = _guard12511;
assign t4_idx_clk = clk;
assign t4_idx_reset = reset;
assign t4_idx_in =
  _guard12514 ? 5'd0 :
  _guard12517 ? t4_add_out :
  'x;
assign t6_idx_write_en = _guard12524;
assign t6_idx_clk = clk;
assign t6_idx_reset = reset;
assign t6_idx_in =
  _guard12527 ? 5'd0 :
  _guard12530 ? t6_add_out :
  'x;
assign t12_idx_write_en = _guard12537;
assign t12_idx_clk = clk;
assign t12_idx_reset = reset;
assign t12_idx_in =
  _guard12540 ? 5'd0 :
  _guard12543 ? t12_add_out :
  'x;
assign t14_idx_write_en = _guard12550;
assign t14_idx_clk = clk;
assign t14_idx_reset = reset;
assign t14_idx_in =
  _guard12553 ? 5'd0 :
  _guard12556 ? t14_add_out :
  'x;
assign l1_idx_write_en = _guard12563;
assign l1_idx_clk = clk;
assign l1_idx_reset = reset;
assign l1_idx_in =
  _guard12566 ? l1_add_out :
  _guard12569 ? 5'd0 :
  'x;
assign l5_add_left = 5'd1;
assign l5_add_right = l5_idx_out;
assign idx_add_left = idx_out;
assign idx_add_right = 6'd1;
assign idx_between_26_30_comb_left = index_ge_26_out;
assign idx_between_26_30_comb_right = index_lt_30_out;
assign index_lt_37_left = idx_add_out;
assign index_lt_37_right = 6'd37;
assign idx_between_31_47_reg_write_en = _guard12586;
assign idx_between_31_47_reg_clk = clk;
assign idx_between_31_47_reg_reset = reset;
assign idx_between_31_47_reg_in =
  _guard12587 ? idx_between_31_47_comb_out :
  _guard12590 ? 1'd0 :
  'x;
assign idx_between_23_27_comb_left = index_ge_23_out;
assign idx_between_23_27_comb_right = index_lt_27_out;
assign index_lt_16_left = idx_add_out;
assign index_lt_16_right = 6'd16;
assign idx_between_1_17_comb_left = index_ge_1_out;
assign idx_between_1_17_comb_right = index_lt_17_out;
assign index_ge_47_left = idx_add_out;
assign index_ge_47_right = 6'd47;
assign index_lt_49_left = idx_add_out;
assign index_lt_49_right = 6'd49;
assign index_ge_38_left = idx_add_out;
assign index_ge_38_right = 6'd38;
assign idx_between_48_49_reg_write_en = _guard12607;
assign idx_between_48_49_reg_clk = clk;
assign idx_between_48_49_reg_reset = reset;
assign idx_between_48_49_reg_in =
  _guard12608 ? idx_between_48_49_comb_out :
  _guard12611 ? 1'd0 :
  'x;
assign index_ge_7_left = idx_add_out;
assign index_ge_7_right = 6'd7;
assign idx_between_50_51_comb_left = index_ge_50_out;
assign idx_between_50_51_comb_right = index_lt_51_out;
assign index_lt_52_left = idx_add_out;
assign index_lt_52_right = 6'd52;
assign idx_between_32_48_reg_write_en = _guard12622;
assign idx_between_32_48_reg_clk = clk;
assign idx_between_32_48_reg_reset = reset;
assign idx_between_32_48_reg_in =
  _guard12623 ? idx_between_32_48_comb_out :
  _guard12626 ? 1'd0 :
  'x;
assign idx_between_21_22_comb_left = index_ge_21_out;
assign idx_between_21_22_comb_right = index_lt_22_out;
assign idx_between_18_34_reg_write_en = _guard12633;
assign idx_between_18_34_reg_clk = clk;
assign idx_between_18_34_reg_reset = reset;
assign idx_between_18_34_reg_in =
  _guard12634 ? idx_between_18_34_comb_out :
  _guard12637 ? 1'd0 :
  'x;
assign idx_between_12_16_comb_left = index_ge_12_out;
assign idx_between_12_16_comb_right = index_lt_16_out;
assign idx_between_8_12_reg_write_en = _guard12644;
assign idx_between_8_12_reg_clk = clk;
assign idx_between_8_12_reg_reset = reset;
assign idx_between_8_12_reg_in =
  _guard12647 ? 1'd0 :
  _guard12648 ? idx_between_8_12_comb_out :
  'x;
assign idx_between_39_40_comb_left = index_ge_39_out;
assign idx_between_39_40_comb_right = index_lt_40_out;
assign cond3_write_en = _guard12651;
assign cond3_clk = clk;
assign cond3_reset = reset;
assign cond3_in =
  _guard12652 ? idx_between_21_22_reg_out :
  1'd0;
assign cond13_write_en = _guard12653;
assign cond13_clk = clk;
assign cond13_reset = reset;
assign cond13_in =
  _guard12654 ? idx_between_23_24_reg_out :
  1'd0;
assign cond29_write_en = _guard12655;
assign cond29_clk = clk;
assign cond29_reset = reset;
assign cond29_in =
  _guard12656 ? idx_between_6_22_reg_out :
  1'd0;
assign cond41_write_en = _guard12657;
assign cond41_clk = clk;
assign cond41_reset = reset;
assign cond41_in =
  _guard12658 ? idx_between_9_25_reg_out :
  1'd0;
assign cond54_write_en = _guard12659;
assign cond54_clk = clk;
assign cond54_reset = reset;
assign cond54_in =
  _guard12660 ? idx_between_11_27_reg_out :
  1'd0;
assign cond64_write_en = _guard12661;
assign cond64_clk = clk;
assign cond64_reset = reset;
assign cond64_in =
  _guard12662 ? idx_between_13_29_reg_out :
  1'd0;
assign cond67_write_en = _guard12663;
assign cond67_clk = clk;
assign cond67_reset = reset;
assign cond67_in =
  _guard12664 ? idx_between_18_34_reg_out :
  1'd0;
assign cond68_write_en = _guard12665;
assign cond68_clk = clk;
assign cond68_reset = reset;
assign cond68_in =
  _guard12666 ? idx_between_34_35_reg_out :
  1'd0;
assign cond77_write_en = _guard12667;
assign cond77_clk = clk;
assign cond77_reset = reset;
assign cond77_in =
  _guard12668 ? idx_between_20_36_reg_out :
  1'd0;
assign cond89_write_en = _guard12669;
assign cond89_clk = clk;
assign cond89_reset = reset;
assign cond89_in =
  _guard12670 ? idx_between_4_20_reg_out :
  1'd0;
assign cond94_write_en = _guard12671;
assign cond94_clk = clk;
assign cond94_reset = reset;
assign cond94_in =
  _guard12672 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire125_in =
  _guard12673 ? idx_between_13_29_reg_out :
  _guard12676 ? cond125_out :
  1'd0;
assign cond128_write_en = _guard12677;
assign cond128_clk = clk;
assign cond128_reset = reset;
assign cond128_in =
  _guard12678 ? idx_between_14_18_reg_out :
  1'd0;
assign cond131_write_en = _guard12679;
assign cond131_clk = clk;
assign cond131_reset = reset;
assign cond131_in =
  _guard12680 ? idx_between_34_35_reg_out :
  1'd0;
assign cond132_write_en = _guard12681;
assign cond132_clk = clk;
assign cond132_reset = reset;
assign cond132_in =
  _guard12682 ? idx_between_15_19_reg_out :
  1'd0;
assign cond_wire132_in =
  _guard12683 ? idx_between_15_19_reg_out :
  _guard12686 ? cond132_out :
  1'd0;
assign cond134_write_en = _guard12687;
assign cond134_clk = clk;
assign cond134_reset = reset;
assign cond134_in =
  _guard12688 ? idx_between_19_35_reg_out :
  1'd0;
assign cond136_write_en = _guard12689;
assign cond136_clk = clk;
assign cond136_reset = reset;
assign cond136_in =
  _guard12690 ? idx_between_16_20_reg_out :
  1'd0;
assign cond139_write_en = _guard12691;
assign cond139_clk = clk;
assign cond139_reset = reset;
assign cond139_in =
  _guard12692 ? idx_between_36_37_reg_out :
  1'd0;
assign cond140_write_en = _guard12693;
assign cond140_clk = clk;
assign cond140_reset = reset;
assign cond140_in =
  _guard12694 ? idx_between_17_21_reg_out :
  1'd0;
assign cond_wire142_in =
  _guard12695 ? idx_between_21_37_reg_out :
  _guard12698 ? cond142_out :
  1'd0;
assign cond_wire148_in =
  _guard12699 ? idx_between_23_24_reg_out :
  _guard12702 ? cond148_out :
  1'd0;
assign cond_wire151_in =
  _guard12705 ? cond151_out :
  _guard12706 ? idx_between_8_24_reg_out :
  1'd0;
assign cond_wire161_in =
  _guard12707 ? idx_between_7_11_reg_out :
  _guard12710 ? cond161_out :
  1'd0;
assign cond_wire162_in =
  _guard12711 ? idx_between_7_23_reg_out :
  _guard12714 ? cond162_out :
  1'd0;
assign cond_wire165_in =
  _guard12715 ? idx_between_8_12_reg_out :
  _guard12718 ? cond165_out :
  1'd0;
assign cond_wire171_in =
  _guard12719 ? idx_between_13_29_reg_out :
  _guard12722 ? cond171_out :
  1'd0;
assign cond172_write_en = _guard12723;
assign cond172_clk = clk;
assign cond172_reset = reset;
assign cond172_in =
  _guard12724 ? idx_between_29_30_reg_out :
  1'd0;
assign cond_wire177_in =
  _guard12727 ? cond177_out :
  _guard12728 ? idx_between_11_15_reg_out :
  1'd0;
assign cond183_write_en = _guard12729;
assign cond183_clk = clk;
assign cond183_reset = reset;
assign cond183_in =
  _guard12730 ? idx_between_16_32_reg_out :
  1'd0;
assign cond187_write_en = _guard12731;
assign cond187_clk = clk;
assign cond187_reset = reset;
assign cond187_in =
  _guard12732 ? idx_between_17_33_reg_out :
  1'd0;
assign cond190_write_en = _guard12733;
assign cond190_clk = clk;
assign cond190_reset = reset;
assign cond190_in =
  _guard12734 ? idx_between_14_30_reg_out :
  1'd0;
assign cond191_write_en = _guard12735;
assign cond191_clk = clk;
assign cond191_reset = reset;
assign cond191_in =
  _guard12736 ? idx_between_18_34_reg_out :
  1'd0;
assign cond223_write_en = _guard12737;
assign cond223_clk = clk;
assign cond223_reset = reset;
assign cond223_in =
  _guard12738 ? idx_between_7_23_reg_out :
  1'd0;
assign cond238_write_en = _guard12739;
assign cond238_clk = clk;
assign cond238_reset = reset;
assign cond238_in =
  _guard12740 ? idx_between_11_15_reg_out :
  1'd0;
assign cond244_write_en = _guard12741;
assign cond244_clk = clk;
assign cond244_reset = reset;
assign cond244_in =
  _guard12742 ? idx_between_16_32_reg_out :
  1'd0;
assign cond_wire252_in =
  _guard12743 ? idx_between_18_34_reg_out :
  _guard12746 ? cond252_out :
  1'd0;
assign cond_wire262_in =
  _guard12747 ? idx_between_17_21_reg_out :
  _guard12750 ? cond262_out :
  1'd0;
assign cond_wire264_in =
  _guard12753 ? cond264_out :
  _guard12754 ? idx_between_21_37_reg_out :
  1'd0;
assign cond265_write_en = _guard12755;
assign cond265_clk = clk;
assign cond265_reset = reset;
assign cond265_in =
  _guard12756 ? idx_between_37_38_reg_out :
  1'd0;
assign cond_wire267_in =
  _guard12757 ? idx_between_18_34_reg_out :
  _guard12760 ? cond267_out :
  1'd0;
assign cond280_write_en = _guard12761;
assign cond280_clk = clk;
assign cond280_reset = reset;
assign cond280_in =
  _guard12762 ? idx_between_6_22_reg_out :
  1'd0;
assign cond_wire289_in =
  _guard12765 ? cond289_out :
  _guard12766 ? idx_between_12_28_reg_out :
  1'd0;
assign cond316_write_en = _guard12767;
assign cond316_clk = clk;
assign cond316_reset = reset;
assign cond316_in =
  _guard12768 ? idx_between_15_31_reg_out :
  1'd0;
assign cond317_write_en = _guard12769;
assign cond317_clk = clk;
assign cond317_reset = reset;
assign cond317_in =
  _guard12770 ? idx_between_19_35_reg_out :
  1'd0;
assign cond321_write_en = _guard12771;
assign cond321_clk = clk;
assign cond321_reset = reset;
assign cond321_in =
  _guard12772 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire363_in =
  _guard12773 ? idx_between_31_32_reg_out :
  _guard12776 ? cond363_out :
  1'd0;
assign cond367_write_en = _guard12777;
assign cond367_clk = clk;
assign cond367_reset = reset;
assign cond367_in =
  _guard12778 ? idx_between_32_33_reg_out :
  1'd0;
assign cond370_write_en = _guard12779;
assign cond370_clk = clk;
assign cond370_reset = reset;
assign cond370_in =
  _guard12780 ? idx_between_17_33_reg_out :
  1'd0;
assign cond371_write_en = _guard12781;
assign cond371_clk = clk;
assign cond371_reset = reset;
assign cond371_in =
  _guard12782 ? idx_between_33_34_reg_out :
  1'd0;
assign cond377_write_en = _guard12783;
assign cond377_clk = clk;
assign cond377_reset = reset;
assign cond377_in =
  _guard12784 ? idx_between_15_31_reg_out :
  1'd0;
assign cond387_write_en = _guard12785;
assign cond387_clk = clk;
assign cond387_reset = reset;
assign cond387_in =
  _guard12786 ? idx_between_37_38_reg_out :
  1'd0;
assign cond391_write_en = _guard12787;
assign cond391_clk = clk;
assign cond391_reset = reset;
assign cond391_in =
  _guard12788 ? idx_between_38_39_reg_out :
  1'd0;
assign cond400_write_en = _guard12789;
assign cond400_clk = clk;
assign cond400_reset = reset;
assign cond400_in =
  _guard12790 ? idx_between_21_25_reg_out :
  1'd0;
assign cond_wire420_in =
  _guard12793 ? cond420_out :
  _guard12794 ? idx_between_30_31_reg_out :
  1'd0;
assign cond429_write_en = _guard12795;
assign cond429_clk = clk;
assign cond429_reset = reset;
assign cond429_in =
  _guard12796 ? idx_between_13_17_reg_out :
  1'd0;
assign cond444_write_en = _guard12797;
assign cond444_clk = clk;
assign cond444_reset = reset;
assign cond444_in =
  _guard12798 ? idx_between_36_37_reg_out :
  1'd0;
assign cond448_write_en = _guard12799;
assign cond448_clk = clk;
assign cond448_reset = reset;
assign cond448_in =
  _guard12800 ? idx_between_37_38_reg_out :
  1'd0;
assign cond453_write_en = _guard12801;
assign cond453_clk = clk;
assign cond453_reset = reset;
assign cond453_in =
  _guard12802 ? idx_between_19_23_reg_out :
  1'd0;
assign cond_wire465_in =
  _guard12805 ? cond465_out :
  _guard12806 ? idx_between_22_26_reg_out :
  1'd0;
assign cond_wire468_in =
  _guard12807 ? idx_between_42_43_reg_out :
  _guard12810 ? cond468_out :
  1'd0;
assign cond_wire476_in =
  _guard12813 ? cond476_out :
  _guard12814 ? idx_between_13_29_reg_out :
  1'd0;
assign cond_wire494_in =
  _guard12817 ? cond494_out :
  _guard12818 ? idx_between_14_18_reg_out :
  1'd0;
assign cond_wire508_in =
  _guard12821 ? cond508_out :
  _guard12822 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire519_in =
  _guard12823 ? idx_between_20_36_reg_out :
  _guard12826 ? cond519_out :
  1'd0;
assign cond_wire530_in =
  _guard12827 ? idx_between_23_27_reg_out :
  _guard12830 ? cond530_out :
  1'd0;
assign cond537_write_en = _guard12831;
assign cond537_clk = clk;
assign cond537_reset = reset;
assign cond537_in =
  _guard12832 ? idx_between_13_29_reg_out :
  1'd0;
assign cond_wire537_in =
  _guard12833 ? idx_between_13_29_reg_out :
  _guard12836 ? cond537_out :
  1'd0;
assign cond538_write_en = _guard12837;
assign cond538_clk = clk;
assign cond538_reset = reset;
assign cond538_in =
  _guard12838 ? idx_between_29_30_reg_out :
  1'd0;
assign cond_wire549_in =
  _guard12839 ? idx_between_16_32_reg_out :
  _guard12842 ? cond549_out :
  1'd0;
assign cond552_write_en = _guard12843;
assign cond552_clk = clk;
assign cond552_reset = reset;
assign cond552_in =
  _guard12844 ? idx_between_13_29_reg_out :
  1'd0;
assign cond_wire558_in =
  _guard12845 ? idx_between_34_35_reg_out :
  _guard12848 ? cond558_out :
  1'd0;
assign cond_wire559_in =
  _guard12849 ? idx_between_15_19_reg_out :
  _guard12852 ? cond559_out :
  1'd0;
assign cond560_write_en = _guard12853;
assign cond560_clk = clk;
assign cond560_reset = reset;
assign cond560_in =
  _guard12854 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire562_in =
  _guard12855 ? idx_between_35_36_reg_out :
  _guard12858 ? cond562_out :
  1'd0;
assign cond_wire567_in =
  _guard12859 ? idx_between_17_21_reg_out :
  _guard12862 ? cond567_out :
  1'd0;
assign cond585_write_en = _guard12863;
assign cond585_clk = clk;
assign cond585_reset = reset;
assign cond585_in =
  _guard12864 ? idx_between_25_41_reg_out :
  1'd0;
assign cond599_write_en = _guard12865;
assign cond599_clk = clk;
assign cond599_reset = reset;
assign cond599_in =
  _guard12866 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire606_in =
  _guard12869 ? cond606_out :
  _guard12870 ? idx_between_15_31_reg_out :
  1'd0;
assign cond617_write_en = _guard12871;
assign cond617_clk = clk;
assign cond617_reset = reset;
assign cond617_in =
  _guard12872 ? idx_between_14_30_reg_out :
  1'd0;
assign cond619_write_en = _guard12873;
assign cond619_clk = clk;
assign cond619_reset = reset;
assign cond619_in =
  _guard12874 ? idx_between_34_35_reg_out :
  1'd0;
assign cond625_write_en = _guard12875;
assign cond625_clk = clk;
assign cond625_reset = reset;
assign cond625_in =
  _guard12876 ? idx_between_16_32_reg_out :
  1'd0;
assign cond_wire625_in =
  _guard12877 ? idx_between_16_32_reg_out :
  _guard12880 ? cond625_out :
  1'd0;
assign cond653_write_en = _guard12881;
assign cond653_clk = clk;
assign cond653_reset = reset;
assign cond653_in =
  _guard12882 ? idx_between_23_39_reg_out :
  1'd0;
assign cond_wire659_in =
  _guard12885 ? cond659_out :
  _guard12886 ? idx_between_44_45_reg_out :
  1'd0;
assign cond685_write_en = _guard12887;
assign cond685_clk = clk;
assign cond685_reset = reset;
assign cond685_in =
  _guard12888 ? idx_between_16_20_reg_out :
  1'd0;
assign cond686_write_en = _guard12889;
assign cond686_clk = clk;
assign cond686_reset = reset;
assign cond686_in =
  _guard12890 ? idx_between_16_32_reg_out :
  1'd0;
assign cond692_write_en = _guard12891;
assign cond692_clk = clk;
assign cond692_reset = reset;
assign cond692_in =
  _guard12892 ? idx_between_37_38_reg_out :
  1'd0;
assign cond696_write_en = _guard12893;
assign cond696_clk = clk;
assign cond696_reset = reset;
assign cond696_in =
  _guard12894 ? idx_between_38_39_reg_out :
  1'd0;
assign cond_wire699_in =
  _guard12895 ? idx_between_23_39_reg_out :
  _guard12898 ? cond699_out :
  1'd0;
assign cond707_write_en = _guard12899;
assign cond707_clk = clk;
assign cond707_reset = reset;
assign cond707_in =
  _guard12900 ? idx_between_25_41_reg_out :
  1'd0;
assign cond714_write_en = _guard12901;
assign cond714_clk = clk;
assign cond714_reset = reset;
assign cond714_in =
  _guard12902 ? idx_between_23_39_reg_out :
  1'd0;
assign cond_wire719_in =
  _guard12903 ? idx_between_28_44_reg_out :
  _guard12906 ? cond719_out :
  1'd0;
assign cond748_write_en = _guard12907;
assign cond748_clk = clk;
assign cond748_reset = reset;
assign cond748_in =
  _guard12908 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire748_in =
  _guard12909 ? idx_between_20_36_reg_out :
  _guard12912 ? cond748_out :
  1'd0;
assign cond759_write_en = _guard12913;
assign cond759_clk = clk;
assign cond759_reset = reset;
assign cond759_in =
  _guard12914 ? idx_between_19_35_reg_out :
  1'd0;
assign cond762_write_en = _guard12915;
assign cond762_clk = clk;
assign cond762_reset = reset;
assign cond762_in =
  _guard12916 ? idx_between_20_24_reg_out :
  1'd0;
assign cond_wire763_in =
  _guard12919 ? cond763_out :
  _guard12920 ? idx_between_20_36_reg_out :
  1'd0;
assign cond773_write_en = _guard12921;
assign cond773_clk = clk;
assign cond773_reset = reset;
assign cond773_in =
  _guard12922 ? idx_between_42_43_reg_out :
  1'd0;
assign cond806_write_en = _guard12923;
assign cond806_clk = clk;
assign cond806_reset = reset;
assign cond806_in =
  _guard12924 ? idx_between_35_36_reg_out :
  1'd0;
assign cond809_write_en = _guard12925;
assign cond809_clk = clk;
assign cond809_reset = reset;
assign cond809_in =
  _guard12926 ? idx_between_20_36_reg_out :
  1'd0;
assign cond833_write_en = _guard12927;
assign cond833_clk = clk;
assign cond833_reset = reset;
assign cond833_in =
  _guard12928 ? idx_between_26_42_reg_out :
  1'd0;
assign cond_wire850_in =
  _guard12931 ? cond850_out :
  _guard12932 ? idx_between_46_47_reg_out :
  1'd0;
assign cond866_write_en = _guard12933;
assign cond866_clk = clk;
assign cond866_reset = reset;
assign cond866_in =
  _guard12934 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire872_in =
  _guard12935 ? idx_between_17_21_reg_out :
  _guard12938 ? cond872_out :
  1'd0;
assign cond887_write_en = _guard12939;
assign cond887_clk = clk;
assign cond887_reset = reset;
assign cond887_in =
  _guard12940 ? idx_between_40_41_reg_out :
  1'd0;
assign cond_wire888_in =
  _guard12943 ? cond888_out :
  _guard12944 ? idx_between_21_25_reg_out :
  1'd0;
assign cond889_write_en = _guard12945;
assign cond889_clk = clk;
assign cond889_reset = reset;
assign cond889_in =
  _guard12946 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire890_in =
  _guard12949 ? cond890_out :
  _guard12950 ? idx_between_25_41_reg_out :
  1'd0;
assign cond895_write_en = _guard12951;
assign cond895_clk = clk;
assign cond895_reset = reset;
assign cond895_in =
  _guard12952 ? idx_between_42_43_reg_out :
  1'd0;
assign cond_wire897_in =
  _guard12953 ? idx_between_23_39_reg_out :
  _guard12956 ? cond897_out :
  1'd0;
assign cond907_write_en = _guard12957;
assign cond907_clk = clk;
assign cond907_reset = reset;
assign cond907_in =
  _guard12958 ? idx_between_45_46_reg_out :
  1'd0;
assign cond909_write_en = _guard12959;
assign cond909_clk = clk;
assign cond909_reset = reset;
assign cond909_in =
  _guard12960 ? idx_between_26_42_reg_out :
  1'd0;
assign cond930_write_en = _guard12961;
assign cond930_clk = clk;
assign cond930_reset = reset;
assign cond930_in =
  _guard12962 ? idx_between_16_32_reg_out :
  1'd0;
assign cond_wire933_in =
  _guard12963 ? idx_between_17_21_reg_out :
  _guard12966 ? cond933_out :
  1'd0;
assign cond940_write_en = _guard12967;
assign cond940_clk = clk;
assign cond940_reset = reset;
assign cond940_in =
  _guard12968 ? idx_between_38_39_reg_out :
  1'd0;
assign cond941_write_en = _guard12969;
assign cond941_clk = clk;
assign cond941_reset = reset;
assign cond941_in =
  _guard12970 ? idx_between_19_23_reg_out :
  1'd0;
assign cond_wire958_in =
  _guard12971 ? idx_between_23_39_reg_out :
  _guard12974 ? cond958_out :
  1'd0;
assign cond960_write_en = _guard12975;
assign cond960_clk = clk;
assign cond960_reset = reset;
assign cond960_in =
  _guard12976 ? idx_between_43_44_reg_out :
  1'd0;
assign cond966_write_en = _guard12977;
assign cond966_clk = clk;
assign cond966_reset = reset;
assign cond966_in =
  _guard12978 ? idx_between_25_41_reg_out :
  1'd0;
assign cond984_write_en = _guard12979;
assign cond984_clk = clk;
assign cond984_reset = reset;
assign cond984_in =
  _guard12980 ? idx_between_49_50_reg_out :
  1'd0;
assign cond986_write_en = _guard12981;
assign cond986_clk = clk;
assign cond986_reset = reset;
assign cond986_in =
  _guard12982 ? idx_between_30_46_reg_out :
  1'd0;
assign cond_wire992_in =
  _guard12983 ? idx_between_20_36_reg_out :
  _guard12986 ? cond992_out :
  1'd0;
assign cond997_write_en = _guard12987;
assign cond997_clk = clk;
assign cond997_reset = reset;
assign cond997_in =
  _guard12988 ? idx_between_37_38_reg_out :
  1'd0;
assign cond_wire998_in =
  _guard12991 ? cond998_out :
  _guard12992 ? idx_between_18_22_reg_out :
  1'd0;
assign cond_wire1013_in =
  _guard12993 ? idx_between_41_42_reg_out :
  _guard12996 ? cond1013_out :
  1'd0;
assign cond_wire1022_in =
  _guard12999 ? cond1022_out :
  _guard13000 ? idx_between_24_28_reg_out :
  1'd0;
assign cond1040_write_en = _guard13001;
assign cond1040_clk = clk;
assign cond1040_reset = reset;
assign cond1040_in =
  _guard13002 ? idx_between_32_48_reg_out :
  1'd0;
assign cond_wire1049_in =
  _guard13005 ? cond1049_out :
  _guard13006 ? idx_between_50_51_reg_out :
  1'd0;
assign early_reset_static_par0_done_in = ud0_out;
assign left_0_7_write_en = _guard13009;
assign left_0_7_clk = clk;
assign left_0_7_reset = reset;
assign left_0_7_in = left_0_6_out;
assign top_0_14_write_en = _guard13015;
assign top_0_14_clk = clk;
assign top_0_14_reset = reset;
assign top_0_14_in = t14_read_data;
assign pe_1_12_mul_ready =
  _guard13021 ? 1'd1 :
  _guard13024 ? 1'd0 :
  1'd0;
assign pe_1_12_clk = clk;
assign pe_1_12_top =
  _guard13037 ? top_1_12_out :
  32'd0;
assign pe_1_12_left =
  _guard13050 ? left_1_12_out :
  32'd0;
assign pe_1_12_reset = reset;
assign pe_1_12_go = _guard13063;
assign pe_2_1_mul_ready =
  _guard13066 ? 1'd1 :
  _guard13069 ? 1'd0 :
  1'd0;
assign pe_2_1_clk = clk;
assign pe_2_1_top =
  _guard13082 ? top_2_1_out :
  32'd0;
assign pe_2_1_left =
  _guard13095 ? left_2_1_out :
  32'd0;
assign pe_2_1_reset = reset;
assign pe_2_1_go = _guard13108;
assign pe_2_3_mul_ready =
  _guard13111 ? 1'd1 :
  _guard13114 ? 1'd0 :
  1'd0;
assign pe_2_3_clk = clk;
assign pe_2_3_top =
  _guard13127 ? top_2_3_out :
  32'd0;
assign pe_2_3_left =
  _guard13140 ? left_2_3_out :
  32'd0;
assign pe_2_3_reset = reset;
assign pe_2_3_go = _guard13153;
assign pe_2_5_mul_ready =
  _guard13156 ? 1'd1 :
  _guard13159 ? 1'd0 :
  1'd0;
assign pe_2_5_clk = clk;
assign pe_2_5_top =
  _guard13172 ? top_2_5_out :
  32'd0;
assign pe_2_5_left =
  _guard13185 ? left_2_5_out :
  32'd0;
assign pe_2_5_reset = reset;
assign pe_2_5_go = _guard13198;
assign pe_3_1_mul_ready =
  _guard13201 ? 1'd1 :
  _guard13204 ? 1'd0 :
  1'd0;
assign pe_3_1_clk = clk;
assign pe_3_1_top =
  _guard13217 ? top_3_1_out :
  32'd0;
assign pe_3_1_left =
  _guard13230 ? left_3_1_out :
  32'd0;
assign pe_3_1_reset = reset;
assign pe_3_1_go = _guard13243;
assign top_3_4_write_en = _guard13246;
assign top_3_4_clk = clk;
assign top_3_4_reset = reset;
assign top_3_4_in = top_2_4_out;
assign pe_3_10_mul_ready =
  _guard13252 ? 1'd1 :
  _guard13255 ? 1'd0 :
  1'd0;
assign pe_3_10_clk = clk;
assign pe_3_10_top =
  _guard13268 ? top_3_10_out :
  32'd0;
assign pe_3_10_left =
  _guard13281 ? left_3_10_out :
  32'd0;
assign pe_3_10_reset = reset;
assign pe_3_10_go = _guard13294;
assign top_4_13_write_en = _guard13297;
assign top_4_13_clk = clk;
assign top_4_13_reset = reset;
assign top_4_13_in = top_3_13_out;
assign pe_4_14_mul_ready =
  _guard13303 ? 1'd1 :
  _guard13306 ? 1'd0 :
  1'd0;
assign pe_4_14_clk = clk;
assign pe_4_14_top =
  _guard13319 ? top_4_14_out :
  32'd0;
assign pe_4_14_left =
  _guard13332 ? left_4_14_out :
  32'd0;
assign pe_4_14_reset = reset;
assign pe_4_14_go = _guard13345;
assign pe_4_15_mul_ready =
  _guard13348 ? 1'd1 :
  _guard13351 ? 1'd0 :
  1'd0;
assign pe_4_15_clk = clk;
assign pe_4_15_top =
  _guard13364 ? top_4_15_out :
  32'd0;
assign pe_4_15_left =
  _guard13377 ? left_4_15_out :
  32'd0;
assign pe_4_15_reset = reset;
assign pe_4_15_go = _guard13390;
assign pe_5_3_mul_ready =
  _guard13393 ? 1'd1 :
  _guard13396 ? 1'd0 :
  1'd0;
assign pe_5_3_clk = clk;
assign pe_5_3_top =
  _guard13409 ? top_5_3_out :
  32'd0;
assign pe_5_3_left =
  _guard13422 ? left_5_3_out :
  32'd0;
assign pe_5_3_reset = reset;
assign pe_5_3_go = _guard13435;
assign pe_5_5_mul_ready =
  _guard13438 ? 1'd1 :
  _guard13441 ? 1'd0 :
  1'd0;
assign pe_5_5_clk = clk;
assign pe_5_5_top =
  _guard13454 ? top_5_5_out :
  32'd0;
assign pe_5_5_left =
  _guard13467 ? left_5_5_out :
  32'd0;
assign pe_5_5_reset = reset;
assign pe_5_5_go = _guard13480;
assign left_5_8_write_en = _guard13483;
assign left_5_8_clk = clk;
assign left_5_8_reset = reset;
assign left_5_8_in = left_5_7_out;
assign left_5_13_write_en = _guard13489;
assign left_5_13_clk = clk;
assign left_5_13_reset = reset;
assign left_5_13_in = left_5_12_out;
assign pe_6_2_mul_ready =
  _guard13495 ? 1'd1 :
  _guard13498 ? 1'd0 :
  1'd0;
assign pe_6_2_clk = clk;
assign pe_6_2_top =
  _guard13511 ? top_6_2_out :
  32'd0;
assign pe_6_2_left =
  _guard13524 ? left_6_2_out :
  32'd0;
assign pe_6_2_reset = reset;
assign pe_6_2_go = _guard13537;
assign pe_6_3_mul_ready =
  _guard13540 ? 1'd1 :
  _guard13543 ? 1'd0 :
  1'd0;
assign pe_6_3_clk = clk;
assign pe_6_3_top =
  _guard13556 ? top_6_3_out :
  32'd0;
assign pe_6_3_left =
  _guard13569 ? left_6_3_out :
  32'd0;
assign pe_6_3_reset = reset;
assign pe_6_3_go = _guard13582;
assign top_6_8_write_en = _guard13585;
assign top_6_8_clk = clk;
assign top_6_8_reset = reset;
assign top_6_8_in = top_5_8_out;
assign pe_6_10_mul_ready =
  _guard13591 ? 1'd1 :
  _guard13594 ? 1'd0 :
  1'd0;
assign pe_6_10_clk = clk;
assign pe_6_10_top =
  _guard13607 ? top_6_10_out :
  32'd0;
assign pe_6_10_left =
  _guard13620 ? left_6_10_out :
  32'd0;
assign pe_6_10_reset = reset;
assign pe_6_10_go = _guard13633;
assign left_6_13_write_en = _guard13636;
assign left_6_13_clk = clk;
assign left_6_13_reset = reset;
assign left_6_13_in = left_6_12_out;
assign left_7_1_write_en = _guard13642;
assign left_7_1_clk = clk;
assign left_7_1_reset = reset;
assign left_7_1_in = left_7_0_out;
assign left_7_3_write_en = _guard13648;
assign left_7_3_clk = clk;
assign left_7_3_reset = reset;
assign left_7_3_in = left_7_2_out;
assign top_7_5_write_en = _guard13654;
assign top_7_5_clk = clk;
assign top_7_5_reset = reset;
assign top_7_5_in = top_6_5_out;
assign pe_8_9_mul_ready =
  _guard13660 ? 1'd1 :
  _guard13663 ? 1'd0 :
  1'd0;
assign pe_8_9_clk = clk;
assign pe_8_9_top =
  _guard13676 ? top_8_9_out :
  32'd0;
assign pe_8_9_left =
  _guard13689 ? left_8_9_out :
  32'd0;
assign pe_8_9_reset = reset;
assign pe_8_9_go = _guard13702;
assign top_8_12_write_en = _guard13705;
assign top_8_12_clk = clk;
assign top_8_12_reset = reset;
assign top_8_12_in = top_7_12_out;
assign pe_8_15_mul_ready =
  _guard13711 ? 1'd1 :
  _guard13714 ? 1'd0 :
  1'd0;
assign pe_8_15_clk = clk;
assign pe_8_15_top =
  _guard13727 ? top_8_15_out :
  32'd0;
assign pe_8_15_left =
  _guard13740 ? left_8_15_out :
  32'd0;
assign pe_8_15_reset = reset;
assign pe_8_15_go = _guard13753;
assign top_9_6_write_en = _guard13756;
assign top_9_6_clk = clk;
assign top_9_6_reset = reset;
assign top_9_6_in = top_8_6_out;
assign top_9_9_write_en = _guard13762;
assign top_9_9_clk = clk;
assign top_9_9_reset = reset;
assign top_9_9_in = top_8_9_out;
assign pe_10_0_mul_ready =
  _guard13768 ? 1'd1 :
  _guard13771 ? 1'd0 :
  1'd0;
assign pe_10_0_clk = clk;
assign pe_10_0_top =
  _guard13784 ? top_10_0_out :
  32'd0;
assign pe_10_0_left =
  _guard13797 ? left_10_0_out :
  32'd0;
assign pe_10_0_reset = reset;
assign pe_10_0_go = _guard13810;
assign left_10_11_write_en = _guard13813;
assign left_10_11_clk = clk;
assign left_10_11_reset = reset;
assign left_10_11_in = left_10_10_out;
assign left_10_13_write_en = _guard13819;
assign left_10_13_clk = clk;
assign left_10_13_reset = reset;
assign left_10_13_in = left_10_12_out;
assign top_10_14_write_en = _guard13825;
assign top_10_14_clk = clk;
assign top_10_14_reset = reset;
assign top_10_14_in = top_9_14_out;
assign left_10_14_write_en = _guard13831;
assign left_10_14_clk = clk;
assign left_10_14_reset = reset;
assign left_10_14_in = left_10_13_out;
assign left_11_4_write_en = _guard13837;
assign left_11_4_clk = clk;
assign left_11_4_reset = reset;
assign left_11_4_in = left_11_3_out;
assign pe_11_9_mul_ready =
  _guard13843 ? 1'd1 :
  _guard13846 ? 1'd0 :
  1'd0;
assign pe_11_9_clk = clk;
assign pe_11_9_top =
  _guard13859 ? top_11_9_out :
  32'd0;
assign pe_11_9_left =
  _guard13872 ? left_11_9_out :
  32'd0;
assign pe_11_9_reset = reset;
assign pe_11_9_go = _guard13885;
assign left_11_9_write_en = _guard13888;
assign left_11_9_clk = clk;
assign left_11_9_reset = reset;
assign left_11_9_in = left_11_8_out;
assign left_11_11_write_en = _guard13894;
assign left_11_11_clk = clk;
assign left_11_11_reset = reset;
assign left_11_11_in = left_11_10_out;
assign left_11_12_write_en = _guard13900;
assign left_11_12_clk = clk;
assign left_11_12_reset = reset;
assign left_11_12_in = left_11_11_out;
assign left_12_11_write_en = _guard13906;
assign left_12_11_clk = clk;
assign left_12_11_reset = reset;
assign left_12_11_in = left_12_10_out;
assign left_13_0_write_en = _guard13912;
assign left_13_0_clk = clk;
assign left_13_0_reset = reset;
assign left_13_0_in = l13_read_data;
assign left_13_1_write_en = _guard13918;
assign left_13_1_clk = clk;
assign left_13_1_reset = reset;
assign left_13_1_in = left_13_0_out;
assign pe_13_5_mul_ready =
  _guard13924 ? 1'd1 :
  _guard13927 ? 1'd0 :
  1'd0;
assign pe_13_5_clk = clk;
assign pe_13_5_top =
  _guard13940 ? top_13_5_out :
  32'd0;
assign pe_13_5_left =
  _guard13953 ? left_13_5_out :
  32'd0;
assign pe_13_5_reset = reset;
assign pe_13_5_go = _guard13966;
assign pe_13_6_mul_ready =
  _guard13969 ? 1'd1 :
  _guard13972 ? 1'd0 :
  1'd0;
assign pe_13_6_clk = clk;
assign pe_13_6_top =
  _guard13985 ? top_13_6_out :
  32'd0;
assign pe_13_6_left =
  _guard13998 ? left_13_6_out :
  32'd0;
assign pe_13_6_reset = reset;
assign pe_13_6_go = _guard14011;
assign left_13_6_write_en = _guard14014;
assign left_13_6_clk = clk;
assign left_13_6_reset = reset;
assign left_13_6_in = left_13_5_out;
assign pe_13_8_mul_ready =
  _guard14020 ? 1'd1 :
  _guard14023 ? 1'd0 :
  1'd0;
assign pe_13_8_clk = clk;
assign pe_13_8_top =
  _guard14036 ? top_13_8_out :
  32'd0;
assign pe_13_8_left =
  _guard14049 ? left_13_8_out :
  32'd0;
assign pe_13_8_reset = reset;
assign pe_13_8_go = _guard14062;
assign pe_13_12_mul_ready =
  _guard14065 ? 1'd1 :
  _guard14068 ? 1'd0 :
  1'd0;
assign pe_13_12_clk = clk;
assign pe_13_12_top =
  _guard14081 ? top_13_12_out :
  32'd0;
assign pe_13_12_left =
  _guard14094 ? left_13_12_out :
  32'd0;
assign pe_13_12_reset = reset;
assign pe_13_12_go = _guard14107;
assign pe_14_4_mul_ready =
  _guard14110 ? 1'd1 :
  _guard14113 ? 1'd0 :
  1'd0;
assign pe_14_4_clk = clk;
assign pe_14_4_top =
  _guard14126 ? top_14_4_out :
  32'd0;
assign pe_14_4_left =
  _guard14139 ? left_14_4_out :
  32'd0;
assign pe_14_4_reset = reset;
assign pe_14_4_go = _guard14152;
assign left_14_6_write_en = _guard14155;
assign left_14_6_clk = clk;
assign left_14_6_reset = reset;
assign left_14_6_in = left_14_5_out;
assign pe_14_12_mul_ready =
  _guard14161 ? 1'd1 :
  _guard14164 ? 1'd0 :
  1'd0;
assign pe_14_12_clk = clk;
assign pe_14_12_top =
  _guard14177 ? top_14_12_out :
  32'd0;
assign pe_14_12_left =
  _guard14190 ? left_14_12_out :
  32'd0;
assign pe_14_12_reset = reset;
assign pe_14_12_go = _guard14203;
assign pe_14_15_mul_ready =
  _guard14206 ? 1'd1 :
  _guard14209 ? 1'd0 :
  1'd0;
assign pe_14_15_clk = clk;
assign pe_14_15_top =
  _guard14222 ? top_14_15_out :
  32'd0;
assign pe_14_15_left =
  _guard14235 ? left_14_15_out :
  32'd0;
assign pe_14_15_reset = reset;
assign pe_14_15_go = _guard14248;
assign pe_15_0_mul_ready =
  _guard14251 ? 1'd1 :
  _guard14254 ? 1'd0 :
  1'd0;
assign pe_15_0_clk = clk;
assign pe_15_0_top =
  _guard14267 ? top_15_0_out :
  32'd0;
assign pe_15_0_left =
  _guard14280 ? left_15_0_out :
  32'd0;
assign pe_15_0_reset = reset;
assign pe_15_0_go = _guard14293;
assign left_15_2_write_en = _guard14296;
assign left_15_2_clk = clk;
assign left_15_2_reset = reset;
assign left_15_2_in = left_15_1_out;
assign top_15_3_write_en = _guard14302;
assign top_15_3_clk = clk;
assign top_15_3_reset = reset;
assign top_15_3_in = top_14_3_out;
assign t4_add_left = 5'd1;
assign t4_add_right = t4_idx_out;
assign t5_idx_write_en = _guard14318;
assign t5_idx_clk = clk;
assign t5_idx_reset = reset;
assign t5_idx_in =
  _guard14321 ? 5'd0 :
  _guard14324 ? t5_add_out :
  'x;
assign t6_add_left = 5'd1;
assign t6_add_right = t6_idx_out;
assign t10_add_left = 5'd1;
assign t10_add_right = t10_idx_out;
assign t15_add_left = 5'd1;
assign t15_add_right = t15_idx_out;
assign l14_idx_write_en = _guard14349;
assign l14_idx_clk = clk;
assign l14_idx_reset = reset;
assign l14_idx_in =
  _guard14352 ? 5'd0 :
  _guard14355 ? l14_add_out :
  'x;
assign idx_between_35_51_reg_write_en = _guard14360;
assign idx_between_35_51_reg_clk = clk;
assign idx_between_35_51_reg_reset = reset;
assign idx_between_35_51_reg_in =
  _guard14361 ? idx_between_35_51_comb_out :
  _guard14364 ? 1'd0 :
  'x;
assign index_ge_17_left = idx_add_out;
assign index_ge_17_right = 6'd17;
assign idx_between_13_17_comb_left = index_ge_13_out;
assign idx_between_13_17_comb_right = index_lt_17_out;
assign idx_between_5_21_reg_write_en = _guard14373;
assign idx_between_5_21_reg_clk = clk;
assign idx_between_5_21_reg_reset = reset;
assign idx_between_5_21_reg_in =
  _guard14376 ? 1'd0 :
  _guard14377 ? idx_between_5_21_comb_out :
  'x;
assign index_lt_24_left = idx_add_out;
assign index_lt_24_right = 6'd24;
assign index_ge_29_left = idx_add_out;
assign index_ge_29_right = 6'd29;
assign idx_between_25_29_reg_write_en = _guard14386;
assign idx_between_25_29_reg_clk = clk;
assign idx_between_25_29_reg_reset = reset;
assign idx_between_25_29_reg_in =
  _guard14387 ? idx_between_25_29_comb_out :
  _guard14390 ? 1'd0 :
  'x;
assign idx_between_29_33_reg_write_en = _guard14395;
assign idx_between_29_33_reg_clk = clk;
assign idx_between_29_33_reg_reset = reset;
assign idx_between_29_33_reg_in =
  _guard14396 ? idx_between_29_33_comb_out :
  _guard14399 ? 1'd0 :
  'x;
assign idx_between_31_32_reg_write_en = _guard14404;
assign idx_between_31_32_reg_clk = clk;
assign idx_between_31_32_reg_reset = reset;
assign idx_between_31_32_reg_in =
  _guard14405 ? idx_between_31_32_comb_out :
  _guard14408 ? 1'd0 :
  'x;
assign idx_between_27_28_reg_write_en = _guard14413;
assign idx_between_27_28_reg_clk = clk;
assign idx_between_27_28_reg_reset = reset;
assign idx_between_27_28_reg_in =
  _guard14416 ? 1'd0 :
  _guard14417 ? idx_between_27_28_comb_out :
  'x;
assign idx_between_14_18_reg_write_en = _guard14422;
assign idx_between_14_18_reg_clk = clk;
assign idx_between_14_18_reg_reset = reset;
assign idx_between_14_18_reg_in =
  _guard14423 ? idx_between_14_18_comb_out :
  _guard14426 ? 1'd0 :
  'x;
assign idx_between_19_35_comb_left = index_ge_19_out;
assign idx_between_19_35_comb_right = index_lt_35_out;
assign idx_between_26_42_comb_left = index_ge_26_out;
assign idx_between_26_42_comb_right = index_lt_42_out;
assign idx_between_17_33_comb_left = index_ge_17_out;
assign idx_between_17_33_comb_right = index_lt_33_out;
assign idx_between_32_33_reg_write_en = _guard14437;
assign idx_between_32_33_reg_clk = clk;
assign idx_between_32_33_reg_reset = reset;
assign idx_between_32_33_reg_in =
  _guard14438 ? idx_between_32_33_comb_out :
  _guard14441 ? 1'd0 :
  'x;
assign idx_between_23_39_comb_left = index_ge_23_out;
assign idx_between_23_39_comb_right = index_lt_39_out;
assign cond17_write_en = _guard14444;
assign cond17_clk = clk;
assign cond17_reset = reset;
assign cond17_in =
  _guard14445 ? idx_between_8_24_reg_out :
  1'd0;
assign cond_wire22_in =
  _guard14446 ? idx_between_9_25_reg_out :
  _guard14449 ? cond22_out :
  1'd0;
assign cond23_write_en = _guard14450;
assign cond23_clk = clk;
assign cond23_reset = reset;
assign cond23_in =
  _guard14451 ? idx_between_25_26_reg_out :
  1'd0;
assign cond25_write_en = _guard14452;
assign cond25_clk = clk;
assign cond25_reset = reset;
assign cond25_in =
  _guard14453 ? idx_between_6_10_reg_out :
  1'd0;
assign cond_wire33_in =
  _guard14454 ? idx_between_27_28_reg_out :
  _guard14457 ? cond33_out :
  1'd0;
assign cond52_write_en = _guard14458;
assign cond52_clk = clk;
assign cond52_reset = reset;
assign cond52_in =
  _guard14459 ? idx_between_15_31_reg_out :
  1'd0;
assign cond56_write_en = _guard14460;
assign cond56_clk = clk;
assign cond56_reset = reset;
assign cond56_in =
  _guard14461 ? idx_between_12_28_reg_out :
  1'd0;
assign cond58_write_en = _guard14462;
assign cond58_clk = clk;
assign cond58_reset = reset;
assign cond58_in =
  _guard14463 ? idx_between_32_33_reg_out :
  1'd0;
assign cond75_write_en = _guard14464;
assign cond75_clk = clk;
assign cond75_reset = reset;
assign cond75_in =
  _guard14465 ? idx_between_16_20_reg_out :
  1'd0;
assign cond88_write_en = _guard14466;
assign cond88_clk = clk;
assign cond88_reset = reset;
assign cond88_in =
  _guard14467 ? idx_between_4_8_reg_out :
  1'd0;
assign cond93_write_en = _guard14468;
assign cond93_clk = clk;
assign cond93_reset = reset;
assign cond93_in =
  _guard14469 ? idx_between_5_21_reg_out :
  1'd0;
assign cond_wire98_in =
  _guard14472 ? cond98_out :
  _guard14473 ? idx_between_10_26_reg_out :
  1'd0;
assign cond_wire106_in =
  _guard14476 ? cond106_out :
  _guard14477 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire120_in =
  _guard14478 ? idx_between_12_16_reg_out :
  _guard14481 ? cond120_out :
  1'd0;
assign cond124_write_en = _guard14482;
assign cond124_clk = clk;
assign cond124_reset = reset;
assign cond124_in =
  _guard14483 ? idx_between_13_17_reg_out :
  1'd0;
assign cond137_write_en = _guard14484;
assign cond137_clk = clk;
assign cond137_reset = reset;
assign cond137_in =
  _guard14485 ? idx_between_16_32_reg_out :
  1'd0;
assign cond155_write_en = _guard14486;
assign cond155_clk = clk;
assign cond155_reset = reset;
assign cond155_in =
  _guard14487 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire176_in =
  _guard14490 ? cond176_out :
  _guard14491 ? idx_between_30_31_reg_out :
  1'd0;
assign cond188_write_en = _guard14492;
assign cond188_clk = clk;
assign cond188_reset = reset;
assign cond188_in =
  _guard14493 ? idx_between_33_34_reg_out :
  1'd0;
assign cond209_write_en = _guard14494;
assign cond209_clk = clk;
assign cond209_reset = reset;
assign cond209_in =
  _guard14495 ? idx_between_3_19_reg_out :
  1'd0;
assign cond_wire213_in =
  _guard14496 ? idx_between_24_25_reg_out :
  _guard14499 ? cond213_out :
  1'd0;
assign cond220_write_en = _guard14500;
assign cond220_clk = clk;
assign cond220_reset = reset;
assign cond220_in =
  _guard14501 ? idx_between_10_26_reg_out :
  1'd0;
assign cond_wire221_in =
  _guard14502 ? idx_between_26_27_reg_out :
  _guard14505 ? cond221_out :
  1'd0;
assign cond228_write_en = _guard14506;
assign cond228_clk = clk;
assign cond228_reset = reset;
assign cond228_in =
  _guard14507 ? idx_between_12_28_reg_out :
  1'd0;
assign cond232_write_en = _guard14508;
assign cond232_clk = clk;
assign cond232_reset = reset;
assign cond232_in =
  _guard14509 ? idx_between_13_29_reg_out :
  1'd0;
assign cond_wire236_in =
  _guard14512 ? cond236_out :
  _guard14513 ? idx_between_14_30_reg_out :
  1'd0;
assign cond258_write_en = _guard14514;
assign cond258_clk = clk;
assign cond258_reset = reset;
assign cond258_in =
  _guard14515 ? idx_between_16_20_reg_out :
  1'd0;
assign cond262_write_en = _guard14516;
assign cond262_clk = clk;
assign cond262_reset = reset;
assign cond262_in =
  _guard14517 ? idx_between_17_21_reg_out :
  1'd0;
assign cond_wire270_in =
  _guard14518 ? idx_between_19_23_reg_out :
  _guard14521 ? cond270_out :
  1'd0;
assign cond272_write_en = _guard14522;
assign cond272_clk = clk;
assign cond272_reset = reset;
assign cond272_in =
  _guard14523 ? idx_between_23_39_reg_out :
  1'd0;
assign cond_wire278_in =
  _guard14524 ? idx_between_25_26_reg_out :
  _guard14527 ? cond278_out :
  1'd0;
assign cond_wire303_in =
  _guard14528 ? idx_between_12_16_reg_out :
  _guard14531 ? cond303_out :
  1'd0;
assign cond311_write_en = _guard14532;
assign cond311_clk = clk;
assign cond311_reset = reset;
assign cond311_in =
  _guard14533 ? idx_between_14_18_reg_out :
  1'd0;
assign cond_wire312_in =
  _guard14534 ? idx_between_14_30_reg_out :
  _guard14537 ? cond312_out :
  1'd0;
assign cond320_write_en = _guard14538;
assign cond320_clk = clk;
assign cond320_reset = reset;
assign cond320_in =
  _guard14539 ? idx_between_16_32_reg_out :
  1'd0;
assign cond323_write_en = _guard14540;
assign cond323_clk = clk;
assign cond323_reset = reset;
assign cond323_in =
  _guard14541 ? idx_between_17_21_reg_out :
  1'd0;
assign cond_wire323_in =
  _guard14542 ? idx_between_17_21_reg_out :
  _guard14545 ? cond323_out :
  1'd0;
assign cond_wire330_in =
  _guard14548 ? cond330_out :
  _guard14549 ? idx_between_38_39_reg_out :
  1'd0;
assign cond331_write_en = _guard14550;
assign cond331_clk = clk;
assign cond331_reset = reset;
assign cond331_in =
  _guard14551 ? idx_between_19_23_reg_out :
  1'd0;
assign cond_wire332_in =
  _guard14554 ? cond332_out :
  _guard14555 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire358_in =
  _guard14556 ? idx_between_14_30_reg_out :
  _guard14559 ? cond358_out :
  1'd0;
assign cond_wire365_in =
  _guard14560 ? idx_between_12_28_reg_out :
  _guard14563 ? cond365_out :
  1'd0;
assign cond369_write_en = _guard14564;
assign cond369_clk = clk;
assign cond369_reset = reset;
assign cond369_in =
  _guard14565 ? idx_between_13_29_reg_out :
  1'd0;
assign cond379_write_en = _guard14566;
assign cond379_clk = clk;
assign cond379_reset = reset;
assign cond379_in =
  _guard14567 ? idx_between_35_36_reg_out :
  1'd0;
assign cond414_write_en = _guard14568;
assign cond414_clk = clk;
assign cond414_reset = reset;
assign cond414_in =
  _guard14569 ? idx_between_9_25_reg_out :
  1'd0;
assign cond415_write_en = _guard14570;
assign cond415_clk = clk;
assign cond415_reset = reset;
assign cond415_in =
  _guard14571 ? idx_between_13_29_reg_out :
  1'd0;
assign cond_wire415_in =
  _guard14572 ? idx_between_13_29_reg_out :
  _guard14575 ? cond415_out :
  1'd0;
assign cond_wire416_in =
  _guard14578 ? cond416_out :
  _guard14579 ? idx_between_29_30_reg_out :
  1'd0;
assign cond_wire423_in =
  _guard14582 ? cond423_out :
  _guard14583 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire430_in =
  _guard14584 ? idx_between_13_29_reg_out :
  _guard14587 ? cond430_out :
  1'd0;
assign cond_wire432_in =
  _guard14590 ? cond432_out :
  _guard14591 ? idx_between_33_34_reg_out :
  1'd0;
assign cond_wire449_in =
  _guard14594 ? cond449_out :
  _guard14595 ? idx_between_18_22_reg_out :
  1'd0;
assign cond_wire451_in =
  _guard14598 ? cond451_out :
  _guard14599 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire453_in =
  _guard14600 ? idx_between_19_23_reg_out :
  _guard14603 ? cond453_out :
  1'd0;
assign cond_wire461_in =
  _guard14604 ? idx_between_21_25_reg_out :
  _guard14607 ? cond461_out :
  1'd0;
assign cond462_write_en = _guard14608;
assign cond462_clk = clk;
assign cond462_reset = reset;
assign cond462_in =
  _guard14609 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire466_in =
  _guard14612 ? cond466_out :
  _guard14613 ? idx_between_22_38_reg_out :
  1'd0;
assign cond484_write_en = _guard14614;
assign cond484_clk = clk;
assign cond484_reset = reset;
assign cond484_in =
  _guard14615 ? idx_between_15_31_reg_out :
  1'd0;
assign cond488_write_en = _guard14616;
assign cond488_clk = clk;
assign cond488_reset = reset;
assign cond488_in =
  _guard14617 ? idx_between_16_32_reg_out :
  1'd0;
assign cond_wire493_in =
  _guard14618 ? idx_between_33_34_reg_out :
  _guard14621 ? cond493_out :
  1'd0;
assign cond496_write_en = _guard14622;
assign cond496_clk = clk;
assign cond496_reset = reset;
assign cond496_in =
  _guard14623 ? idx_between_18_34_reg_out :
  1'd0;
assign cond_wire497_in =
  _guard14624 ? idx_between_34_35_reg_out :
  _guard14627 ? cond497_out :
  1'd0;
assign cond500_write_en = _guard14628;
assign cond500_clk = clk;
assign cond500_reset = reset;
assign cond500_in =
  _guard14629 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire503_in =
  _guard14630 ? idx_between_16_32_reg_out :
  _guard14633 ? cond503_out :
  1'd0;
assign cond510_write_en = _guard14634;
assign cond510_clk = clk;
assign cond510_reset = reset;
assign cond510_in =
  _guard14635 ? idx_between_18_22_reg_out :
  1'd0;
assign cond511_write_en = _guard14636;
assign cond511_clk = clk;
assign cond511_reset = reset;
assign cond511_in =
  _guard14637 ? idx_between_18_34_reg_out :
  1'd0;
assign cond532_write_en = _guard14638;
assign cond532_clk = clk;
assign cond532_reset = reset;
assign cond532_in =
  _guard14639 ? idx_between_27_43_reg_out :
  1'd0;
assign cond533_write_en = _guard14640;
assign cond533_clk = clk;
assign cond533_reset = reset;
assign cond533_in =
  _guard14641 ? idx_between_43_44_reg_out :
  1'd0;
assign cond551_write_en = _guard14642;
assign cond551_clk = clk;
assign cond551_reset = reset;
assign cond551_in =
  _guard14643 ? idx_between_13_17_reg_out :
  1'd0;
assign cond_wire561_in =
  _guard14646 ? cond561_out :
  _guard14647 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire566_in =
  _guard14648 ? idx_between_36_37_reg_out :
  _guard14651 ? cond566_out :
  1'd0;
assign cond569_write_en = _guard14652;
assign cond569_clk = clk;
assign cond569_reset = reset;
assign cond569_in =
  _guard14653 ? idx_between_21_37_reg_out :
  1'd0;
assign cond582_write_en = _guard14654;
assign cond582_clk = clk;
assign cond582_reset = reset;
assign cond582_in =
  _guard14655 ? idx_between_40_41_reg_out :
  1'd0;
assign cond594_write_en = _guard14656;
assign cond594_clk = clk;
assign cond594_reset = reset;
assign cond594_in =
  _guard14657 ? idx_between_43_44_reg_out :
  1'd0;
assign cond596_write_en = _guard14658;
assign cond596_clk = clk;
assign cond596_reset = reset;
assign cond596_in =
  _guard14659 ? idx_between_24_40_reg_out :
  1'd0;
assign cond603_write_en = _guard14660;
assign cond603_clk = clk;
assign cond603_reset = reset;
assign cond603_in =
  _guard14661 ? idx_between_30_31_reg_out :
  1'd0;
assign cond610_write_en = _guard14662;
assign cond610_clk = clk;
assign cond610_reset = reset;
assign cond610_in =
  _guard14663 ? idx_between_16_32_reg_out :
  1'd0;
assign cond_wire611_in =
  _guard14664 ? idx_between_32_33_reg_out :
  _guard14667 ? cond611_out :
  1'd0;
assign cond_wire618_in =
  _guard14668 ? idx_between_18_34_reg_out :
  _guard14671 ? cond618_out :
  1'd0;
assign cond634_write_en = _guard14672;
assign cond634_clk = clk;
assign cond634_reset = reset;
assign cond634_in =
  _guard14673 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire640_in =
  _guard14674 ? idx_between_20_24_reg_out :
  _guard14677 ? cond640_out :
  1'd0;
assign cond648_write_en = _guard14678;
assign cond648_clk = clk;
assign cond648_reset = reset;
assign cond648_in =
  _guard14679 ? idx_between_22_26_reg_out :
  1'd0;
assign cond_wire657_in =
  _guard14682 ? cond657_out :
  _guard14683 ? idx_between_24_40_reg_out :
  1'd0;
assign cond662_write_en = _guard14684;
assign cond662_clk = clk;
assign cond662_reset = reset;
assign cond662_in =
  _guard14685 ? idx_between_29_45_reg_out :
  1'd0;
assign cond668_write_en = _guard14686;
assign cond668_clk = clk;
assign cond668_reset = reset;
assign cond668_in =
  _guard14687 ? idx_between_31_32_reg_out :
  1'd0;
assign cond_wire672_in =
  _guard14688 ? idx_between_32_33_reg_out :
  _guard14691 ? cond672_out :
  1'd0;
assign cond674_write_en = _guard14692;
assign cond674_clk = clk;
assign cond674_reset = reset;
assign cond674_in =
  _guard14693 ? idx_between_13_29_reg_out :
  1'd0;
assign cond682_write_en = _guard14694;
assign cond682_clk = clk;
assign cond682_reset = reset;
assign cond682_in =
  _guard14695 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire703_in =
  _guard14696 ? idx_between_24_40_reg_out :
  _guard14699 ? cond703_out :
  1'd0;
assign cond709_write_en = _guard14700;
assign cond709_clk = clk;
assign cond709_reset = reset;
assign cond709_in =
  _guard14701 ? idx_between_22_26_reg_out :
  1'd0;
assign cond_wire715_in =
  _guard14704 ? cond715_out :
  _guard14705 ? idx_between_27_43_reg_out :
  1'd0;
assign cond_wire739_in =
  _guard14706 ? idx_between_14_30_reg_out :
  _guard14709 ? cond739_out :
  1'd0;
assign cond_wire764_in =
  _guard14712 ? cond764_out :
  _guard14713 ? idx_between_24_40_reg_out :
  1'd0;
assign cond_wire769_in =
  _guard14716 ? cond769_out :
  _guard14717 ? idx_between_41_42_reg_out :
  1'd0;
assign cond774_write_en = _guard14718;
assign cond774_clk = clk;
assign cond774_reset = reset;
assign cond774_in =
  _guard14719 ? idx_between_23_27_reg_out :
  1'd0;
assign cond_wire784_in =
  _guard14722 ? cond784_out :
  _guard14723 ? idx_between_29_45_reg_out :
  1'd0;
assign cond785_write_en = _guard14724;
assign cond785_clk = clk;
assign cond785_reset = reset;
assign cond785_in =
  _guard14725 ? idx_between_45_46_reg_out :
  1'd0;
assign cond_wire787_in =
  _guard14728 ? cond787_out :
  _guard14729 ? idx_between_26_42_reg_out :
  1'd0;
assign cond790_write_en = _guard14730;
assign cond790_clk = clk;
assign cond790_reset = reset;
assign cond790_in =
  _guard14731 ? idx_between_27_31_reg_out :
  1'd0;
assign cond794_write_en = _guard14732;
assign cond794_clk = clk;
assign cond794_reset = reset;
assign cond794_in =
  _guard14733 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire805_in =
  _guard14736 ? cond805_out :
  _guard14737 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire817_in =
  _guard14740 ? cond817_out :
  _guard14741 ? idx_between_22_38_reg_out :
  1'd0;
assign cond830_write_en = _guard14742;
assign cond830_clk = clk;
assign cond830_reset = reset;
assign cond830_in =
  _guard14743 ? idx_between_41_42_reg_out :
  1'd0;
assign cond_wire833_in =
  _guard14746 ? cond833_out :
  _guard14747 ? idx_between_26_42_reg_out :
  1'd0;
assign cond841_write_en = _guard14748;
assign cond841_clk = clk;
assign cond841_reset = reset;
assign cond841_in =
  _guard14749 ? idx_between_28_44_reg_out :
  1'd0;
assign cond851_write_en = _guard14750;
assign cond851_clk = clk;
assign cond851_reset = reset;
assign cond851_in =
  _guard14751 ? idx_between_27_31_reg_out :
  1'd0;
assign cond_wire858_in =
  _guard14754 ? cond858_out :
  _guard14755 ? idx_between_48_49_reg_out :
  1'd0;
assign cond860_write_en = _guard14756;
assign cond860_clk = clk;
assign cond860_reset = reset;
assign cond860_in =
  _guard14757 ? idx_between_14_18_reg_out :
  1'd0;
assign cond_wire860_in =
  _guard14758 ? idx_between_14_18_reg_out :
  _guard14761 ? cond860_out :
  1'd0;
assign cond863_write_en = _guard14762;
assign cond863_clk = clk;
assign cond863_reset = reset;
assign cond863_in =
  _guard14763 ? idx_between_34_35_reg_out :
  1'd0;
assign cond865_write_en = _guard14764;
assign cond865_clk = clk;
assign cond865_reset = reset;
assign cond865_in =
  _guard14765 ? idx_between_15_31_reg_out :
  1'd0;
assign cond871_write_en = _guard14766;
assign cond871_clk = clk;
assign cond871_reset = reset;
assign cond871_in =
  _guard14767 ? idx_between_36_37_reg_out :
  1'd0;
assign cond_wire874_in =
  _guard14770 ? cond874_out :
  _guard14771 ? idx_between_21_37_reg_out :
  1'd0;
assign cond878_write_en = _guard14772;
assign cond878_clk = clk;
assign cond878_reset = reset;
assign cond878_in =
  _guard14773 ? idx_between_22_38_reg_out :
  1'd0;
assign cond892_write_en = _guard14774;
assign cond892_clk = clk;
assign cond892_reset = reset;
assign cond892_in =
  _guard14775 ? idx_between_22_26_reg_out :
  1'd0;
assign cond893_write_en = _guard14776;
assign cond893_clk = clk;
assign cond893_reset = reset;
assign cond893_in =
  _guard14777 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire910_in =
  _guard14778 ? idx_between_30_46_reg_out :
  _guard14781 ? cond910_out :
  1'd0;
assign cond_wire912_in =
  _guard14784 ? cond912_out :
  _guard14785 ? idx_between_27_31_reg_out :
  1'd0;
assign cond_wire917_in =
  _guard14788 ? cond917_out :
  _guard14789 ? idx_between_28_44_reg_out :
  1'd0;
assign cond_wire918_in =
  _guard14792 ? cond918_out :
  _guard14793 ? idx_between_32_48_reg_out :
  1'd0;
assign cond922_write_en = _guard14794;
assign cond922_clk = clk;
assign cond922_reset = reset;
assign cond922_in =
  _guard14795 ? idx_between_33_49_reg_out :
  1'd0;
assign cond923_write_en = _guard14796;
assign cond923_clk = clk;
assign cond923_reset = reset;
assign cond923_in =
  _guard14797 ? idx_between_49_50_reg_out :
  1'd0;
assign cond929_write_en = _guard14798;
assign cond929_clk = clk;
assign cond929_reset = reset;
assign cond929_in =
  _guard14799 ? idx_between_16_20_reg_out :
  1'd0;
assign cond_wire934_in =
  _guard14800 ? idx_between_17_33_reg_out :
  _guard14803 ? cond934_out :
  1'd0;
assign cond936_write_en = _guard14804;
assign cond936_clk = clk;
assign cond936_reset = reset;
assign cond936_in =
  _guard14805 ? idx_between_37_38_reg_out :
  1'd0;
assign cond_wire936_in =
  _guard14808 ? cond936_out :
  _guard14809 ? idx_between_37_38_reg_out :
  1'd0;
assign cond939_write_en = _guard14810;
assign cond939_clk = clk;
assign cond939_reset = reset;
assign cond939_in =
  _guard14811 ? idx_between_22_38_reg_out :
  1'd0;
assign cond958_write_en = _guard14812;
assign cond958_clk = clk;
assign cond958_reset = reset;
assign cond958_in =
  _guard14813 ? idx_between_23_39_reg_out :
  1'd0;
assign cond972_write_en = _guard14814;
assign cond972_clk = clk;
assign cond972_reset = reset;
assign cond972_in =
  _guard14815 ? idx_between_46_47_reg_out :
  1'd0;
assign cond_wire990_in =
  _guard14816 ? idx_between_16_20_reg_out :
  _guard14819 ? cond990_out :
  1'd0;
assign cond991_write_en = _guard14820;
assign cond991_clk = clk;
assign cond991_reset = reset;
assign cond991_in =
  _guard14821 ? idx_between_16_32_reg_out :
  1'd0;
assign cond_wire995_in =
  _guard14822 ? idx_between_17_33_reg_out :
  _guard14825 ? cond995_out :
  1'd0;
assign cond_wire1002_in =
  _guard14826 ? idx_between_19_23_reg_out :
  _guard14829 ? cond1002_out :
  1'd0;
assign cond1016_write_en = _guard14830;
assign cond1016_clk = clk;
assign cond1016_reset = reset;
assign cond1016_in =
  _guard14831 ? idx_between_26_42_reg_out :
  1'd0;
assign cond_wire1020_in =
  _guard14832 ? idx_between_27_43_reg_out :
  _guard14835 ? cond1020_out :
  1'd0;
assign cond1021_write_en = _guard14836;
assign cond1021_clk = clk;
assign cond1021_reset = reset;
assign cond1021_in =
  _guard14837 ? idx_between_43_44_reg_out :
  1'd0;
assign cond1033_write_en = _guard14838;
assign cond1033_clk = clk;
assign cond1033_reset = reset;
assign cond1033_in =
  _guard14839 ? idx_between_46_47_reg_out :
  1'd0;
assign cond_wire1037_in =
  _guard14842 ? cond1037_out :
  _guard14843 ? idx_between_47_48_reg_out :
  1'd0;
assign cond_wire1039_in =
  _guard14846 ? cond1039_out :
  _guard14847 ? idx_between_28_44_reg_out :
  1'd0;
assign cond1050_write_en = _guard14848;
assign cond1050_clk = clk;
assign cond1050_reset = reset;
assign cond1050_in =
  _guard14849 ? idx_between_31_35_reg_out :
  1'd0;
assign fsm0_write_en = _guard14850;
assign fsm0_clk = clk;
assign fsm0_reset = reset;
assign fsm0_in =
  _guard14853 ? adder_out :
  _guard14856 ? 6'd0 :
  6'd0;
assign left_0_9_write_en = _guard14859;
assign left_0_9_clk = clk;
assign left_0_9_reset = reset;
assign left_0_9_in = left_0_8_out;
assign pe_1_5_mul_ready =
  _guard14865 ? 1'd1 :
  _guard14868 ? 1'd0 :
  1'd0;
assign pe_1_5_clk = clk;
assign pe_1_5_top =
  _guard14881 ? top_1_5_out :
  32'd0;
assign pe_1_5_left =
  _guard14894 ? left_1_5_out :
  32'd0;
assign pe_1_5_reset = reset;
assign pe_1_5_go = _guard14907;
assign top_1_6_write_en = _guard14910;
assign top_1_6_clk = clk;
assign top_1_6_reset = reset;
assign top_1_6_in = top_0_6_out;
assign left_1_10_write_en = _guard14916;
assign left_1_10_clk = clk;
assign left_1_10_reset = reset;
assign left_1_10_in = left_1_9_out;
assign top_1_11_write_en = _guard14922;
assign top_1_11_clk = clk;
assign top_1_11_reset = reset;
assign top_1_11_in = top_0_11_out;
assign top_2_0_write_en = _guard14928;
assign top_2_0_clk = clk;
assign top_2_0_reset = reset;
assign top_2_0_in = top_1_0_out;
assign left_2_12_write_en = _guard14934;
assign left_2_12_clk = clk;
assign left_2_12_reset = reset;
assign left_2_12_in = left_2_11_out;
assign top_3_0_write_en = _guard14940;
assign top_3_0_clk = clk;
assign top_3_0_reset = reset;
assign top_3_0_in = top_2_0_out;
assign top_3_1_write_en = _guard14946;
assign top_3_1_clk = clk;
assign top_3_1_reset = reset;
assign top_3_1_in = top_2_1_out;
assign top_3_9_write_en = _guard14952;
assign top_3_9_clk = clk;
assign top_3_9_reset = reset;
assign top_3_9_in = top_2_9_out;
assign top_3_10_write_en = _guard14958;
assign top_3_10_clk = clk;
assign top_3_10_reset = reset;
assign top_3_10_in = top_2_10_out;
assign top_3_15_write_en = _guard14964;
assign top_3_15_clk = clk;
assign top_3_15_reset = reset;
assign top_3_15_in = top_2_15_out;
assign pe_4_6_mul_ready =
  _guard14970 ? 1'd1 :
  _guard14973 ? 1'd0 :
  1'd0;
assign pe_4_6_clk = clk;
assign pe_4_6_top =
  _guard14986 ? top_4_6_out :
  32'd0;
assign pe_4_6_left =
  _guard14999 ? left_4_6_out :
  32'd0;
assign pe_4_6_reset = reset;
assign pe_4_6_go = _guard15012;
assign left_4_10_write_en = _guard15015;
assign left_4_10_clk = clk;
assign left_4_10_reset = reset;
assign left_4_10_in = left_4_9_out;
assign pe_4_11_mul_ready =
  _guard15021 ? 1'd1 :
  _guard15024 ? 1'd0 :
  1'd0;
assign pe_4_11_clk = clk;
assign pe_4_11_top =
  _guard15037 ? top_4_11_out :
  32'd0;
assign pe_4_11_left =
  _guard15050 ? left_4_11_out :
  32'd0;
assign pe_4_11_reset = reset;
assign pe_4_11_go = _guard15063;
assign top_5_2_write_en = _guard15066;
assign top_5_2_clk = clk;
assign top_5_2_reset = reset;
assign top_5_2_in = top_4_2_out;
assign top_5_4_write_en = _guard15072;
assign top_5_4_clk = clk;
assign top_5_4_reset = reset;
assign top_5_4_in = top_4_4_out;
assign left_5_10_write_en = _guard15078;
assign left_5_10_clk = clk;
assign left_5_10_reset = reset;
assign left_5_10_in = left_5_9_out;
assign top_5_13_write_en = _guard15084;
assign top_5_13_clk = clk;
assign top_5_13_reset = reset;
assign top_5_13_in = top_4_13_out;
assign top_6_14_write_en = _guard15090;
assign top_6_14_clk = clk;
assign top_6_14_reset = reset;
assign top_6_14_in = top_5_14_out;
assign left_6_14_write_en = _guard15096;
assign left_6_14_clk = clk;
assign left_6_14_reset = reset;
assign left_6_14_in = left_6_13_out;
assign left_6_15_write_en = _guard15102;
assign left_6_15_clk = clk;
assign left_6_15_reset = reset;
assign left_6_15_in = left_6_14_out;
assign left_7_7_write_en = _guard15108;
assign left_7_7_clk = clk;
assign left_7_7_reset = reset;
assign left_7_7_in = left_7_6_out;
assign left_8_9_write_en = _guard15114;
assign left_8_9_clk = clk;
assign left_8_9_reset = reset;
assign left_8_9_in = left_8_8_out;
assign left_8_12_write_en = _guard15120;
assign left_8_12_clk = clk;
assign left_8_12_reset = reset;
assign left_8_12_in = left_8_11_out;
assign top_8_13_write_en = _guard15126;
assign top_8_13_clk = clk;
assign top_8_13_reset = reset;
assign top_8_13_in = top_7_13_out;
assign pe_9_10_mul_ready =
  _guard15132 ? 1'd1 :
  _guard15135 ? 1'd0 :
  1'd0;
assign pe_9_10_clk = clk;
assign pe_9_10_top =
  _guard15148 ? top_9_10_out :
  32'd0;
assign pe_9_10_left =
  _guard15161 ? left_9_10_out :
  32'd0;
assign pe_9_10_reset = reset;
assign pe_9_10_go = _guard15174;
assign pe_9_12_mul_ready =
  _guard15177 ? 1'd1 :
  _guard15180 ? 1'd0 :
  1'd0;
assign pe_9_12_clk = clk;
assign pe_9_12_top =
  _guard15193 ? top_9_12_out :
  32'd0;
assign pe_9_12_left =
  _guard15206 ? left_9_12_out :
  32'd0;
assign pe_9_12_reset = reset;
assign pe_9_12_go = _guard15219;
assign top_10_1_write_en = _guard15222;
assign top_10_1_clk = clk;
assign top_10_1_reset = reset;
assign top_10_1_in = top_9_1_out;
assign pe_10_14_mul_ready =
  _guard15228 ? 1'd1 :
  _guard15231 ? 1'd0 :
  1'd0;
assign pe_10_14_clk = clk;
assign pe_10_14_top =
  _guard15244 ? top_10_14_out :
  32'd0;
assign pe_10_14_left =
  _guard15257 ? left_10_14_out :
  32'd0;
assign pe_10_14_reset = reset;
assign pe_10_14_go = _guard15270;
assign left_10_15_write_en = _guard15273;
assign left_10_15_clk = clk;
assign left_10_15_reset = reset;
assign left_10_15_in = left_10_14_out;
assign pe_11_2_mul_ready =
  _guard15279 ? 1'd1 :
  _guard15282 ? 1'd0 :
  1'd0;
assign pe_11_2_clk = clk;
assign pe_11_2_top =
  _guard15295 ? top_11_2_out :
  32'd0;
assign pe_11_2_left =
  _guard15308 ? left_11_2_out :
  32'd0;
assign pe_11_2_reset = reset;
assign pe_11_2_go = _guard15321;
assign top_11_2_write_en = _guard15324;
assign top_11_2_clk = clk;
assign top_11_2_reset = reset;
assign top_11_2_in = top_10_2_out;
assign pe_11_3_mul_ready =
  _guard15330 ? 1'd1 :
  _guard15333 ? 1'd0 :
  1'd0;
assign pe_11_3_clk = clk;
assign pe_11_3_top =
  _guard15346 ? top_11_3_out :
  32'd0;
assign pe_11_3_left =
  _guard15359 ? left_11_3_out :
  32'd0;
assign pe_11_3_reset = reset;
assign pe_11_3_go = _guard15372;
assign top_11_6_write_en = _guard15375;
assign top_11_6_clk = clk;
assign top_11_6_reset = reset;
assign top_11_6_in = top_10_6_out;
assign top_11_14_write_en = _guard15381;
assign top_11_14_clk = clk;
assign top_11_14_reset = reset;
assign top_11_14_in = top_10_14_out;
assign left_12_3_write_en = _guard15387;
assign left_12_3_clk = clk;
assign left_12_3_reset = reset;
assign left_12_3_in = left_12_2_out;
assign top_12_13_write_en = _guard15393;
assign top_12_13_clk = clk;
assign top_12_13_reset = reset;
assign top_12_13_in = top_11_13_out;
assign pe_13_1_mul_ready =
  _guard15399 ? 1'd1 :
  _guard15402 ? 1'd0 :
  1'd0;
assign pe_13_1_clk = clk;
assign pe_13_1_top =
  _guard15415 ? top_13_1_out :
  32'd0;
assign pe_13_1_left =
  _guard15428 ? left_13_1_out :
  32'd0;
assign pe_13_1_reset = reset;
assign pe_13_1_go = _guard15441;
assign top_13_1_write_en = _guard15444;
assign top_13_1_clk = clk;
assign top_13_1_reset = reset;
assign top_13_1_in = top_12_1_out;
assign pe_14_0_mul_ready =
  _guard15450 ? 1'd1 :
  _guard15453 ? 1'd0 :
  1'd0;
assign pe_14_0_clk = clk;
assign pe_14_0_top =
  _guard15466 ? top_14_0_out :
  32'd0;
assign pe_14_0_left =
  _guard15479 ? left_14_0_out :
  32'd0;
assign pe_14_0_reset = reset;
assign pe_14_0_go = _guard15492;
assign pe_14_5_mul_ready =
  _guard15495 ? 1'd1 :
  _guard15498 ? 1'd0 :
  1'd0;
assign pe_14_5_clk = clk;
assign pe_14_5_top =
  _guard15511 ? top_14_5_out :
  32'd0;
assign pe_14_5_left =
  _guard15524 ? left_14_5_out :
  32'd0;
assign pe_14_5_reset = reset;
assign pe_14_5_go = _guard15537;
assign top_14_5_write_en = _guard15540;
assign top_14_5_clk = clk;
assign top_14_5_reset = reset;
assign top_14_5_in = top_13_5_out;
assign left_15_5_write_en = _guard15546;
assign left_15_5_clk = clk;
assign left_15_5_reset = reset;
assign left_15_5_in = left_15_4_out;
assign pe_15_12_mul_ready =
  _guard15552 ? 1'd1 :
  _guard15555 ? 1'd0 :
  1'd0;
assign pe_15_12_clk = clk;
assign pe_15_12_top =
  _guard15568 ? top_15_12_out :
  32'd0;
assign pe_15_12_left =
  _guard15581 ? left_15_12_out :
  32'd0;
assign pe_15_12_reset = reset;
assign pe_15_12_go = _guard15594;
assign t7_add_left = 5'd1;
assign t7_add_right = t7_idx_out;
assign t13_add_left = 5'd1;
assign t13_add_right = t13_idx_out;
assign l4_idx_write_en = _guard15613;
assign l4_idx_clk = clk;
assign l4_idx_reset = reset;
assign l4_idx_in =
  _guard15616 ? 5'd0 :
  _guard15619 ? l4_add_out :
  'x;
assign l10_add_left = 5'd1;
assign l10_add_right = l10_idx_out;
assign l15_idx_write_en = _guard15632;
assign l15_idx_clk = clk;
assign l15_idx_reset = reset;
assign l15_idx_in =
  _guard15635 ? l15_add_out :
  _guard15638 ? 5'd0 :
  'x;
assign idx_write_en = _guard15643;
assign idx_clk = clk;
assign idx_reset = reset;
assign idx_in =
  _guard15644 ? idx_add_out :
  _guard15647 ? 6'd0 :
  'x;
assign idx_between_22_26_reg_write_en = _guard15652;
assign idx_between_22_26_reg_clk = clk;
assign idx_between_22_26_reg_reset = reset;
assign idx_between_22_26_reg_in =
  _guard15653 ? idx_between_22_26_comb_out :
  _guard15656 ? 1'd0 :
  'x;
assign idx_between_21_37_reg_write_en = _guard15661;
assign idx_between_21_37_reg_clk = clk;
assign idx_between_21_37_reg_reset = reset;
assign idx_between_21_37_reg_in =
  _guard15662 ? idx_between_21_37_comb_out :
  _guard15665 ? 1'd0 :
  'x;
assign index_ge_21_left = idx_add_out;
assign index_ge_21_right = 6'd21;
assign index_ge_31_left = idx_add_out;
assign index_ge_31_right = 6'd31;
assign idx_between_33_49_reg_write_en = _guard15674;
assign idx_between_33_49_reg_clk = clk;
assign idx_between_33_49_reg_reset = reset;
assign idx_between_33_49_reg_in =
  _guard15677 ? 1'd0 :
  _guard15678 ? idx_between_33_49_comb_out :
  'x;
assign idx_between_20_24_comb_left = index_ge_20_out;
assign idx_between_20_24_comb_right = index_lt_24_out;
assign idx_between_38_39_comb_left = index_ge_38_out;
assign idx_between_38_39_comb_right = index_lt_39_out;
assign idx_between_48_49_comb_left = index_ge_48_out;
assign idx_between_48_49_comb_right = index_lt_49_out;
assign idx_between_25_29_comb_left = index_ge_25_out;
assign idx_between_25_29_comb_right = index_lt_29_out;
assign idx_between_7_23_comb_left = index_ge_7_out;
assign idx_between_7_23_comb_right = index_lt_23_out;
assign index_lt_35_left = idx_add_out;
assign index_lt_35_right = 6'd35;
assign index_ge_49_left = idx_add_out;
assign index_ge_49_right = 6'd49;
assign idx_between_5_9_reg_write_en = _guard15697;
assign idx_between_5_9_reg_clk = clk;
assign idx_between_5_9_reg_reset = reset;
assign idx_between_5_9_reg_in =
  _guard15698 ? idx_between_5_9_comb_out :
  _guard15701 ? 1'd0 :
  'x;
assign index_ge_34_left = idx_add_out;
assign index_ge_34_right = 6'd34;
assign idx_between_28_29_comb_left = index_ge_28_out;
assign idx_between_28_29_comb_right = index_lt_29_out;
assign index_lt_15_left = idx_add_out;
assign index_lt_15_right = 6'd15;
assign idx_between_32_33_comb_left = index_ge_32_out;
assign idx_between_32_33_comb_right = index_lt_33_out;
assign idx_between_19_23_comb_left = index_ge_19_out;
assign idx_between_19_23_comb_right = index_lt_23_out;
assign cond7_write_en = _guard15712;
assign cond7_clk = clk;
assign cond7_reset = reset;
assign cond7_in =
  _guard15713 ? idx_between_6_22_reg_out :
  1'd0;
assign cond_wire8_in =
  _guard15714 ? idx_between_22_23_reg_out :
  _guard15717 ? cond8_out :
  1'd0;
assign cond9_write_en = _guard15718;
assign cond9_clk = clk;
assign cond9_reset = reset;
assign cond9_in =
  _guard15719 ? idx_between_2_18_reg_out :
  1'd0;
assign cond14_write_en = _guard15720;
assign cond14_clk = clk;
assign cond14_reset = reset;
assign cond14_in =
  _guard15721 ? idx_between_3_19_reg_out :
  1'd0;
assign cond_wire20_in =
  _guard15722 ? idx_between_5_9_reg_out :
  _guard15725 ? cond20_out :
  1'd0;
assign cond27_write_en = _guard15726;
assign cond27_clk = clk;
assign cond27_reset = reset;
assign cond27_in =
  _guard15727 ? idx_between_10_26_reg_out :
  1'd0;
assign cond32_write_en = _guard15728;
assign cond32_clk = clk;
assign cond32_reset = reset;
assign cond32_in =
  _guard15729 ? idx_between_11_27_reg_out :
  1'd0;
assign cond_wire37_in =
  _guard15730 ? idx_between_12_28_reg_out :
  _guard15733 ? cond37_out :
  1'd0;
assign cond50_write_en = _guard15734;
assign cond50_clk = clk;
assign cond50_reset = reset;
assign cond50_in =
  _guard15735 ? idx_between_11_15_reg_out :
  1'd0;
assign cond_wire60_in =
  _guard15738 ? cond60_out :
  _guard15739 ? idx_between_13_17_reg_out :
  1'd0;
assign cond_wire64_in =
  _guard15740 ? idx_between_13_29_reg_out :
  _guard15743 ? cond64_out :
  1'd0;
assign cond_wire81_in =
  _guard15746 ? cond81_out :
  _guard15747 ? idx_between_2_18_reg_out :
  1'd0;
assign cond_wire82_in =
  _guard15748 ? idx_between_6_22_reg_out :
  _guard15751 ? cond82_out :
  1'd0;
assign cond83_write_en = _guard15752;
assign cond83_clk = clk;
assign cond83_reset = reset;
assign cond83_in =
  _guard15753 ? idx_between_22_23_reg_out :
  1'd0;
assign cond_wire86_in =
  _guard15754 ? idx_between_7_23_reg_out :
  _guard15757 ? cond86_out :
  1'd0;
assign cond_wire87_in =
  _guard15758 ? idx_between_23_24_reg_out :
  _guard15761 ? cond87_out :
  1'd0;
assign cond91_write_en = _guard15762;
assign cond91_clk = clk;
assign cond91_reset = reset;
assign cond91_in =
  _guard15763 ? idx_between_24_25_reg_out :
  1'd0;
assign cond_wire105_in =
  _guard15766 ? cond105_out :
  _guard15767 ? idx_between_8_24_reg_out :
  1'd0;
assign cond116_write_en = _guard15768;
assign cond116_clk = clk;
assign cond116_reset = reset;
assign cond116_in =
  _guard15769 ? idx_between_11_15_reg_out :
  1'd0;
assign cond_wire117_in =
  _guard15770 ? idx_between_11_27_reg_out :
  _guard15773 ? cond117_out :
  1'd0;
assign cond_wire138_in =
  _guard15774 ? idx_between_20_36_reg_out :
  _guard15777 ? cond138_out :
  1'd0;
assign cond_wire140_in =
  _guard15778 ? idx_between_17_21_reg_out :
  _guard15781 ? cond140_out :
  1'd0;
assign cond_wire156_in =
  _guard15782 ? idx_between_25_26_reg_out :
  _guard15785 ? cond156_out :
  1'd0;
assign cond161_write_en = _guard15786;
assign cond161_clk = clk;
assign cond161_reset = reset;
assign cond161_in =
  _guard15787 ? idx_between_7_11_reg_out :
  1'd0;
assign cond174_write_en = _guard15788;
assign cond174_clk = clk;
assign cond174_reset = reset;
assign cond174_in =
  _guard15789 ? idx_between_10_26_reg_out :
  1'd0;
assign cond176_write_en = _guard15790;
assign cond176_clk = clk;
assign cond176_reset = reset;
assign cond176_in =
  _guard15791 ? idx_between_30_31_reg_out :
  1'd0;
assign cond_wire187_in =
  _guard15792 ? idx_between_17_33_reg_out :
  _guard15795 ? cond187_out :
  1'd0;
assign cond_wire190_in =
  _guard15796 ? idx_between_14_30_reg_out :
  _guard15799 ? cond190_out :
  1'd0;
assign cond194_write_en = _guard15800;
assign cond194_clk = clk;
assign cond194_reset = reset;
assign cond194_in =
  _guard15801 ? idx_between_15_31_reg_out :
  1'd0;
assign cond201_write_en = _guard15802;
assign cond201_clk = clk;
assign cond201_reset = reset;
assign cond201_in =
  _guard15803 ? idx_between_17_21_reg_out :
  1'd0;
assign cond205_write_en = _guard15804;
assign cond205_clk = clk;
assign cond205_reset = reset;
assign cond205_in =
  _guard15805 ? idx_between_18_22_reg_out :
  1'd0;
assign cond_wire207_in =
  _guard15808 ? cond207_out :
  _guard15809 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire209_in =
  _guard15810 ? idx_between_3_19_reg_out :
  _guard15813 ? cond209_out :
  1'd0;
assign cond219_write_en = _guard15814;
assign cond219_clk = clk;
assign cond219_reset = reset;
assign cond219_in =
  _guard15815 ? idx_between_6_22_reg_out :
  1'd0;
assign cond221_write_en = _guard15816;
assign cond221_clk = clk;
assign cond221_reset = reset;
assign cond221_in =
  _guard15817 ? idx_between_26_27_reg_out :
  1'd0;
assign cond225_write_en = _guard15818;
assign cond225_clk = clk;
assign cond225_reset = reset;
assign cond225_in =
  _guard15819 ? idx_between_27_28_reg_out :
  1'd0;
assign cond256_write_en = _guard15820;
assign cond256_clk = clk;
assign cond256_reset = reset;
assign cond256_in =
  _guard15821 ? idx_between_19_35_reg_out :
  1'd0;
assign cond275_write_en = _guard15822;
assign cond275_clk = clk;
assign cond275_reset = reset;
assign cond275_in =
  _guard15823 ? idx_between_5_9_reg_out :
  1'd0;
assign cond286_write_en = _guard15824;
assign cond286_clk = clk;
assign cond286_reset = reset;
assign cond286_in =
  _guard15825 ? idx_between_27_28_reg_out :
  1'd0;
assign cond_wire287_in =
  _guard15828 ? cond287_out :
  _guard15829 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire319_in =
  _guard15830 ? idx_between_16_20_reg_out :
  _guard15833 ? cond319_out :
  1'd0;
assign cond_wire345_in =
  _guard15834 ? idx_between_7_23_reg_out :
  _guard15837 ? cond345_out :
  1'd0;
assign cond363_write_en = _guard15838;
assign cond363_clk = clk;
assign cond363_reset = reset;
assign cond363_in =
  _guard15839 ? idx_between_31_32_reg_out :
  1'd0;
assign cond368_write_en = _guard15840;
assign cond368_clk = clk;
assign cond368_reset = reset;
assign cond368_in =
  _guard15841 ? idx_between_13_17_reg_out :
  1'd0;
assign cond385_write_en = _guard15842;
assign cond385_clk = clk;
assign cond385_reset = reset;
assign cond385_in =
  _guard15843 ? idx_between_17_33_reg_out :
  1'd0;
assign cond_wire409_in =
  _guard15844 ? idx_between_8_12_reg_out :
  _guard15847 ? cond409_out :
  1'd0;
assign cond419_write_en = _guard15848;
assign cond419_clk = clk;
assign cond419_reset = reset;
assign cond419_in =
  _guard15849 ? idx_between_14_30_reg_out :
  1'd0;
assign cond428_write_en = _guard15850;
assign cond428_clk = clk;
assign cond428_reset = reset;
assign cond428_in =
  _guard15851 ? idx_between_32_33_reg_out :
  1'd0;
assign cond_wire428_in =
  _guard15852 ? idx_between_32_33_reg_out :
  _guard15855 ? cond428_out :
  1'd0;
assign cond_wire433_in =
  _guard15858 ? cond433_out :
  _guard15859 ? idx_between_14_18_reg_out :
  1'd0;
assign cond442_write_en = _guard15860;
assign cond442_clk = clk;
assign cond442_reset = reset;
assign cond442_in =
  _guard15861 ? idx_between_16_32_reg_out :
  1'd0;
assign cond_wire442_in =
  _guard15862 ? idx_between_16_32_reg_out :
  _guard15865 ? cond442_out :
  1'd0;
assign cond_wire446_in =
  _guard15866 ? idx_between_17_33_reg_out :
  _guard15869 ? cond446_out :
  1'd0;
assign cond450_write_en = _guard15870;
assign cond450_clk = clk;
assign cond450_reset = reset;
assign cond450_in =
  _guard15871 ? idx_between_18_34_reg_out :
  1'd0;
assign cond481_write_en = _guard15872;
assign cond481_clk = clk;
assign cond481_reset = reset;
assign cond481_in =
  _guard15873 ? idx_between_30_31_reg_out :
  1'd0;
assign cond_wire486_in =
  _guard15876 ? cond486_out :
  _guard15877 ? idx_between_12_16_reg_out :
  1'd0;
assign cond_wire487_in =
  _guard15878 ? idx_between_12_28_reg_out :
  _guard15881 ? cond487_out :
  1'd0;
assign cond501_write_en = _guard15882;
assign cond501_clk = clk;
assign cond501_reset = reset;
assign cond501_in =
  _guard15883 ? idx_between_35_36_reg_out :
  1'd0;
assign cond_wire502_in =
  _guard15884 ? idx_between_16_20_reg_out :
  _guard15887 ? cond502_out :
  1'd0;
assign cond_wire524_in =
  _guard15890 ? cond524_out :
  _guard15891 ? idx_between_25_41_reg_out :
  1'd0;
assign cond525_write_en = _guard15892;
assign cond525_clk = clk;
assign cond525_reset = reset;
assign cond525_in =
  _guard15893 ? idx_between_41_42_reg_out :
  1'd0;
assign cond557_write_en = _guard15894;
assign cond557_clk = clk;
assign cond557_reset = reset;
assign cond557_in =
  _guard15895 ? idx_between_18_34_reg_out :
  1'd0;
assign cond567_write_en = _guard15896;
assign cond567_clk = clk;
assign cond567_reset = reset;
assign cond567_in =
  _guard15897 ? idx_between_17_21_reg_out :
  1'd0;
assign cond_wire583_in =
  _guard15898 ? idx_between_21_25_reg_out :
  _guard15901 ? cond583_out :
  1'd0;
assign cond_wire585_in =
  _guard15904 ? cond585_out :
  _guard15905 ? idx_between_25_41_reg_out :
  1'd0;
assign cond622_write_en = _guard15906;
assign cond622_clk = clk;
assign cond622_reset = reset;
assign cond622_in =
  _guard15907 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire628_in =
  _guard15910 ? cond628_out :
  _guard15911 ? idx_between_17_21_reg_out :
  1'd0;
assign cond651_write_en = _guard15912;
assign cond651_clk = clk;
assign cond651_reset = reset;
assign cond651_in =
  _guard15913 ? idx_between_42_43_reg_out :
  1'd0;
assign cond657_write_en = _guard15914;
assign cond657_clk = clk;
assign cond657_reset = reset;
assign cond657_in =
  _guard15915 ? idx_between_24_40_reg_out :
  1'd0;
assign cond664_write_en = _guard15916;
assign cond664_clk = clk;
assign cond664_reset = reset;
assign cond664_in =
  _guard15917 ? idx_between_10_26_reg_out :
  1'd0;
assign cond669_write_en = _guard15918;
assign cond669_clk = clk;
assign cond669_reset = reset;
assign cond669_in =
  _guard15919 ? idx_between_12_16_reg_out :
  1'd0;
assign cond_wire687_in =
  _guard15920 ? idx_between_20_36_reg_out :
  _guard15923 ? cond687_out :
  1'd0;
assign cond699_write_en = _guard15924;
assign cond699_clk = clk;
assign cond699_reset = reset;
assign cond699_in =
  _guard15925 ? idx_between_23_39_reg_out :
  1'd0;
assign cond706_write_en = _guard15926;
assign cond706_clk = clk;
assign cond706_reset = reset;
assign cond706_in =
  _guard15927 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire729_in =
  _guard15928 ? idx_between_11_27_reg_out :
  _guard15931 ? cond729_out :
  1'd0;
assign cond_wire750_in =
  _guard15932 ? idx_between_17_21_reg_out :
  _guard15935 ? cond750_out :
  1'd0;
assign cond783_write_en = _guard15936;
assign cond783_clk = clk;
assign cond783_reset = reset;
assign cond783_in =
  _guard15937 ? idx_between_25_41_reg_out :
  1'd0;
assign cond_wire783_in =
  _guard15940 ? cond783_out :
  _guard15941 ? idx_between_25_41_reg_out :
  1'd0;
assign cond788_write_en = _guard15942;
assign cond788_clk = clk;
assign cond788_reset = reset;
assign cond788_in =
  _guard15943 ? idx_between_30_46_reg_out :
  1'd0;
assign cond793_write_en = _guard15944;
assign cond793_clk = clk;
assign cond793_reset = reset;
assign cond793_in =
  _guard15945 ? idx_between_47_48_reg_out :
  1'd0;
assign cond798_write_en = _guard15946;
assign cond798_clk = clk;
assign cond798_reset = reset;
assign cond798_in =
  _guard15947 ? idx_between_33_34_reg_out :
  1'd0;
assign cond_wire810_in =
  _guard15948 ? idx_between_36_37_reg_out :
  _guard15951 ? cond810_out :
  1'd0;
assign cond_wire811_in =
  _guard15954 ? cond811_out :
  _guard15955 ? idx_between_17_21_reg_out :
  1'd0;
assign cond817_write_en = _guard15956;
assign cond817_clk = clk;
assign cond817_reset = reset;
assign cond817_in =
  _guard15957 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire830_in =
  _guard15960 ? cond830_out :
  _guard15961 ? idx_between_41_42_reg_out :
  1'd0;
assign cond_wire840_in =
  _guard15964 ? cond840_out :
  _guard15965 ? idx_between_24_40_reg_out :
  1'd0;
assign cond_wire866_in =
  _guard15968 ? cond866_out :
  _guard15969 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire869_in =
  _guard15970 ? idx_between_16_32_reg_out :
  _guard15973 ? cond869_out :
  1'd0;
assign cond_wire876_in =
  _guard15976 ? cond876_out :
  _guard15977 ? idx_between_18_22_reg_out :
  1'd0;
assign cond_wire884_in =
  _guard15980 ? cond884_out :
  _guard15981 ? idx_between_20_24_reg_out :
  1'd0;
assign cond885_write_en = _guard15982;
assign cond885_clk = clk;
assign cond885_reset = reset;
assign cond885_in =
  _guard15983 ? idx_between_20_36_reg_out :
  1'd0;
assign cond896_write_en = _guard15984;
assign cond896_clk = clk;
assign cond896_reset = reset;
assign cond896_in =
  _guard15985 ? idx_between_23_27_reg_out :
  1'd0;
assign cond904_write_en = _guard15986;
assign cond904_clk = clk;
assign cond904_reset = reset;
assign cond904_in =
  _guard15987 ? idx_between_25_29_reg_out :
  1'd0;
assign cond_wire924_in =
  _guard15990 ? cond924_out :
  _guard15991 ? idx_between_14_30_reg_out :
  1'd0;
assign cond934_write_en = _guard15992;
assign cond934_clk = clk;
assign cond934_reset = reset;
assign cond934_in =
  _guard15993 ? idx_between_17_33_reg_out :
  1'd0;
assign cond938_write_en = _guard15994;
assign cond938_clk = clk;
assign cond938_reset = reset;
assign cond938_in =
  _guard15995 ? idx_between_18_34_reg_out :
  1'd0;
assign cond942_write_en = _guard15996;
assign cond942_clk = clk;
assign cond942_reset = reset;
assign cond942_in =
  _guard15997 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire945_in =
  _guard16000 ? cond945_out :
  _guard16001 ? idx_between_20_24_reg_out :
  1'd0;
assign cond_wire959_in =
  _guard16002 ? idx_between_27_43_reg_out :
  _guard16005 ? cond959_out :
  1'd0;
assign cond971_write_en = _guard16006;
assign cond971_clk = clk;
assign cond971_reset = reset;
assign cond971_in =
  _guard16007 ? idx_between_30_46_reg_out :
  1'd0;
assign cond_wire993_in =
  _guard16010 ? cond993_out :
  _guard16011 ? idx_between_36_37_reg_out :
  1'd0;
assign cond1011_write_en = _guard16012;
assign cond1011_clk = clk;
assign cond1011_reset = reset;
assign cond1011_in =
  _guard16013 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire1016_in =
  _guard16016 ? cond1016_out :
  _guard16017 ? idx_between_26_42_reg_out :
  1'd0;
assign cond_wire1019_in =
  _guard16018 ? idx_between_23_39_reg_out :
  _guard16021 ? cond1019_out :
  1'd0;
assign cond_wire1033_in =
  _guard16024 ? cond1033_out :
  _guard16025 ? idx_between_46_47_reg_out :
  1'd0;
assign cond_wire1034_in =
  _guard16028 ? cond1034_out :
  _guard16029 ? idx_between_27_31_reg_out :
  1'd0;
assign wrapper_early_reset_static_seq_done_in = _guard16032;
assign top_0_1_write_en = _guard16035;
assign top_0_1_clk = clk;
assign top_0_1_reset = reset;
assign top_0_1_in = t1_read_data;
assign left_0_2_write_en = _guard16041;
assign left_0_2_clk = clk;
assign left_0_2_reset = reset;
assign left_0_2_in = left_0_1_out;
assign pe_0_4_mul_ready =
  _guard16047 ? 1'd1 :
  _guard16050 ? 1'd0 :
  1'd0;
assign pe_0_4_clk = clk;
assign pe_0_4_top =
  _guard16063 ? top_0_4_out :
  32'd0;
assign pe_0_4_left =
  _guard16076 ? left_0_4_out :
  32'd0;
assign pe_0_4_reset = reset;
assign pe_0_4_go = _guard16089;
assign top_0_9_write_en = _guard16092;
assign top_0_9_clk = clk;
assign top_0_9_reset = reset;
assign top_0_9_in = t9_read_data;
assign left_0_10_write_en = _guard16098;
assign left_0_10_clk = clk;
assign left_0_10_reset = reset;
assign left_0_10_in = left_0_9_out;
assign pe_0_14_mul_ready =
  _guard16104 ? 1'd1 :
  _guard16107 ? 1'd0 :
  1'd0;
assign pe_0_14_clk = clk;
assign pe_0_14_top =
  _guard16120 ? top_0_14_out :
  32'd0;
assign pe_0_14_left =
  _guard16133 ? left_0_14_out :
  32'd0;
assign pe_0_14_reset = reset;
assign pe_0_14_go = _guard16146;
assign pe_1_9_mul_ready =
  _guard16149 ? 1'd1 :
  _guard16152 ? 1'd0 :
  1'd0;
assign pe_1_9_clk = clk;
assign pe_1_9_top =
  _guard16165 ? top_1_9_out :
  32'd0;
assign pe_1_9_left =
  _guard16178 ? left_1_9_out :
  32'd0;
assign pe_1_9_reset = reset;
assign pe_1_9_go = _guard16191;
assign top_2_3_write_en = _guard16194;
assign top_2_3_clk = clk;
assign top_2_3_reset = reset;
assign top_2_3_in = top_1_3_out;
assign pe_2_6_mul_ready =
  _guard16200 ? 1'd1 :
  _guard16203 ? 1'd0 :
  1'd0;
assign pe_2_6_clk = clk;
assign pe_2_6_top =
  _guard16216 ? top_2_6_out :
  32'd0;
assign pe_2_6_left =
  _guard16229 ? left_2_6_out :
  32'd0;
assign pe_2_6_reset = reset;
assign pe_2_6_go = _guard16242;
assign pe_2_8_mul_ready =
  _guard16245 ? 1'd1 :
  _guard16248 ? 1'd0 :
  1'd0;
assign pe_2_8_clk = clk;
assign pe_2_8_top =
  _guard16261 ? top_2_8_out :
  32'd0;
assign pe_2_8_left =
  _guard16274 ? left_2_8_out :
  32'd0;
assign pe_2_8_reset = reset;
assign pe_2_8_go = _guard16287;
assign top_2_13_write_en = _guard16290;
assign top_2_13_clk = clk;
assign top_2_13_reset = reset;
assign top_2_13_in = top_1_13_out;
assign left_3_0_write_en = _guard16296;
assign left_3_0_clk = clk;
assign left_3_0_reset = reset;
assign left_3_0_in = l3_read_data;
assign pe_3_9_mul_ready =
  _guard16302 ? 1'd1 :
  _guard16305 ? 1'd0 :
  1'd0;
assign pe_3_9_clk = clk;
assign pe_3_9_top =
  _guard16318 ? top_3_9_out :
  32'd0;
assign pe_3_9_left =
  _guard16331 ? left_3_9_out :
  32'd0;
assign pe_3_9_reset = reset;
assign pe_3_9_go = _guard16344;
assign pe_3_11_mul_ready =
  _guard16347 ? 1'd1 :
  _guard16350 ? 1'd0 :
  1'd0;
assign pe_3_11_clk = clk;
assign pe_3_11_top =
  _guard16363 ? top_3_11_out :
  32'd0;
assign pe_3_11_left =
  _guard16376 ? left_3_11_out :
  32'd0;
assign pe_3_11_reset = reset;
assign pe_3_11_go = _guard16389;
assign pe_4_2_mul_ready =
  _guard16392 ? 1'd1 :
  _guard16395 ? 1'd0 :
  1'd0;
assign pe_4_2_clk = clk;
assign pe_4_2_top =
  _guard16408 ? top_4_2_out :
  32'd0;
assign pe_4_2_left =
  _guard16421 ? left_4_2_out :
  32'd0;
assign pe_4_2_reset = reset;
assign pe_4_2_go = _guard16434;
assign pe_4_8_mul_ready =
  _guard16437 ? 1'd1 :
  _guard16440 ? 1'd0 :
  1'd0;
assign pe_4_8_clk = clk;
assign pe_4_8_top =
  _guard16453 ? top_4_8_out :
  32'd0;
assign pe_4_8_left =
  _guard16466 ? left_4_8_out :
  32'd0;
assign pe_4_8_reset = reset;
assign pe_4_8_go = _guard16479;
assign top_5_1_write_en = _guard16482;
assign top_5_1_clk = clk;
assign top_5_1_reset = reset;
assign top_5_1_in = top_4_1_out;
assign left_5_4_write_en = _guard16488;
assign left_5_4_clk = clk;
assign left_5_4_reset = reset;
assign left_5_4_in = left_5_3_out;
assign left_5_14_write_en = _guard16494;
assign left_5_14_clk = clk;
assign left_5_14_reset = reset;
assign left_5_14_in = left_5_13_out;
assign pe_6_7_mul_ready =
  _guard16500 ? 1'd1 :
  _guard16503 ? 1'd0 :
  1'd0;
assign pe_6_7_clk = clk;
assign pe_6_7_top =
  _guard16516 ? top_6_7_out :
  32'd0;
assign pe_6_7_left =
  _guard16529 ? left_6_7_out :
  32'd0;
assign pe_6_7_reset = reset;
assign pe_6_7_go = _guard16542;
assign top_6_11_write_en = _guard16545;
assign top_6_11_clk = clk;
assign top_6_11_reset = reset;
assign top_6_11_in = top_5_11_out;
assign pe_6_13_mul_ready =
  _guard16551 ? 1'd1 :
  _guard16554 ? 1'd0 :
  1'd0;
assign pe_6_13_clk = clk;
assign pe_6_13_top =
  _guard16567 ? top_6_13_out :
  32'd0;
assign pe_6_13_left =
  _guard16580 ? left_6_13_out :
  32'd0;
assign pe_6_13_reset = reset;
assign pe_6_13_go = _guard16593;
assign pe_6_14_mul_ready =
  _guard16596 ? 1'd1 :
  _guard16599 ? 1'd0 :
  1'd0;
assign pe_6_14_clk = clk;
assign pe_6_14_top =
  _guard16612 ? top_6_14_out :
  32'd0;
assign pe_6_14_left =
  _guard16625 ? left_6_14_out :
  32'd0;
assign pe_6_14_reset = reset;
assign pe_6_14_go = _guard16638;
assign pe_6_15_mul_ready =
  _guard16641 ? 1'd1 :
  _guard16644 ? 1'd0 :
  1'd0;
assign pe_6_15_clk = clk;
assign pe_6_15_top =
  _guard16657 ? top_6_15_out :
  32'd0;
assign pe_6_15_left =
  _guard16670 ? left_6_15_out :
  32'd0;
assign pe_6_15_reset = reset;
assign pe_6_15_go = _guard16683;
assign left_8_3_write_en = _guard16686;
assign left_8_3_clk = clk;
assign left_8_3_reset = reset;
assign left_8_3_in = left_8_2_out;
assign pe_9_0_mul_ready =
  _guard16692 ? 1'd1 :
  _guard16695 ? 1'd0 :
  1'd0;
assign pe_9_0_clk = clk;
assign pe_9_0_top =
  _guard16708 ? top_9_0_out :
  32'd0;
assign pe_9_0_left =
  _guard16721 ? left_9_0_out :
  32'd0;
assign pe_9_0_reset = reset;
assign pe_9_0_go = _guard16734;
assign left_9_1_write_en = _guard16737;
assign left_9_1_clk = clk;
assign left_9_1_reset = reset;
assign left_9_1_in = left_9_0_out;
assign left_9_2_write_en = _guard16743;
assign left_9_2_clk = clk;
assign left_9_2_reset = reset;
assign left_9_2_in = left_9_1_out;
assign pe_9_4_mul_ready =
  _guard16749 ? 1'd1 :
  _guard16752 ? 1'd0 :
  1'd0;
assign pe_9_4_clk = clk;
assign pe_9_4_top =
  _guard16765 ? top_9_4_out :
  32'd0;
assign pe_9_4_left =
  _guard16778 ? left_9_4_out :
  32'd0;
assign pe_9_4_reset = reset;
assign pe_9_4_go = _guard16791;
assign left_9_14_write_en = _guard16794;
assign left_9_14_clk = clk;
assign left_9_14_reset = reset;
assign left_9_14_in = left_9_13_out;
assign left_9_15_write_en = _guard16800;
assign left_9_15_clk = clk;
assign left_9_15_reset = reset;
assign left_9_15_in = left_9_14_out;
assign pe_10_10_mul_ready =
  _guard16806 ? 1'd1 :
  _guard16809 ? 1'd0 :
  1'd0;
assign pe_10_10_clk = clk;
assign pe_10_10_top =
  _guard16822 ? top_10_10_out :
  32'd0;
assign pe_10_10_left =
  _guard16835 ? left_10_10_out :
  32'd0;
assign pe_10_10_reset = reset;
assign pe_10_10_go = _guard16848;
assign top_10_10_write_en = _guard16851;
assign top_10_10_clk = clk;
assign top_10_10_reset = reset;
assign top_10_10_in = top_9_10_out;
assign pe_12_1_mul_ready =
  _guard16857 ? 1'd1 :
  _guard16860 ? 1'd0 :
  1'd0;
assign pe_12_1_clk = clk;
assign pe_12_1_top =
  _guard16873 ? top_12_1_out :
  32'd0;
assign pe_12_1_left =
  _guard16886 ? left_12_1_out :
  32'd0;
assign pe_12_1_reset = reset;
assign pe_12_1_go = _guard16899;
assign left_12_1_write_en = _guard16902;
assign left_12_1_clk = clk;
assign left_12_1_reset = reset;
assign left_12_1_in = left_12_0_out;
assign top_12_5_write_en = _guard16908;
assign top_12_5_clk = clk;
assign top_12_5_reset = reset;
assign top_12_5_in = top_11_5_out;
assign pe_12_7_mul_ready =
  _guard16914 ? 1'd1 :
  _guard16917 ? 1'd0 :
  1'd0;
assign pe_12_7_clk = clk;
assign pe_12_7_top =
  _guard16930 ? top_12_7_out :
  32'd0;
assign pe_12_7_left =
  _guard16943 ? left_12_7_out :
  32'd0;
assign pe_12_7_reset = reset;
assign pe_12_7_go = _guard16956;
assign pe_12_11_mul_ready =
  _guard16959 ? 1'd1 :
  _guard16962 ? 1'd0 :
  1'd0;
assign pe_12_11_clk = clk;
assign pe_12_11_top =
  _guard16975 ? top_12_11_out :
  32'd0;
assign pe_12_11_left =
  _guard16988 ? left_12_11_out :
  32'd0;
assign pe_12_11_reset = reset;
assign pe_12_11_go = _guard17001;
assign top_13_3_write_en = _guard17004;
assign top_13_3_clk = clk;
assign top_13_3_reset = reset;
assign top_13_3_in = top_12_3_out;
assign top_13_8_write_en = _guard17010;
assign top_13_8_clk = clk;
assign top_13_8_reset = reset;
assign top_13_8_in = top_12_8_out;
assign pe_13_11_mul_ready =
  _guard17016 ? 1'd1 :
  _guard17019 ? 1'd0 :
  1'd0;
assign pe_13_11_clk = clk;
assign pe_13_11_top =
  _guard17032 ? top_13_11_out :
  32'd0;
assign pe_13_11_left =
  _guard17045 ? left_13_11_out :
  32'd0;
assign pe_13_11_reset = reset;
assign pe_13_11_go = _guard17058;
assign left_13_14_write_en = _guard17061;
assign left_13_14_clk = clk;
assign left_13_14_reset = reset;
assign left_13_14_in = left_13_13_out;
assign top_14_7_write_en = _guard17067;
assign top_14_7_clk = clk;
assign top_14_7_reset = reset;
assign top_14_7_in = top_13_7_out;
assign left_14_12_write_en = _guard17073;
assign left_14_12_clk = clk;
assign left_14_12_reset = reset;
assign left_14_12_in = left_14_11_out;
assign left_14_13_write_en = _guard17079;
assign left_14_13_clk = clk;
assign left_14_13_reset = reset;
assign left_14_13_in = left_14_12_out;
assign left_15_0_write_en = _guard17085;
assign left_15_0_clk = clk;
assign left_15_0_reset = reset;
assign left_15_0_in = l15_read_data;
assign top_15_6_write_en = _guard17091;
assign top_15_6_clk = clk;
assign top_15_6_reset = reset;
assign top_15_6_in = top_14_6_out;
assign top_15_10_write_en = _guard17097;
assign top_15_10_clk = clk;
assign top_15_10_reset = reset;
assign top_15_10_in = top_14_10_out;
assign pe_15_11_mul_ready =
  _guard17103 ? 1'd1 :
  _guard17106 ? 1'd0 :
  1'd0;
assign pe_15_11_clk = clk;
assign pe_15_11_top =
  _guard17119 ? top_15_11_out :
  32'd0;
assign pe_15_11_left =
  _guard17132 ? left_15_11_out :
  32'd0;
assign pe_15_11_reset = reset;
assign pe_15_11_go = _guard17145;
assign t14_add_left = 5'd1;
assign t14_add_right = t14_idx_out;
assign l7_add_left = 5'd1;
assign l7_add_right = l7_idx_out;
assign l12_add_left = 5'd1;
assign l12_add_right = l12_idx_out;
assign idx_between_30_46_comb_left = index_ge_30_out;
assign idx_between_30_46_comb_right = index_lt_46_out;
assign index_lt_47_left = idx_add_out;
assign index_lt_47_right = 6'd47;
assign index_ge_1_left = idx_add_out;
assign index_ge_1_right = 6'd1;
assign idx_between_50_51_reg_write_en = _guard17174;
assign idx_between_50_51_reg_clk = clk;
assign idx_between_50_51_reg_reset = reset;
assign idx_between_50_51_reg_in =
  _guard17175 ? idx_between_50_51_comb_out :
  _guard17178 ? 1'd0 :
  'x;
assign idx_between_51_52_reg_write_en = _guard17183;
assign idx_between_51_52_reg_clk = clk;
assign idx_between_51_52_reg_reset = reset;
assign idx_between_51_52_reg_in =
  _guard17184 ? idx_between_51_52_comb_out :
  _guard17187 ? 1'd0 :
  'x;
assign idx_between_51_52_comb_left = index_ge_51_out;
assign idx_between_51_52_comb_right = index_lt_52_out;
assign index_ge_32_left = idx_add_out;
assign index_ge_32_right = 6'd32;
assign index_lt_9_left = idx_add_out;
assign index_lt_9_right = 6'd9;
assign index_ge_4_left = idx_add_out;
assign index_ge_4_right = 6'd4;
assign idx_between_1_5_reg_write_en = _guard17200;
assign idx_between_1_5_reg_clk = clk;
assign idx_between_1_5_reg_reset = reset;
assign idx_between_1_5_reg_in =
  _guard17203 ? 1'd0 :
  _guard17204 ? idx_between_1_5_comb_out :
  'x;
assign idx_between_24_25_reg_write_en = _guard17209;
assign idx_between_24_25_reg_clk = clk;
assign idx_between_24_25_reg_reset = reset;
assign idx_between_24_25_reg_in =
  _guard17210 ? idx_between_24_25_comb_out :
  _guard17213 ? 1'd0 :
  'x;
assign index_lt_6_left = idx_add_out;
assign index_lt_6_right = 6'd6;
assign idx_between_3_7_comb_left = index_ge_3_out;
assign idx_between_3_7_comb_right = index_lt_7_out;
assign index_lt_8_left = idx_add_out;
assign index_lt_8_right = 6'd8;
assign idx_between_29_30_reg_write_en = _guard17224;
assign idx_between_29_30_reg_clk = clk;
assign idx_between_29_30_reg_reset = reset;
assign idx_between_29_30_reg_in =
  _guard17227 ? 1'd0 :
  _guard17228 ? idx_between_29_30_comb_out :
  'x;
assign index_lt_36_left = idx_add_out;
assign index_lt_36_right = 6'd36;
assign index_lt_44_left = idx_add_out;
assign index_lt_44_right = 6'd44;
assign cond4_write_en = _guard17233;
assign cond4_clk = clk;
assign cond4_reset = reset;
assign cond4_in =
  _guard17234 ? idx_between_1_17_reg_out :
  1'd0;
assign cond5_write_en = _guard17235;
assign cond5_clk = clk;
assign cond5_reset = reset;
assign cond5_in =
  _guard17236 ? idx_between_2_6_reg_out :
  1'd0;
assign cond_wire6_in =
  _guard17239 ? cond6_out :
  _guard17240 ? idx_between_2_18_reg_out :
  1'd0;
assign cond20_write_en = _guard17241;
assign cond20_clk = clk;
assign cond20_reset = reset;
assign cond20_in =
  _guard17242 ? idx_between_5_9_reg_out :
  1'd0;
assign cond_wire36_in =
  _guard17245 ? cond36_out :
  _guard17246 ? idx_between_8_24_reg_out :
  1'd0;
assign cond46_write_en = _guard17247;
assign cond46_clk = clk;
assign cond46_reset = reset;
assign cond46_in =
  _guard17248 ? idx_between_10_26_reg_out :
  1'd0;
assign cond_wire62_in =
  _guard17249 ? idx_between_17_33_reg_out :
  _guard17252 ? cond62_out :
  1'd0;
assign cond63_write_en = _guard17253;
assign cond63_clk = clk;
assign cond63_reset = reset;
assign cond63_in =
  _guard17254 ? idx_between_33_34_reg_out :
  1'd0;
assign cond_wire66_in =
  _guard17255 ? idx_between_14_30_reg_out :
  _guard17258 ? cond66_out :
  1'd0;
assign cond_wire74_in =
  _guard17261 ? cond74_out :
  _guard17262 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire75_in =
  _guard17263 ? idx_between_16_20_reg_out :
  _guard17266 ? cond75_out :
  1'd0;
assign cond78_write_en = _guard17267;
assign cond78_clk = clk;
assign cond78_reset = reset;
assign cond78_in =
  _guard17268 ? idx_between_36_37_reg_out :
  1'd0;
assign cond90_write_en = _guard17269;
assign cond90_clk = clk;
assign cond90_reset = reset;
assign cond90_in =
  _guard17270 ? idx_between_8_24_reg_out :
  1'd0;
assign cond_wire92_in =
  _guard17273 ? cond92_out :
  _guard17274 ? idx_between_5_9_reg_out :
  1'd0;
assign cond101_write_en = _guard17275;
assign cond101_clk = clk;
assign cond101_reset = reset;
assign cond101_in =
  _guard17276 ? idx_between_7_23_reg_out :
  1'd0;
assign cond106_write_en = _guard17277;
assign cond106_clk = clk;
assign cond106_reset = reset;
assign cond106_in =
  _guard17278 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire108_in =
  _guard17281 ? cond108_out :
  _guard17282 ? idx_between_9_13_reg_out :
  1'd0;
assign cond112_write_en = _guard17283;
assign cond112_clk = clk;
assign cond112_reset = reset;
assign cond112_in =
  _guard17284 ? idx_between_10_14_reg_out :
  1'd0;
assign cond122_write_en = _guard17285;
assign cond122_clk = clk;
assign cond122_reset = reset;
assign cond122_in =
  _guard17286 ? idx_between_16_32_reg_out :
  1'd0;
assign cond_wire122_in =
  _guard17287 ? idx_between_16_32_reg_out :
  _guard17290 ? cond122_out :
  1'd0;
assign cond_wire128_in =
  _guard17293 ? cond128_out :
  _guard17294 ? idx_between_14_18_reg_out :
  1'd0;
assign cond_wire139_in =
  _guard17295 ? idx_between_36_37_reg_out :
  _guard17298 ? cond139_out :
  1'd0;
assign cond143_write_en = _guard17299;
assign cond143_clk = clk;
assign cond143_reset = reset;
assign cond143_in =
  _guard17300 ? idx_between_37_38_reg_out :
  1'd0;
assign cond_wire143_in =
  _guard17303 ? cond143_out :
  _guard17304 ? idx_between_37_38_reg_out :
  1'd0;
assign cond148_write_en = _guard17305;
assign cond148_clk = clk;
assign cond148_reset = reset;
assign cond148_in =
  _guard17306 ? idx_between_23_24_reg_out :
  1'd0;
assign cond152_write_en = _guard17307;
assign cond152_clk = clk;
assign cond152_reset = reset;
assign cond152_in =
  _guard17308 ? idx_between_24_25_reg_out :
  1'd0;
assign cond_wire172_in =
  _guard17311 ? cond172_out :
  _guard17312 ? idx_between_29_30_reg_out :
  1'd0;
assign cond_wire178_in =
  _guard17313 ? idx_between_11_27_reg_out :
  _guard17316 ? cond178_out :
  1'd0;
assign cond_wire181_in =
  _guard17319 ? cond181_out :
  _guard17320 ? idx_between_12_16_reg_out :
  1'd0;
assign cond_wire189_in =
  _guard17323 ? cond189_out :
  _guard17324 ? idx_between_14_18_reg_out :
  1'd0;
assign cond192_write_en = _guard17325;
assign cond192_clk = clk;
assign cond192_reset = reset;
assign cond192_in =
  _guard17326 ? idx_between_34_35_reg_out :
  1'd0;
assign cond196_write_en = _guard17327;
assign cond196_clk = clk;
assign cond196_reset = reset;
assign cond196_in =
  _guard17328 ? idx_between_35_36_reg_out :
  1'd0;
assign cond203_write_en = _guard17329;
assign cond203_clk = clk;
assign cond203_reset = reset;
assign cond203_in =
  _guard17330 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire203_in =
  _guard17331 ? idx_between_21_37_reg_out :
  _guard17334 ? cond203_out :
  1'd0;
assign cond208_write_en = _guard17335;
assign cond208_clk = clk;
assign cond208_reset = reset;
assign cond208_in =
  _guard17336 ? idx_between_38_39_reg_out :
  1'd0;
assign cond_wire210_in =
  _guard17337 ? idx_between_4_8_reg_out :
  _guard17340 ? cond210_out :
  1'd0;
assign cond_wire214_in =
  _guard17343 ? cond214_out :
  _guard17344 ? idx_between_5_9_reg_out :
  1'd0;
assign cond_wire233_in =
  _guard17347 ? cond233_out :
  _guard17348 ? idx_between_29_30_reg_out :
  1'd0;
assign cond235_write_en = _guard17349;
assign cond235_clk = clk;
assign cond235_reset = reset;
assign cond235_in =
  _guard17350 ? idx_between_10_26_reg_out :
  1'd0;
assign cond_wire248_in =
  _guard17351 ? idx_between_17_33_reg_out :
  _guard17354 ? cond248_out :
  1'd0;
assign cond250_write_en = _guard17355;
assign cond250_clk = clk;
assign cond250_reset = reset;
assign cond250_in =
  _guard17356 ? idx_between_14_18_reg_out :
  1'd0;
assign cond252_write_en = _guard17357;
assign cond252_clk = clk;
assign cond252_reset = reset;
assign cond252_in =
  _guard17358 ? idx_between_18_34_reg_out :
  1'd0;
assign cond_wire253_in =
  _guard17359 ? idx_between_34_35_reg_out :
  _guard17362 ? cond253_out :
  1'd0;
assign cond_wire256_in =
  _guard17365 ? cond256_out :
  _guard17366 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire258_in =
  _guard17367 ? idx_between_16_20_reg_out :
  _guard17370 ? cond258_out :
  1'd0;
assign cond_wire268_in =
  _guard17373 ? cond268_out :
  _guard17374 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire276_in =
  _guard17377 ? cond276_out :
  _guard17378 ? idx_between_5_21_reg_out :
  1'd0;
assign cond_wire281_in =
  _guard17381 ? cond281_out :
  _guard17382 ? idx_between_10_26_reg_out :
  1'd0;
assign cond_wire282_in =
  _guard17383 ? idx_between_26_27_reg_out :
  _guard17386 ? cond282_out :
  1'd0;
assign cond283_write_en = _guard17387;
assign cond283_clk = clk;
assign cond283_reset = reset;
assign cond283_in =
  _guard17388 ? idx_between_7_11_reg_out :
  1'd0;
assign cond_wire286_in =
  _guard17389 ? idx_between_27_28_reg_out :
  _guard17392 ? cond286_out :
  1'd0;
assign cond307_write_en = _guard17393;
assign cond307_clk = clk;
assign cond307_reset = reset;
assign cond307_in =
  _guard17394 ? idx_between_13_17_reg_out :
  1'd0;
assign cond_wire311_in =
  _guard17395 ? idx_between_14_18_reg_out :
  _guard17398 ? cond311_out :
  1'd0;
assign cond314_write_en = _guard17399;
assign cond314_clk = clk;
assign cond314_reset = reset;
assign cond314_in =
  _guard17400 ? idx_between_34_35_reg_out :
  1'd0;
assign cond_wire314_in =
  _guard17401 ? idx_between_34_35_reg_out :
  _guard17404 ? cond314_out :
  1'd0;
assign cond_wire326_in =
  _guard17407 ? cond326_out :
  _guard17408 ? idx_between_37_38_reg_out :
  1'd0;
assign cond_wire337_in =
  _guard17409 ? idx_between_24_40_reg_out :
  _guard17412 ? cond337_out :
  1'd0;
assign cond_wire349_in =
  _guard17415 ? cond349_out :
  _guard17416 ? idx_between_8_24_reg_out :
  1'd0;
assign cond_wire357_in =
  _guard17419 ? cond357_out :
  _guard17420 ? idx_between_10_26_reg_out :
  1'd0;
assign cond_wire377_in =
  _guard17423 ? cond377_out :
  _guard17424 ? idx_between_15_31_reg_out :
  1'd0;
assign cond378_write_en = _guard17425;
assign cond378_clk = clk;
assign cond378_reset = reset;
assign cond378_in =
  _guard17426 ? idx_between_19_35_reg_out :
  1'd0;
assign cond380_write_en = _guard17427;
assign cond380_clk = clk;
assign cond380_reset = reset;
assign cond380_in =
  _guard17428 ? idx_between_16_20_reg_out :
  1'd0;
assign cond_wire398_in =
  _guard17431 ? cond398_out :
  _guard17432 ? idx_between_24_40_reg_out :
  1'd0;
assign cond411_write_en = _guard17433;
assign cond411_clk = clk;
assign cond411_reset = reset;
assign cond411_in =
  _guard17434 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire418_in =
  _guard17435 ? idx_between_10_26_reg_out :
  _guard17438 ? cond418_out :
  1'd0;
assign cond434_write_en = _guard17439;
assign cond434_clk = clk;
assign cond434_reset = reset;
assign cond434_in =
  _guard17440 ? idx_between_14_30_reg_out :
  1'd0;
assign cond436_write_en = _guard17441;
assign cond436_clk = clk;
assign cond436_reset = reset;
assign cond436_in =
  _guard17442 ? idx_between_34_35_reg_out :
  1'd0;
assign cond_wire436_in =
  _guard17443 ? idx_between_34_35_reg_out :
  _guard17446 ? cond436_out :
  1'd0;
assign cond452_write_en = _guard17447;
assign cond452_clk = clk;
assign cond452_reset = reset;
assign cond452_in =
  _guard17448 ? idx_between_38_39_reg_out :
  1'd0;
assign cond459_write_en = _guard17449;
assign cond459_clk = clk;
assign cond459_reset = reset;
assign cond459_in =
  _guard17450 ? idx_between_24_40_reg_out :
  1'd0;
assign cond461_write_en = _guard17451;
assign cond461_clk = clk;
assign cond461_reset = reset;
assign cond461_in =
  _guard17452 ? idx_between_21_25_reg_out :
  1'd0;
assign cond467_write_en = _guard17453;
assign cond467_clk = clk;
assign cond467_reset = reset;
assign cond467_in =
  _guard17454 ? idx_between_26_42_reg_out :
  1'd0;
assign cond472_write_en = _guard17455;
assign cond472_clk = clk;
assign cond472_reset = reset;
assign cond472_in =
  _guard17456 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire474_in =
  _guard17459 ? cond474_out :
  _guard17460 ? idx_between_9_13_reg_out :
  1'd0;
assign cond482_write_en = _guard17461;
assign cond482_clk = clk;
assign cond482_reset = reset;
assign cond482_in =
  _guard17462 ? idx_between_11_15_reg_out :
  1'd0;
assign cond486_write_en = _guard17463;
assign cond486_clk = clk;
assign cond486_reset = reset;
assign cond486_in =
  _guard17464 ? idx_between_12_16_reg_out :
  1'd0;
assign cond_wire506_in =
  _guard17467 ? cond506_out :
  _guard17468 ? idx_between_17_21_reg_out :
  1'd0;
assign cond507_write_en = _guard17469;
assign cond507_clk = clk;
assign cond507_reset = reset;
assign cond507_in =
  _guard17470 ? idx_between_17_33_reg_out :
  1'd0;
assign cond524_write_en = _guard17471;
assign cond524_clk = clk;
assign cond524_reset = reset;
assign cond524_in =
  _guard17472 ? idx_between_25_41_reg_out :
  1'd0;
assign cond526_write_en = _guard17473;
assign cond526_clk = clk;
assign cond526_reset = reset;
assign cond526_in =
  _guard17474 ? idx_between_22_26_reg_out :
  1'd0;
assign cond_wire526_in =
  _guard17475 ? idx_between_22_26_reg_out :
  _guard17478 ? cond526_out :
  1'd0;
assign cond_wire527_in =
  _guard17481 ? cond527_out :
  _guard17482 ? idx_between_22_38_reg_out :
  1'd0;
assign cond529_write_en = _guard17483;
assign cond529_clk = clk;
assign cond529_reset = reset;
assign cond529_in =
  _guard17484 ? idx_between_42_43_reg_out :
  1'd0;
assign cond_wire532_in =
  _guard17487 ? cond532_out :
  _guard17488 ? idx_between_27_43_reg_out :
  1'd0;
assign cond541_write_en = _guard17489;
assign cond541_clk = clk;
assign cond541_reset = reset;
assign cond541_in =
  _guard17490 ? idx_between_14_30_reg_out :
  1'd0;
assign cond543_write_en = _guard17491;
assign cond543_clk = clk;
assign cond543_reset = reset;
assign cond543_in =
  _guard17492 ? idx_between_11_15_reg_out :
  1'd0;
assign cond545_write_en = _guard17493;
assign cond545_clk = clk;
assign cond545_reset = reset;
assign cond545_in =
  _guard17494 ? idx_between_15_31_reg_out :
  1'd0;
assign cond546_write_en = _guard17495;
assign cond546_clk = clk;
assign cond546_reset = reset;
assign cond546_in =
  _guard17496 ? idx_between_31_32_reg_out :
  1'd0;
assign cond_wire546_in =
  _guard17497 ? idx_between_31_32_reg_out :
  _guard17500 ? cond546_out :
  1'd0;
assign cond568_write_en = _guard17501;
assign cond568_clk = clk;
assign cond568_reset = reset;
assign cond568_in =
  _guard17502 ? idx_between_17_33_reg_out :
  1'd0;
assign cond570_write_en = _guard17503;
assign cond570_clk = clk;
assign cond570_reset = reset;
assign cond570_in =
  _guard17504 ? idx_between_37_38_reg_out :
  1'd0;
assign cond_wire574_in =
  _guard17505 ? idx_between_38_39_reg_out :
  _guard17508 ? cond574_out :
  1'd0;
assign cond586_write_en = _guard17509;
assign cond586_clk = clk;
assign cond586_reset = reset;
assign cond586_in =
  _guard17510 ? idx_between_41_42_reg_out :
  1'd0;
assign cond_wire597_in =
  _guard17513 ? cond597_out :
  _guard17514 ? idx_between_28_44_reg_out :
  1'd0;
assign cond_wire620_in =
  _guard17515 ? idx_between_15_19_reg_out :
  _guard17518 ? cond620_out :
  1'd0;
assign cond_wire634_in =
  _guard17521 ? cond634_out :
  _guard17522 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire639_in =
  _guard17523 ? idx_between_39_40_reg_out :
  _guard17526 ? cond639_out :
  1'd0;
assign cond_wire649_in =
  _guard17527 ? idx_between_22_38_reg_out :
  _guard17530 ? cond649_out :
  1'd0;
assign cond650_write_en = _guard17531;
assign cond650_clk = clk;
assign cond650_reset = reset;
assign cond650_in =
  _guard17532 ? idx_between_26_42_reg_out :
  1'd0;
assign cond_wire654_in =
  _guard17533 ? idx_between_27_43_reg_out :
  _guard17536 ? cond654_out :
  1'd0;
assign cond_wire668_in =
  _guard17537 ? idx_between_31_32_reg_out :
  _guard17540 ? cond668_out :
  1'd0;
assign cond672_write_en = _guard17541;
assign cond672_clk = clk;
assign cond672_reset = reset;
assign cond672_in =
  _guard17542 ? idx_between_32_33_reg_out :
  1'd0;
assign cond677_write_en = _guard17543;
assign cond677_clk = clk;
assign cond677_reset = reset;
assign cond677_in =
  _guard17544 ? idx_between_14_18_reg_out :
  1'd0;
assign cond_wire684_in =
  _guard17547 ? cond684_out :
  _guard17548 ? idx_between_35_36_reg_out :
  1'd0;
assign cond_wire692_in =
  _guard17551 ? cond692_out :
  _guard17552 ? idx_between_37_38_reg_out :
  1'd0;
assign cond_wire693_in =
  _guard17555 ? cond693_out :
  _guard17556 ? idx_between_18_22_reg_out :
  1'd0;
assign cond695_write_en = _guard17557;
assign cond695_clk = clk;
assign cond695_reset = reset;
assign cond695_in =
  _guard17558 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire698_in =
  _guard17559 ? idx_between_19_35_reg_out :
  _guard17562 ? cond698_out :
  1'd0;
assign cond_wire700_in =
  _guard17565 ? cond700_out :
  _guard17566 ? idx_between_39_40_reg_out :
  1'd0;
assign cond702_write_en = _guard17567;
assign cond702_clk = clk;
assign cond702_reset = reset;
assign cond702_in =
  _guard17568 ? idx_between_20_36_reg_out :
  1'd0;
assign cond713_write_en = _guard17569;
assign cond713_clk = clk;
assign cond713_reset = reset;
assign cond713_in =
  _guard17570 ? idx_between_23_27_reg_out :
  1'd0;
assign cond720_write_en = _guard17571;
assign cond720_clk = clk;
assign cond720_reset = reset;
assign cond720_in =
  _guard17572 ? idx_between_44_45_reg_out :
  1'd0;
assign cond_wire725_in =
  _guard17575 ? cond725_out :
  _guard17576 ? idx_between_26_30_reg_out :
  1'd0;
assign cond_wire733_in =
  _guard17577 ? idx_between_32_33_reg_out :
  _guard17580 ? cond733_out :
  1'd0;
assign cond_wire735_in =
  _guard17581 ? idx_between_13_29_reg_out :
  _guard17584 ? cond735_out :
  1'd0;
assign cond752_write_en = _guard17585;
assign cond752_clk = clk;
assign cond752_reset = reset;
assign cond752_in =
  _guard17586 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire752_in =
  _guard17587 ? idx_between_21_37_reg_out :
  _guard17590 ? cond752_out :
  1'd0;
assign cond754_write_en = _guard17591;
assign cond754_clk = clk;
assign cond754_reset = reset;
assign cond754_in =
  _guard17592 ? idx_between_18_22_reg_out :
  1'd0;
assign cond758_write_en = _guard17593;
assign cond758_clk = clk;
assign cond758_reset = reset;
assign cond758_in =
  _guard17594 ? idx_between_19_23_reg_out :
  1'd0;
assign cond_wire788_in =
  _guard17595 ? idx_between_30_46_reg_out :
  _guard17598 ? cond788_out :
  1'd0;
assign cond803_write_en = _guard17599;
assign cond803_clk = clk;
assign cond803_reset = reset;
assign cond803_in =
  _guard17600 ? idx_between_15_19_reg_out :
  1'd0;
assign cond812_write_en = _guard17601;
assign cond812_clk = clk;
assign cond812_reset = reset;
assign cond812_in =
  _guard17602 ? idx_between_17_33_reg_out :
  1'd0;
assign cond_wire815_in =
  _guard17605 ? cond815_out :
  _guard17606 ? idx_between_18_22_reg_out :
  1'd0;
assign cond816_write_en = _guard17607;
assign cond816_clk = clk;
assign cond816_reset = reset;
assign cond816_in =
  _guard17608 ? idx_between_18_34_reg_out :
  1'd0;
assign cond823_write_en = _guard17609;
assign cond823_clk = clk;
assign cond823_reset = reset;
assign cond823_in =
  _guard17610 ? idx_between_20_24_reg_out :
  1'd0;
assign cond_wire832_in =
  _guard17613 ? cond832_out :
  _guard17614 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire837_in =
  _guard17617 ? cond837_out :
  _guard17618 ? idx_between_27_43_reg_out :
  1'd0;
assign cond_wire839_in =
  _guard17621 ? cond839_out :
  _guard17622 ? idx_between_24_28_reg_out :
  1'd0;
assign cond850_write_en = _guard17623;
assign cond850_clk = clk;
assign cond850_reset = reset;
assign cond850_in =
  _guard17624 ? idx_between_46_47_reg_out :
  1'd0;
assign cond857_write_en = _guard17625;
assign cond857_clk = clk;
assign cond857_reset = reset;
assign cond857_in =
  _guard17626 ? idx_between_32_48_reg_out :
  1'd0;
assign cond876_write_en = _guard17627;
assign cond876_clk = clk;
assign cond876_reset = reset;
assign cond876_in =
  _guard17628 ? idx_between_18_22_reg_out :
  1'd0;
assign cond884_write_en = _guard17629;
assign cond884_clk = clk;
assign cond884_reset = reset;
assign cond884_in =
  _guard17630 ? idx_between_20_24_reg_out :
  1'd0;
assign cond_wire885_in =
  _guard17631 ? idx_between_20_36_reg_out :
  _guard17634 ? cond885_out :
  1'd0;
assign cond891_write_en = _guard17635;
assign cond891_clk = clk;
assign cond891_reset = reset;
assign cond891_in =
  _guard17636 ? idx_between_41_42_reg_out :
  1'd0;
assign cond_wire909_in =
  _guard17639 ? cond909_out :
  _guard17640 ? idx_between_26_42_reg_out :
  1'd0;
assign cond910_write_en = _guard17641;
assign cond910_clk = clk;
assign cond910_reset = reset;
assign cond910_in =
  _guard17642 ? idx_between_30_46_reg_out :
  1'd0;
assign cond912_write_en = _guard17643;
assign cond912_clk = clk;
assign cond912_reset = reset;
assign cond912_in =
  _guard17644 ? idx_between_27_31_reg_out :
  1'd0;
assign cond_wire931_in =
  _guard17647 ? cond931_out :
  _guard17648 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire935_in =
  _guard17649 ? idx_between_21_37_reg_out :
  _guard17652 ? cond935_out :
  1'd0;
assign cond946_write_en = _guard17653;
assign cond946_clk = clk;
assign cond946_reset = reset;
assign cond946_in =
  _guard17654 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire952_in =
  _guard17655 ? idx_between_41_42_reg_out :
  _guard17658 ? cond952_out :
  1'd0;
assign cond_wire964_in =
  _guard17659 ? idx_between_44_45_reg_out :
  _guard17662 ? cond964_out :
  1'd0;
assign cond_wire965_in =
  _guard17663 ? idx_between_25_29_reg_out :
  _guard17666 ? cond965_out :
  1'd0;
assign cond_wire989_in =
  _guard17669 ? cond989_out :
  _guard17670 ? idx_between_15_31_reg_out :
  1'd0;
assign cond998_write_en = _guard17671;
assign cond998_clk = clk;
assign cond998_reset = reset;
assign cond998_in =
  _guard17672 ? idx_between_18_22_reg_out :
  1'd0;
assign cond_wire1004_in =
  _guard17673 ? idx_between_23_39_reg_out :
  _guard17676 ? cond1004_out :
  1'd0;
assign cond1007_write_en = _guard17677;
assign cond1007_clk = clk;
assign cond1007_reset = reset;
assign cond1007_in =
  _guard17678 ? idx_between_20_36_reg_out :
  1'd0;
assign cond1008_write_en = _guard17679;
assign cond1008_clk = clk;
assign cond1008_reset = reset;
assign cond1008_in =
  _guard17680 ? idx_between_24_40_reg_out :
  1'd0;
assign cond_wire1010_in =
  _guard17681 ? idx_between_21_25_reg_out :
  _guard17684 ? cond1010_out :
  1'd0;
assign cond_wire1014_in =
  _guard17685 ? idx_between_22_26_reg_out :
  _guard17688 ? cond1014_out :
  1'd0;
assign cond1018_write_en = _guard17689;
assign cond1018_clk = clk;
assign cond1018_reset = reset;
assign cond1018_in =
  _guard17690 ? idx_between_23_27_reg_out :
  1'd0;
assign cond_wire1024_in =
  _guard17693 ? cond1024_out :
  _guard17694 ? idx_between_28_44_reg_out :
  1'd0;
assign cond_wire1027_in =
  _guard17697 ? cond1027_out :
  _guard17698 ? idx_between_25_41_reg_out :
  1'd0;
assign cond1029_write_en = _guard17699;
assign cond1029_clk = clk;
assign cond1029_reset = reset;
assign cond1029_in =
  _guard17700 ? idx_between_45_46_reg_out :
  1'd0;
assign cond_wire1031_in =
  _guard17703 ? cond1031_out :
  _guard17704 ? idx_between_26_42_reg_out :
  1'd0;
assign cond1036_write_en = _guard17705;
assign cond1036_clk = clk;
assign cond1036_reset = reset;
assign cond1036_in =
  _guard17706 ? idx_between_31_47_reg_out :
  1'd0;
assign cond_wire1038_in =
  _guard17707 ? idx_between_28_32_reg_out :
  _guard17710 ? cond1038_out :
  1'd0;
assign adder0_left =
  _guard17711 ? fsm_out :
  1'd0;
assign adder0_right = _guard17712;
assign early_reset_static_seq_go_in = _guard17713;
assign top_0_2_write_en = _guard17716;
assign top_0_2_clk = clk;
assign top_0_2_reset = reset;
assign top_0_2_in = t2_read_data;
assign left_0_8_write_en = _guard17722;
assign left_0_8_clk = clk;
assign left_0_8_reset = reset;
assign left_0_8_in = left_0_7_out;
assign pe_0_11_mul_ready =
  _guard17728 ? 1'd1 :
  _guard17731 ? 1'd0 :
  1'd0;
assign pe_0_11_clk = clk;
assign pe_0_11_top =
  _guard17744 ? top_0_11_out :
  32'd0;
assign pe_0_11_left =
  _guard17757 ? left_0_11_out :
  32'd0;
assign pe_0_11_reset = reset;
assign pe_0_11_go = _guard17770;
assign left_0_14_write_en = _guard17773;
assign left_0_14_clk = clk;
assign left_0_14_reset = reset;
assign left_0_14_in = left_0_13_out;
assign top_1_1_write_en = _guard17779;
assign top_1_1_clk = clk;
assign top_1_1_reset = reset;
assign top_1_1_in = top_0_1_out;
assign left_3_2_write_en = _guard17785;
assign left_3_2_clk = clk;
assign left_3_2_reset = reset;
assign left_3_2_in = left_3_1_out;
assign left_3_4_write_en = _guard17791;
assign left_3_4_clk = clk;
assign left_3_4_reset = reset;
assign left_3_4_in = left_3_3_out;
assign top_4_1_write_en = _guard17797;
assign top_4_1_clk = clk;
assign top_4_1_reset = reset;
assign top_4_1_in = top_3_1_out;
assign top_4_2_write_en = _guard17803;
assign top_4_2_clk = clk;
assign top_4_2_reset = reset;
assign top_4_2_in = top_3_2_out;
assign left_4_15_write_en = _guard17809;
assign left_4_15_clk = clk;
assign left_4_15_reset = reset;
assign left_4_15_in = left_4_14_out;
assign top_5_9_write_en = _guard17815;
assign top_5_9_clk = clk;
assign top_5_9_reset = reset;
assign top_5_9_in = top_4_9_out;
assign top_5_11_write_en = _guard17821;
assign top_5_11_clk = clk;
assign top_5_11_reset = reset;
assign top_5_11_in = top_4_11_out;
assign top_6_4_write_en = _guard17827;
assign top_6_4_clk = clk;
assign top_6_4_reset = reset;
assign top_6_4_in = top_5_4_out;
assign top_6_5_write_en = _guard17833;
assign top_6_5_clk = clk;
assign top_6_5_reset = reset;
assign top_6_5_in = top_5_5_out;
assign left_6_6_write_en = _guard17839;
assign left_6_6_clk = clk;
assign left_6_6_reset = reset;
assign left_6_6_in = left_6_5_out;
assign left_7_2_write_en = _guard17845;
assign left_7_2_clk = clk;
assign left_7_2_reset = reset;
assign left_7_2_in = left_7_1_out;
assign pe_7_5_mul_ready =
  _guard17851 ? 1'd1 :
  _guard17854 ? 1'd0 :
  1'd0;
assign pe_7_5_clk = clk;
assign pe_7_5_top =
  _guard17867 ? top_7_5_out :
  32'd0;
assign pe_7_5_left =
  _guard17880 ? left_7_5_out :
  32'd0;
assign pe_7_5_reset = reset;
assign pe_7_5_go = _guard17893;
assign pe_7_6_mul_ready =
  _guard17896 ? 1'd1 :
  _guard17899 ? 1'd0 :
  1'd0;
assign pe_7_6_clk = clk;
assign pe_7_6_top =
  _guard17912 ? top_7_6_out :
  32'd0;
assign pe_7_6_left =
  _guard17925 ? left_7_6_out :
  32'd0;
assign pe_7_6_reset = reset;
assign pe_7_6_go = _guard17938;
assign top_7_8_write_en = _guard17941;
assign top_7_8_clk = clk;
assign top_7_8_reset = reset;
assign top_7_8_in = top_6_8_out;
assign pe_7_14_mul_ready =
  _guard17947 ? 1'd1 :
  _guard17950 ? 1'd0 :
  1'd0;
assign pe_7_14_clk = clk;
assign pe_7_14_top =
  _guard17963 ? top_7_14_out :
  32'd0;
assign pe_7_14_left =
  _guard17976 ? left_7_14_out :
  32'd0;
assign pe_7_14_reset = reset;
assign pe_7_14_go = _guard17989;
assign pe_8_11_mul_ready =
  _guard17992 ? 1'd1 :
  _guard17995 ? 1'd0 :
  1'd0;
assign pe_8_11_clk = clk;
assign pe_8_11_top =
  _guard18008 ? top_8_11_out :
  32'd0;
assign pe_8_11_left =
  _guard18021 ? left_8_11_out :
  32'd0;
assign pe_8_11_reset = reset;
assign pe_8_11_go = _guard18034;
assign top_8_15_write_en = _guard18037;
assign top_8_15_clk = clk;
assign top_8_15_reset = reset;
assign top_8_15_in = top_7_15_out;
assign pe_9_5_mul_ready =
  _guard18043 ? 1'd1 :
  _guard18046 ? 1'd0 :
  1'd0;
assign pe_9_5_clk = clk;
assign pe_9_5_top =
  _guard18059 ? top_9_5_out :
  32'd0;
assign pe_9_5_left =
  _guard18072 ? left_9_5_out :
  32'd0;
assign pe_9_5_reset = reset;
assign pe_9_5_go = _guard18085;
assign left_9_8_write_en = _guard18088;
assign left_9_8_clk = clk;
assign left_9_8_reset = reset;
assign left_9_8_in = left_9_7_out;
assign pe_10_2_mul_ready =
  _guard18094 ? 1'd1 :
  _guard18097 ? 1'd0 :
  1'd0;
assign pe_10_2_clk = clk;
assign pe_10_2_top =
  _guard18110 ? top_10_2_out :
  32'd0;
assign pe_10_2_left =
  _guard18123 ? left_10_2_out :
  32'd0;
assign pe_10_2_reset = reset;
assign pe_10_2_go = _guard18136;
assign left_10_7_write_en = _guard18139;
assign left_10_7_clk = clk;
assign left_10_7_reset = reset;
assign left_10_7_in = left_10_6_out;
assign pe_11_1_mul_ready =
  _guard18145 ? 1'd1 :
  _guard18148 ? 1'd0 :
  1'd0;
assign pe_11_1_clk = clk;
assign pe_11_1_top =
  _guard18161 ? top_11_1_out :
  32'd0;
assign pe_11_1_left =
  _guard18174 ? left_11_1_out :
  32'd0;
assign pe_11_1_reset = reset;
assign pe_11_1_go = _guard18187;
assign top_11_13_write_en = _guard18190;
assign top_11_13_clk = clk;
assign top_11_13_reset = reset;
assign top_11_13_in = top_10_13_out;
assign left_11_14_write_en = _guard18196;
assign left_11_14_clk = clk;
assign left_11_14_reset = reset;
assign left_11_14_in = left_11_13_out;
assign pe_12_6_mul_ready =
  _guard18202 ? 1'd1 :
  _guard18205 ? 1'd0 :
  1'd0;
assign pe_12_6_clk = clk;
assign pe_12_6_top =
  _guard18218 ? top_12_6_out :
  32'd0;
assign pe_12_6_left =
  _guard18231 ? left_12_6_out :
  32'd0;
assign pe_12_6_reset = reset;
assign pe_12_6_go = _guard18244;
assign top_12_6_write_en = _guard18247;
assign top_12_6_clk = clk;
assign top_12_6_reset = reset;
assign top_12_6_in = top_11_6_out;
assign top_12_8_write_en = _guard18253;
assign top_12_8_clk = clk;
assign top_12_8_reset = reset;
assign top_12_8_in = top_11_8_out;
assign left_12_15_write_en = _guard18259;
assign left_12_15_clk = clk;
assign left_12_15_reset = reset;
assign left_12_15_in = left_12_14_out;
assign pe_13_4_mul_ready =
  _guard18265 ? 1'd1 :
  _guard18268 ? 1'd0 :
  1'd0;
assign pe_13_4_clk = clk;
assign pe_13_4_top =
  _guard18281 ? top_13_4_out :
  32'd0;
assign pe_13_4_left =
  _guard18294 ? left_13_4_out :
  32'd0;
assign pe_13_4_reset = reset;
assign pe_13_4_go = _guard18307;
assign top_13_11_write_en = _guard18310;
assign top_13_11_clk = clk;
assign top_13_11_reset = reset;
assign top_13_11_in = top_12_11_out;
assign top_13_13_write_en = _guard18316;
assign top_13_13_clk = clk;
assign top_13_13_reset = reset;
assign top_13_13_in = top_12_13_out;
assign pe_14_6_mul_ready =
  _guard18322 ? 1'd1 :
  _guard18325 ? 1'd0 :
  1'd0;
assign pe_14_6_clk = clk;
assign pe_14_6_top =
  _guard18338 ? top_14_6_out :
  32'd0;
assign pe_14_6_left =
  _guard18351 ? left_14_6_out :
  32'd0;
assign pe_14_6_reset = reset;
assign pe_14_6_go = _guard18364;
assign pe_15_4_mul_ready =
  _guard18367 ? 1'd1 :
  _guard18370 ? 1'd0 :
  1'd0;
assign pe_15_4_clk = clk;
assign pe_15_4_top =
  _guard18383 ? top_15_4_out :
  32'd0;
assign pe_15_4_left =
  _guard18396 ? left_15_4_out :
  32'd0;
assign pe_15_4_reset = reset;
assign pe_15_4_go = _guard18409;
assign left_15_6_write_en = _guard18412;
assign left_15_6_clk = clk;
assign left_15_6_reset = reset;
assign left_15_6_in = left_15_5_out;
assign top_15_14_write_en = _guard18418;
assign top_15_14_clk = clk;
assign top_15_14_reset = reset;
assign top_15_14_in = top_14_14_out;
assign t0_add_left = 5'd1;
assign t0_add_right = t0_idx_out;
assign l0_add_left = 5'd1;
assign l0_add_right = l0_idx_out;
assign index_lt_20_left = idx_add_out;
assign index_lt_20_right = 6'd20;
assign index_lt_46_left = idx_add_out;
assign index_lt_46_right = 6'd46;
assign index_lt_21_left = idx_add_out;
assign index_lt_21_right = 6'd21;
assign idx_between_23_27_reg_write_en = _guard18444;
assign idx_between_23_27_reg_clk = clk;
assign idx_between_23_27_reg_reset = reset;
assign idx_between_23_27_reg_in =
  _guard18445 ? idx_between_23_27_comb_out :
  _guard18448 ? 1'd0 :
  'x;
assign index_ge_23_left = idx_add_out;
assign index_ge_23_right = 6'd23;
assign index_ge_33_left = idx_add_out;
assign index_ge_33_right = 6'd33;
assign idx_between_20_24_reg_write_en = _guard18457;
assign idx_between_20_24_reg_clk = clk;
assign idx_between_20_24_reg_reset = reset;
assign idx_between_20_24_reg_in =
  _guard18458 ? idx_between_20_24_comb_out :
  _guard18461 ? 1'd0 :
  'x;
assign index_lt_39_left = idx_add_out;
assign index_lt_39_right = 6'd39;
assign idx_between_30_34_reg_write_en = _guard18468;
assign idx_between_30_34_reg_clk = clk;
assign idx_between_30_34_reg_reset = reset;
assign idx_between_30_34_reg_in =
  _guard18469 ? idx_between_30_34_comb_out :
  _guard18472 ? 1'd0 :
  'x;
assign idx_between_14_30_comb_left = index_ge_14_out;
assign idx_between_14_30_comb_right = index_lt_30_out;
assign index_ge_28_left = idx_add_out;
assign index_ge_28_right = 6'd28;
assign index_lt_33_left = idx_add_out;
assign index_lt_33_right = 6'd33;
assign index_ge_11_left = idx_add_out;
assign index_ge_11_right = 6'd11;
assign idx_between_12_28_reg_write_en = _guard18485;
assign idx_between_12_28_reg_clk = clk;
assign idx_between_12_28_reg_reset = reset;
assign idx_between_12_28_reg_in =
  _guard18488 ? 1'd0 :
  _guard18489 ? idx_between_12_28_comb_out :
  'x;
assign idx_between_4_8_comb_left = index_ge_4_out;
assign idx_between_4_8_comb_right = index_lt_8_out;
assign index_ge_9_left = idx_add_out;
assign index_ge_9_right = 6'd9;
assign idx_between_9_25_comb_left = index_ge_9_out;
assign idx_between_9_25_comb_right = index_lt_25_out;
assign idx_between_11_15_comb_left = index_ge_11_out;
assign idx_between_11_15_comb_right = index_lt_15_out;
assign cond_wire2_in =
  _guard18498 ? idx_between_5_21_reg_out :
  _guard18501 ? cond2_out :
  1'd0;
assign cond_wire9_in =
  _guard18502 ? idx_between_2_18_reg_out :
  _guard18505 ? cond9_out :
  1'd0;
assign cond10_write_en = _guard18506;
assign cond10_clk = clk;
assign cond10_reset = reset;
assign cond10_in =
  _guard18507 ? idx_between_3_7_reg_out :
  1'd0;
assign cond_wire11_in =
  _guard18510 ? cond11_out :
  _guard18511 ? idx_between_3_19_reg_out :
  1'd0;
assign cond21_write_en = _guard18512;
assign cond21_clk = clk;
assign cond21_reset = reset;
assign cond21_in =
  _guard18513 ? idx_between_5_21_reg_out :
  1'd0;
assign cond24_write_en = _guard18514;
assign cond24_clk = clk;
assign cond24_reset = reset;
assign cond24_in =
  _guard18515 ? idx_between_5_21_reg_out :
  1'd0;
assign cond31_write_en = _guard18516;
assign cond31_clk = clk;
assign cond31_reset = reset;
assign cond31_in =
  _guard18517 ? idx_between_7_23_reg_out :
  1'd0;
assign cond36_write_en = _guard18518;
assign cond36_clk = clk;
assign cond36_reset = reset;
assign cond36_in =
  _guard18519 ? idx_between_8_24_reg_out :
  1'd0;
assign cond_wire41_in =
  _guard18522 ? cond41_out :
  _guard18523 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire45_in =
  _guard18526 ? cond45_out :
  _guard18527 ? idx_between_10_14_reg_out :
  1'd0;
assign cond51_write_en = _guard18528;
assign cond51_clk = clk;
assign cond51_reset = reset;
assign cond51_in =
  _guard18529 ? idx_between_11_27_reg_out :
  1'd0;
assign cond_wire57_in =
  _guard18530 ? idx_between_16_32_reg_out :
  _guard18533 ? cond57_out :
  1'd0;
assign cond_wire58_in =
  _guard18534 ? idx_between_32_33_reg_out :
  _guard18537 ? cond58_out :
  1'd0;
assign cond61_write_en = _guard18538;
assign cond61_clk = clk;
assign cond61_reset = reset;
assign cond61_in =
  _guard18539 ? idx_between_13_29_reg_out :
  1'd0;
assign cond80_write_en = _guard18540;
assign cond80_clk = clk;
assign cond80_reset = reset;
assign cond80_in =
  _guard18541 ? idx_between_2_6_reg_out :
  1'd0;
assign cond_wire80_in =
  _guard18544 ? cond80_out :
  _guard18545 ? idx_between_2_6_reg_out :
  1'd0;
assign cond86_write_en = _guard18546;
assign cond86_clk = clk;
assign cond86_reset = reset;
assign cond86_in =
  _guard18547 ? idx_between_7_23_reg_out :
  1'd0;
assign cond97_write_en = _guard18548;
assign cond97_clk = clk;
assign cond97_reset = reset;
assign cond97_in =
  _guard18549 ? idx_between_6_22_reg_out :
  1'd0;
assign cond_wire123_in =
  _guard18552 ? cond123_out :
  _guard18553 ? idx_between_32_33_reg_out :
  1'd0;
assign cond127_write_en = _guard18554;
assign cond127_clk = clk;
assign cond127_reset = reset;
assign cond127_in =
  _guard18555 ? idx_between_33_34_reg_out :
  1'd0;
assign cond129_write_en = _guard18556;
assign cond129_clk = clk;
assign cond129_reset = reset;
assign cond129_in =
  _guard18557 ? idx_between_14_30_reg_out :
  1'd0;
assign cond_wire129_in =
  _guard18558 ? idx_between_14_30_reg_out :
  _guard18561 ? cond129_out :
  1'd0;
assign cond_wire136_in =
  _guard18562 ? idx_between_16_20_reg_out :
  _guard18565 ? cond136_out :
  1'd0;
assign cond_wire145_in =
  _guard18566 ? idx_between_3_7_reg_out :
  _guard18569 ? cond145_out :
  1'd0;
assign cond170_write_en = _guard18570;
assign cond170_clk = clk;
assign cond170_reset = reset;
assign cond170_in =
  _guard18571 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire184_in =
  _guard18572 ? idx_between_32_33_reg_out :
  _guard18575 ? cond184_out :
  1'd0;
assign cond_wire194_in =
  _guard18578 ? cond194_out :
  _guard18579 ? idx_between_15_31_reg_out :
  1'd0;
assign cond199_write_en = _guard18580;
assign cond199_clk = clk;
assign cond199_reset = reset;
assign cond199_in =
  _guard18581 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire201_in =
  _guard18582 ? idx_between_17_21_reg_out :
  _guard18585 ? cond201_out :
  1'd0;
assign cond211_write_en = _guard18586;
assign cond211_clk = clk;
assign cond211_reset = reset;
assign cond211_in =
  _guard18587 ? idx_between_4_20_reg_out :
  1'd0;
assign cond_wire220_in =
  _guard18590 ? cond220_out :
  _guard18591 ? idx_between_10_26_reg_out :
  1'd0;
assign cond242_write_en = _guard18592;
assign cond242_clk = clk;
assign cond242_reset = reset;
assign cond242_in =
  _guard18593 ? idx_between_12_16_reg_out :
  1'd0;
assign cond_wire242_in =
  _guard18596 ? cond242_out :
  _guard18597 ? idx_between_12_16_reg_out :
  1'd0;
assign cond_wire246_in =
  _guard18598 ? idx_between_13_17_reg_out :
  _guard18601 ? cond246_out :
  1'd0;
assign cond249_write_en = _guard18602;
assign cond249_clk = clk;
assign cond249_reset = reset;
assign cond249_in =
  _guard18603 ? idx_between_33_34_reg_out :
  1'd0;
assign cond_wire249_in =
  _guard18606 ? cond249_out :
  _guard18607 ? idx_between_33_34_reg_out :
  1'd0;
assign cond_wire250_in =
  _guard18608 ? idx_between_14_18_reg_out :
  _guard18611 ? cond250_out :
  1'd0;
assign cond_wire251_in =
  _guard18614 ? cond251_out :
  _guard18615 ? idx_between_14_30_reg_out :
  1'd0;
assign cond268_write_en = _guard18616;
assign cond268_clk = clk;
assign cond268_reset = reset;
assign cond268_in =
  _guard18617 ? idx_between_22_38_reg_out :
  1'd0;
assign cond269_write_en = _guard18618;
assign cond269_clk = clk;
assign cond269_reset = reset;
assign cond269_in =
  _guard18619 ? idx_between_38_39_reg_out :
  1'd0;
assign cond274_write_en = _guard18620;
assign cond274_clk = clk;
assign cond274_reset = reset;
assign cond274_in =
  _guard18621 ? idx_between_4_20_reg_out :
  1'd0;
assign cond_wire288_in =
  _guard18624 ? cond288_out :
  _guard18625 ? idx_between_8_24_reg_out :
  1'd0;
assign cond292_write_en = _guard18626;
assign cond292_clk = clk;
assign cond292_reset = reset;
assign cond292_in =
  _guard18627 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire294_in =
  _guard18628 ? idx_between_29_30_reg_out :
  _guard18631 ? cond294_out :
  1'd0;
assign cond_wire299_in =
  _guard18634 ? cond299_out :
  _guard18635 ? idx_between_11_15_reg_out :
  1'd0;
assign cond301_write_en = _guard18636;
assign cond301_clk = clk;
assign cond301_reset = reset;
assign cond301_in =
  _guard18637 ? idx_between_15_31_reg_out :
  1'd0;
assign cond332_write_en = _guard18638;
assign cond332_clk = clk;
assign cond332_reset = reset;
assign cond332_in =
  _guard18639 ? idx_between_19_35_reg_out :
  1'd0;
assign cond335_write_en = _guard18640;
assign cond335_clk = clk;
assign cond335_reset = reset;
assign cond335_in =
  _guard18641 ? idx_between_20_24_reg_out :
  1'd0;
assign cond344_write_en = _guard18642;
assign cond344_clk = clk;
assign cond344_reset = reset;
assign cond344_in =
  _guard18643 ? idx_between_7_11_reg_out :
  1'd0;
assign cond_wire347_in =
  _guard18644 ? idx_between_27_28_reg_out :
  _guard18647 ? cond347_out :
  1'd0;
assign cond_wire379_in =
  _guard18650 ? cond379_out :
  _guard18651 ? idx_between_35_36_reg_out :
  1'd0;
assign cond_wire385_in =
  _guard18652 ? idx_between_17_33_reg_out :
  _guard18655 ? cond385_out :
  1'd0;
assign cond396_write_en = _guard18656;
assign cond396_clk = clk;
assign cond396_reset = reset;
assign cond396_in =
  _guard18657 ? idx_between_20_24_reg_out :
  1'd0;
assign cond405_write_en = _guard18658;
assign cond405_clk = clk;
assign cond405_reset = reset;
assign cond405_in =
  _guard18659 ? idx_between_7_11_reg_out :
  1'd0;
assign cond_wire434_in =
  _guard18660 ? idx_between_14_30_reg_out :
  _guard18663 ? cond434_out :
  1'd0;
assign cond_wire440_in =
  _guard18666 ? cond440_out :
  _guard18667 ? idx_between_35_36_reg_out :
  1'd0;
assign cond441_write_en = _guard18668;
assign cond441_clk = clk;
assign cond441_reset = reset;
assign cond441_in =
  _guard18669 ? idx_between_16_20_reg_out :
  1'd0;
assign cond454_write_en = _guard18670;
assign cond454_clk = clk;
assign cond454_reset = reset;
assign cond454_in =
  _guard18671 ? idx_between_19_35_reg_out :
  1'd0;
assign cond466_write_en = _guard18672;
assign cond466_clk = clk;
assign cond466_reset = reset;
assign cond466_in =
  _guard18673 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire484_in =
  _guard18676 ? cond484_out :
  _guard18677 ? idx_between_15_31_reg_out :
  1'd0;
assign cond497_write_en = _guard18678;
assign cond497_clk = clk;
assign cond497_reset = reset;
assign cond497_in =
  _guard18679 ? idx_between_34_35_reg_out :
  1'd0;
assign cond_wire501_in =
  _guard18682 ? cond501_out :
  _guard18683 ? idx_between_35_36_reg_out :
  1'd0;
assign cond502_write_en = _guard18684;
assign cond502_clk = clk;
assign cond502_reset = reset;
assign cond502_in =
  _guard18685 ? idx_between_16_20_reg_out :
  1'd0;
assign cond514_write_en = _guard18686;
assign cond514_clk = clk;
assign cond514_reset = reset;
assign cond514_in =
  _guard18687 ? idx_between_19_23_reg_out :
  1'd0;
assign cond515_write_en = _guard18688;
assign cond515_clk = clk;
assign cond515_reset = reset;
assign cond515_in =
  _guard18689 ? idx_between_19_35_reg_out :
  1'd0;
assign cond531_write_en = _guard18690;
assign cond531_clk = clk;
assign cond531_reset = reset;
assign cond531_in =
  _guard18691 ? idx_between_23_39_reg_out :
  1'd0;
assign cond_wire534_in =
  _guard18692 ? idx_between_8_24_reg_out :
  _guard18695 ? cond534_out :
  1'd0;
assign cond548_write_en = _guard18696;
assign cond548_clk = clk;
assign cond548_reset = reset;
assign cond548_in =
  _guard18697 ? idx_between_12_28_reg_out :
  1'd0;
assign cond553_write_en = _guard18698;
assign cond553_clk = clk;
assign cond553_reset = reset;
assign cond553_in =
  _guard18699 ? idx_between_17_33_reg_out :
  1'd0;
assign cond556_write_en = _guard18700;
assign cond556_clk = clk;
assign cond556_reset = reset;
assign cond556_in =
  _guard18701 ? idx_between_14_30_reg_out :
  1'd0;
assign cond558_write_en = _guard18702;
assign cond558_clk = clk;
assign cond558_reset = reset;
assign cond558_in =
  _guard18703 ? idx_between_34_35_reg_out :
  1'd0;
assign cond559_write_en = _guard18704;
assign cond559_clk = clk;
assign cond559_reset = reset;
assign cond559_in =
  _guard18705 ? idx_between_15_19_reg_out :
  1'd0;
assign cond_wire572_in =
  _guard18708 ? cond572_out :
  _guard18709 ? idx_between_18_34_reg_out :
  1'd0;
assign cond579_write_en = _guard18710;
assign cond579_clk = clk;
assign cond579_reset = reset;
assign cond579_in =
  _guard18711 ? idx_between_20_24_reg_out :
  1'd0;
assign cond_wire588_in =
  _guard18714 ? cond588_out :
  _guard18715 ? idx_between_22_38_reg_out :
  1'd0;
assign cond604_write_en = _guard18716;
assign cond604_clk = clk;
assign cond604_reset = reset;
assign cond604_in =
  _guard18717 ? idx_between_11_15_reg_out :
  1'd0;
assign cond607_write_en = _guard18718;
assign cond607_clk = clk;
assign cond607_reset = reset;
assign cond607_in =
  _guard18719 ? idx_between_31_32_reg_out :
  1'd0;
assign cond608_write_en = _guard18720;
assign cond608_clk = clk;
assign cond608_reset = reset;
assign cond608_in =
  _guard18721 ? idx_between_12_16_reg_out :
  1'd0;
assign cond_wire616_in =
  _guard18722 ? idx_between_14_18_reg_out :
  _guard18725 ? cond616_out :
  1'd0;
assign cond618_write_en = _guard18726;
assign cond618_clk = clk;
assign cond618_reset = reset;
assign cond618_in =
  _guard18727 ? idx_between_18_34_reg_out :
  1'd0;
assign cond626_write_en = _guard18728;
assign cond626_clk = clk;
assign cond626_reset = reset;
assign cond626_in =
  _guard18729 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire632_in =
  _guard18732 ? cond632_out :
  _guard18733 ? idx_between_18_22_reg_out :
  1'd0;
assign cond638_write_en = _guard18734;
assign cond638_clk = clk;
assign cond638_reset = reset;
assign cond638_in =
  _guard18735 ? idx_between_23_39_reg_out :
  1'd0;
assign cond643_write_en = _guard18736;
assign cond643_clk = clk;
assign cond643_reset = reset;
assign cond643_in =
  _guard18737 ? idx_between_40_41_reg_out :
  1'd0;
assign cond644_write_en = _guard18738;
assign cond644_clk = clk;
assign cond644_reset = reset;
assign cond644_in =
  _guard18739 ? idx_between_21_25_reg_out :
  1'd0;
assign cond_wire646_in =
  _guard18742 ? cond646_out :
  _guard18743 ? idx_between_25_41_reg_out :
  1'd0;
assign cond_wire660_in =
  _guard18746 ? cond660_out :
  _guard18747 ? idx_between_25_29_reg_out :
  1'd0;
assign cond_wire662_in =
  _guard18748 ? idx_between_29_45_reg_out :
  _guard18751 ? cond662_out :
  1'd0;
assign cond_wire663_in =
  _guard18754 ? cond663_out :
  _guard18755 ? idx_between_45_46_reg_out :
  1'd0;
assign cond_wire667_in =
  _guard18758 ? cond667_out :
  _guard18759 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire670_in =
  _guard18762 ? cond670_out :
  _guard18763 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire681_in =
  _guard18764 ? idx_between_15_19_reg_out :
  _guard18767 ? cond681_out :
  1'd0;
assign cond_wire683_in =
  _guard18770 ? cond683_out :
  _guard18771 ? idx_between_19_35_reg_out :
  1'd0;
assign cond694_write_en = _guard18772;
assign cond694_clk = clk;
assign cond694_reset = reset;
assign cond694_in =
  _guard18773 ? idx_between_18_34_reg_out :
  1'd0;
assign cond_wire696_in =
  _guard18776 ? cond696_out :
  _guard18777 ? idx_between_38_39_reg_out :
  1'd0;
assign cond705_write_en = _guard18778;
assign cond705_clk = clk;
assign cond705_reset = reset;
assign cond705_in =
  _guard18779 ? idx_between_21_25_reg_out :
  1'd0;
assign cond_wire713_in =
  _guard18782 ? cond713_out :
  _guard18783 ? idx_between_23_27_reg_out :
  1'd0;
assign cond_wire720_in =
  _guard18784 ? idx_between_44_45_reg_out :
  _guard18787 ? cond720_out :
  1'd0;
assign cond_wire723_in =
  _guard18790 ? cond723_out :
  _guard18791 ? idx_between_29_45_reg_out :
  1'd0;
assign cond_wire726_in =
  _guard18792 ? idx_between_26_42_reg_out :
  _guard18795 ? cond726_out :
  1'd0;
assign cond727_write_en = _guard18796;
assign cond727_clk = clk;
assign cond727_reset = reset;
assign cond727_in =
  _guard18797 ? idx_between_30_46_reg_out :
  1'd0;
assign cond734_write_en = _guard18798;
assign cond734_clk = clk;
assign cond734_reset = reset;
assign cond734_in =
  _guard18799 ? idx_between_13_17_reg_out :
  1'd0;
assign cond740_write_en = _guard18800;
assign cond740_clk = clk;
assign cond740_reset = reset;
assign cond740_in =
  _guard18801 ? idx_between_18_34_reg_out :
  1'd0;
assign cond_wire741_in =
  _guard18802 ? idx_between_34_35_reg_out :
  _guard18805 ? cond741_out :
  1'd0;
assign cond744_write_en = _guard18806;
assign cond744_clk = clk;
assign cond744_reset = reset;
assign cond744_in =
  _guard18807 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire751_in =
  _guard18808 ? idx_between_17_33_reg_out :
  _guard18811 ? cond751_out :
  1'd0;
assign cond772_write_en = _guard18812;
assign cond772_clk = clk;
assign cond772_reset = reset;
assign cond772_in =
  _guard18813 ? idx_between_26_42_reg_out :
  1'd0;
assign cond_wire773_in =
  _guard18814 ? idx_between_42_43_reg_out :
  _guard18817 ? cond773_out :
  1'd0;
assign cond_wire776_in =
  _guard18820 ? cond776_out :
  _guard18821 ? idx_between_27_43_reg_out :
  1'd0;
assign cond_wire808_in =
  _guard18822 ? idx_between_16_32_reg_out :
  _guard18825 ? cond808_out :
  1'd0;
assign cond813_write_en = _guard18826;
assign cond813_clk = clk;
assign cond813_reset = reset;
assign cond813_in =
  _guard18827 ? idx_between_21_37_reg_out :
  1'd0;
assign cond821_write_en = _guard18828;
assign cond821_clk = clk;
assign cond821_reset = reset;
assign cond821_in =
  _guard18829 ? idx_between_23_39_reg_out :
  1'd0;
assign cond832_write_en = _guard18830;
assign cond832_clk = clk;
assign cond832_reset = reset;
assign cond832_in =
  _guard18831 ? idx_between_22_38_reg_out :
  1'd0;
assign cond845_write_en = _guard18832;
assign cond845_clk = clk;
assign cond845_reset = reset;
assign cond845_in =
  _guard18833 ? idx_between_29_45_reg_out :
  1'd0;
assign cond_wire856_in =
  _guard18836 ? cond856_out :
  _guard18837 ? idx_between_28_44_reg_out :
  1'd0;
assign cond_wire865_in =
  _guard18840 ? cond865_out :
  _guard18841 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire915_in =
  _guard18842 ? idx_between_47_48_reg_out :
  _guard18845 ? cond915_out :
  1'd0;
assign cond926_write_en = _guard18846;
assign cond926_clk = clk;
assign cond926_reset = reset;
assign cond926_in =
  _guard18847 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire943_in =
  _guard18850 ? cond943_out :
  _guard18851 ? idx_between_23_39_reg_out :
  1'd0;
assign cond_wire948_in =
  _guard18852 ? idx_between_40_41_reg_out :
  _guard18855 ? cond948_out :
  1'd0;
assign cond_wire956_in =
  _guard18856 ? idx_between_42_43_reg_out :
  _guard18859 ? cond956_out :
  1'd0;
assign cond961_write_en = _guard18860;
assign cond961_clk = clk;
assign cond961_reset = reset;
assign cond961_in =
  _guard18861 ? idx_between_24_28_reg_out :
  1'd0;
assign cond_wire961_in =
  _guard18864 ? cond961_out :
  _guard18865 ? idx_between_24_28_reg_out :
  1'd0;
assign cond_wire979_in =
  _guard18868 ? cond979_out :
  _guard18869 ? idx_between_32_48_reg_out :
  1'd0;
assign cond_wire983_in =
  _guard18870 ? idx_between_33_49_reg_out :
  _guard18873 ? cond983_out :
  1'd0;
assign cond_wire985_in =
  _guard18876 ? cond985_out :
  _guard18877 ? idx_between_30_34_reg_out :
  1'd0;
assign cond_wire999_in =
  _guard18878 ? idx_between_18_34_reg_out :
  _guard18881 ? cond999_out :
  1'd0;
assign cond_wire1003_in =
  _guard18884 ? cond1003_out :
  _guard18885 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire1006_in =
  _guard18888 ? cond1006_out :
  _guard18889 ? idx_between_20_24_reg_out :
  1'd0;
assign cond1026_write_en = _guard18890;
assign cond1026_clk = clk;
assign cond1026_reset = reset;
assign cond1026_in =
  _guard18891 ? idx_between_25_29_reg_out :
  1'd0;
assign cond1037_write_en = _guard18892;
assign cond1037_clk = clk;
assign cond1037_reset = reset;
assign cond1037_in =
  _guard18893 ? idx_between_47_48_reg_out :
  1'd0;
assign cond_wire1044_in =
  _guard18896 ? cond1044_out :
  _guard18897 ? idx_between_33_49_reg_out :
  1'd0;
assign cond_wire1048_in =
  _guard18898 ? idx_between_34_50_reg_out :
  _guard18901 ? cond1048_out :
  1'd0;
assign cond1051_write_en = _guard18902;
assign cond1051_clk = clk;
assign cond1051_reset = reset;
assign cond1051_in =
  _guard18903 ? idx_between_35_51_reg_out :
  1'd0;
assign signal_reg_write_en = _guard18913;
assign signal_reg_clk = clk;
assign signal_reg_reset = reset;
assign signal_reg_in =
  _guard18919 ? 1'd1 :
  _guard18922 ? 1'd0 :
  1'd0;
assign top_0_4_write_en = _guard18925;
assign top_0_4_clk = clk;
assign top_0_4_reset = reset;
assign top_0_4_in = t4_read_data;
assign left_0_5_write_en = _guard18931;
assign left_0_5_clk = clk;
assign left_0_5_reset = reset;
assign left_0_5_in = left_0_4_out;
assign top_0_10_write_en = _guard18937;
assign top_0_10_clk = clk;
assign top_0_10_reset = reset;
assign top_0_10_in = t10_read_data;
assign pe_1_11_mul_ready =
  _guard18943 ? 1'd1 :
  _guard18946 ? 1'd0 :
  1'd0;
assign pe_1_11_clk = clk;
assign pe_1_11_top =
  _guard18959 ? top_1_11_out :
  32'd0;
assign pe_1_11_left =
  _guard18972 ? left_1_11_out :
  32'd0;
assign pe_1_11_reset = reset;
assign pe_1_11_go = _guard18985;
assign left_1_12_write_en = _guard18988;
assign left_1_12_clk = clk;
assign left_1_12_reset = reset;
assign left_1_12_in = left_1_11_out;
assign pe_2_0_mul_ready =
  _guard18994 ? 1'd1 :
  _guard18997 ? 1'd0 :
  1'd0;
assign pe_2_0_clk = clk;
assign pe_2_0_top =
  _guard19010 ? top_2_0_out :
  32'd0;
assign pe_2_0_left =
  _guard19023 ? left_2_0_out :
  32'd0;
assign pe_2_0_reset = reset;
assign pe_2_0_go = _guard19036;
assign left_2_1_write_en = _guard19039;
assign left_2_1_clk = clk;
assign left_2_1_reset = reset;
assign left_2_1_in = left_2_0_out;
assign top_2_2_write_en = _guard19045;
assign top_2_2_clk = clk;
assign top_2_2_reset = reset;
assign top_2_2_in = top_1_2_out;
assign left_2_5_write_en = _guard19051;
assign left_2_5_clk = clk;
assign left_2_5_reset = reset;
assign left_2_5_in = left_2_4_out;
assign left_3_6_write_en = _guard19057;
assign left_3_6_clk = clk;
assign left_3_6_reset = reset;
assign left_3_6_in = left_3_5_out;
assign left_3_8_write_en = _guard19063;
assign left_3_8_clk = clk;
assign left_3_8_reset = reset;
assign left_3_8_in = left_3_7_out;
assign pe_3_12_mul_ready =
  _guard19069 ? 1'd1 :
  _guard19072 ? 1'd0 :
  1'd0;
assign pe_3_12_clk = clk;
assign pe_3_12_top =
  _guard19085 ? top_3_12_out :
  32'd0;
assign pe_3_12_left =
  _guard19098 ? left_3_12_out :
  32'd0;
assign pe_3_12_reset = reset;
assign pe_3_12_go = _guard19111;
assign top_3_12_write_en = _guard19114;
assign top_3_12_clk = clk;
assign top_3_12_reset = reset;
assign top_3_12_in = top_2_12_out;
assign left_3_15_write_en = _guard19120;
assign left_3_15_clk = clk;
assign left_3_15_reset = reset;
assign left_3_15_in = left_3_14_out;
assign pe_4_4_mul_ready =
  _guard19126 ? 1'd1 :
  _guard19129 ? 1'd0 :
  1'd0;
assign pe_4_4_clk = clk;
assign pe_4_4_top =
  _guard19142 ? top_4_4_out :
  32'd0;
assign pe_4_4_left =
  _guard19155 ? left_4_4_out :
  32'd0;
assign pe_4_4_reset = reset;
assign pe_4_4_go = _guard19168;
assign left_4_4_write_en = _guard19171;
assign left_4_4_clk = clk;
assign left_4_4_reset = reset;
assign left_4_4_in = left_4_3_out;
assign pe_4_7_mul_ready =
  _guard19177 ? 1'd1 :
  _guard19180 ? 1'd0 :
  1'd0;
assign pe_4_7_clk = clk;
assign pe_4_7_top =
  _guard19193 ? top_4_7_out :
  32'd0;
assign pe_4_7_left =
  _guard19206 ? left_4_7_out :
  32'd0;
assign pe_4_7_reset = reset;
assign pe_4_7_go = _guard19219;
assign top_4_11_write_en = _guard19222;
assign top_4_11_clk = clk;
assign top_4_11_reset = reset;
assign top_4_11_in = top_3_11_out;
assign top_4_12_write_en = _guard19228;
assign top_4_12_clk = clk;
assign top_4_12_reset = reset;
assign top_4_12_in = top_3_12_out;
assign pe_4_13_mul_ready =
  _guard19234 ? 1'd1 :
  _guard19237 ? 1'd0 :
  1'd0;
assign pe_4_13_clk = clk;
assign pe_4_13_top =
  _guard19250 ? top_4_13_out :
  32'd0;
assign pe_4_13_left =
  _guard19263 ? left_4_13_out :
  32'd0;
assign pe_4_13_reset = reset;
assign pe_4_13_go = _guard19276;
assign left_5_5_write_en = _guard19279;
assign left_5_5_clk = clk;
assign left_5_5_reset = reset;
assign left_5_5_in = left_5_4_out;
assign left_5_9_write_en = _guard19285;
assign left_5_9_clk = clk;
assign left_5_9_reset = reset;
assign left_5_9_in = left_5_8_out;
assign top_5_10_write_en = _guard19291;
assign top_5_10_clk = clk;
assign top_5_10_reset = reset;
assign top_5_10_in = top_4_10_out;
assign pe_5_14_mul_ready =
  _guard19297 ? 1'd1 :
  _guard19300 ? 1'd0 :
  1'd0;
assign pe_5_14_clk = clk;
assign pe_5_14_top =
  _guard19313 ? top_5_14_out :
  32'd0;
assign pe_5_14_left =
  _guard19326 ? left_5_14_out :
  32'd0;
assign pe_5_14_reset = reset;
assign pe_5_14_go = _guard19339;
assign left_5_15_write_en = _guard19342;
assign left_5_15_clk = clk;
assign left_5_15_reset = reset;
assign left_5_15_in = left_5_14_out;
assign left_6_10_write_en = _guard19348;
assign left_6_10_clk = clk;
assign left_6_10_reset = reset;
assign left_6_10_in = left_6_9_out;
assign left_7_0_write_en = _guard19354;
assign left_7_0_clk = clk;
assign left_7_0_reset = reset;
assign left_7_0_in = l7_read_data;
assign top_7_3_write_en = _guard19360;
assign top_7_3_clk = clk;
assign top_7_3_reset = reset;
assign top_7_3_in = top_6_3_out;
assign top_7_6_write_en = _guard19366;
assign top_7_6_clk = clk;
assign top_7_6_reset = reset;
assign top_7_6_in = top_6_6_out;
assign left_7_10_write_en = _guard19372;
assign left_7_10_clk = clk;
assign left_7_10_reset = reset;
assign left_7_10_in = left_7_9_out;
assign left_8_0_write_en = _guard19378;
assign left_8_0_clk = clk;
assign left_8_0_reset = reset;
assign left_8_0_in = l8_read_data;
assign left_8_6_write_en = _guard19384;
assign left_8_6_clk = clk;
assign left_8_6_reset = reset;
assign left_8_6_in = left_8_5_out;
assign pe_9_1_mul_ready =
  _guard19390 ? 1'd1 :
  _guard19393 ? 1'd0 :
  1'd0;
assign pe_9_1_clk = clk;
assign pe_9_1_top =
  _guard19406 ? top_9_1_out :
  32'd0;
assign pe_9_1_left =
  _guard19419 ? left_9_1_out :
  32'd0;
assign pe_9_1_reset = reset;
assign pe_9_1_go = _guard19432;
assign top_9_3_write_en = _guard19435;
assign top_9_3_clk = clk;
assign top_9_3_reset = reset;
assign top_9_3_in = top_8_3_out;
assign left_9_7_write_en = _guard19441;
assign left_9_7_clk = clk;
assign left_9_7_reset = reset;
assign left_9_7_in = left_9_6_out;
assign pe_9_8_mul_ready =
  _guard19447 ? 1'd1 :
  _guard19450 ? 1'd0 :
  1'd0;
assign pe_9_8_clk = clk;
assign pe_9_8_top =
  _guard19463 ? top_9_8_out :
  32'd0;
assign pe_9_8_left =
  _guard19476 ? left_9_8_out :
  32'd0;
assign pe_9_8_reset = reset;
assign pe_9_8_go = _guard19489;
assign pe_10_3_mul_ready =
  _guard19492 ? 1'd1 :
  _guard19495 ? 1'd0 :
  1'd0;
assign pe_10_3_clk = clk;
assign pe_10_3_top =
  _guard19508 ? top_10_3_out :
  32'd0;
assign pe_10_3_left =
  _guard19521 ? left_10_3_out :
  32'd0;
assign pe_10_3_reset = reset;
assign pe_10_3_go = _guard19534;
assign left_10_5_write_en = _guard19537;
assign left_10_5_clk = clk;
assign left_10_5_reset = reset;
assign left_10_5_in = left_10_4_out;
assign top_10_9_write_en = _guard19543;
assign top_10_9_clk = clk;
assign top_10_9_reset = reset;
assign top_10_9_in = top_9_9_out;
assign top_11_7_write_en = _guard19549;
assign top_11_7_clk = clk;
assign top_11_7_reset = reset;
assign top_11_7_in = top_10_7_out;
assign left_13_3_write_en = _guard19555;
assign left_13_3_clk = clk;
assign left_13_3_reset = reset;
assign left_13_3_in = left_13_2_out;
assign top_13_6_write_en = _guard19561;
assign top_13_6_clk = clk;
assign top_13_6_reset = reset;
assign top_13_6_in = top_12_6_out;
assign left_14_4_write_en = _guard19567;
assign left_14_4_clk = clk;
assign left_14_4_reset = reset;
assign left_14_4_in = left_14_3_out;
assign left_14_9_write_en = _guard19573;
assign left_14_9_clk = clk;
assign left_14_9_reset = reset;
assign left_14_9_in = left_14_8_out;
assign t1_add_left = 5'd1;
assign t1_add_right = t1_idx_out;
assign t3_idx_write_en = _guard19589;
assign t3_idx_clk = clk;
assign t3_idx_reset = reset;
assign t3_idx_in =
  _guard19592 ? t3_add_out :
  _guard19595 ? 5'd0 :
  'x;
assign t12_add_left = 5'd1;
assign t12_add_right = t12_idx_out;
assign l4_add_left = 5'd1;
assign l4_add_right = l4_idx_out;
assign index_ge_16_left = idx_add_out;
assign index_ge_16_right = 6'd16;
assign index_ge_44_left = idx_add_out;
assign index_ge_44_right = 6'd44;
assign index_ge_22_left = idx_add_out;
assign index_ge_22_right = 6'd22;
assign idx_between_13_17_reg_write_en = _guard19618;
assign idx_between_13_17_reg_clk = clk;
assign idx_between_13_17_reg_reset = reset;
assign idx_between_13_17_reg_in =
  _guard19619 ? idx_between_13_17_comb_out :
  _guard19622 ? 1'd0 :
  'x;
assign idx_between_27_43_reg_write_en = _guard19627;
assign idx_between_27_43_reg_clk = clk;
assign idx_between_27_43_reg_reset = reset;
assign idx_between_27_43_reg_in =
  _guard19628 ? idx_between_27_43_comb_out :
  _guard19631 ? 1'd0 :
  'x;
assign idx_between_41_42_reg_write_en = _guard19636;
assign idx_between_41_42_reg_clk = clk;
assign idx_between_41_42_reg_reset = reset;
assign idx_between_41_42_reg_in =
  _guard19637 ? idx_between_41_42_comb_out :
  _guard19640 ? 1'd0 :
  'x;
assign idx_between_47_48_reg_write_en = _guard19645;
assign idx_between_47_48_reg_clk = clk;
assign idx_between_47_48_reg_reset = reset;
assign idx_between_47_48_reg_in =
  _guard19648 ? 1'd0 :
  _guard19649 ? idx_between_47_48_comb_out :
  'x;
assign idx_between_47_48_comb_left = index_ge_47_out;
assign idx_between_47_48_comb_right = index_lt_48_out;
assign idx_between_33_49_comb_left = index_ge_33_out;
assign idx_between_33_49_comb_right = index_lt_49_out;
assign index_ge_48_left = idx_add_out;
assign index_ge_48_right = 6'd48;
assign idx_between_22_23_comb_left = index_ge_22_out;
assign idx_between_22_23_comb_right = index_lt_23_out;
assign idx_between_49_50_reg_write_en = _guard19662;
assign idx_between_49_50_reg_clk = clk;
assign idx_between_49_50_reg_reset = reset;
assign idx_between_49_50_reg_in =
  _guard19663 ? idx_between_49_50_comb_out :
  _guard19666 ? 1'd0 :
  'x;
assign idx_between_4_20_comb_left = index_ge_4_out;
assign idx_between_4_20_comb_right = index_lt_20_out;
assign index_lt_22_left = idx_add_out;
assign index_lt_22_right = 6'd22;
assign index_ge_2_left = idx_add_out;
assign index_ge_2_right = 6'd2;
assign index_ge_19_left = idx_add_out;
assign index_ge_19_right = 6'd19;
assign index_lt_10_left = idx_add_out;
assign index_lt_10_right = 6'd10;
assign idx_between_35_36_reg_write_en = _guard19681;
assign idx_between_35_36_reg_clk = clk;
assign idx_between_35_36_reg_reset = reset;
assign idx_between_35_36_reg_in =
  _guard19684 ? 1'd0 :
  _guard19685 ? idx_between_35_36_comb_out :
  'x;
assign idx_between_12_16_reg_write_en = _guard19690;
assign idx_between_12_16_reg_clk = clk;
assign idx_between_12_16_reg_reset = reset;
assign idx_between_12_16_reg_in =
  _guard19691 ? idx_between_12_16_comb_out :
  _guard19694 ? 1'd0 :
  'x;
assign idx_between_26_42_reg_write_en = _guard19699;
assign idx_between_26_42_reg_clk = clk;
assign idx_between_26_42_reg_reset = reset;
assign idx_between_26_42_reg_in =
  _guard19700 ? idx_between_26_42_comb_out :
  _guard19703 ? 1'd0 :
  'x;
assign idx_between_43_44_comb_left = index_ge_43_out;
assign idx_between_43_44_comb_right = index_lt_44_out;
assign cond_wire_in =
  _guard19708 ? cond_out :
  _guard19709 ? idx_between_0_16_reg_out :
  1'd0;
assign cond_wire15_in =
  _guard19712 ? cond15_out :
  _guard19713 ? idx_between_4_8_reg_out :
  1'd0;
assign cond16_write_en = _guard19714;
assign cond16_clk = clk;
assign cond16_reset = reset;
assign cond16_in =
  _guard19715 ? idx_between_4_20_reg_out :
  1'd0;
assign cond37_write_en = _guard19716;
assign cond37_clk = clk;
assign cond37_reset = reset;
assign cond37_in =
  _guard19717 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire49_in =
  _guard19718 ? idx_between_10_26_reg_out :
  _guard19721 ? cond49_out :
  1'd0;
assign cond_wire55_in =
  _guard19722 ? idx_between_12_16_reg_out :
  _guard19725 ? cond55_out :
  1'd0;
assign cond_wire93_in =
  _guard19726 ? idx_between_5_21_reg_out :
  _guard19729 ? cond93_out :
  1'd0;
assign cond_wire95_in =
  _guard19730 ? idx_between_25_26_reg_out :
  _guard19733 ? cond95_out :
  1'd0;
assign cond_wire96_in =
  _guard19734 ? idx_between_6_10_reg_out :
  _guard19737 ? cond96_out :
  1'd0;
assign cond_wire99_in =
  _guard19738 ? idx_between_26_27_reg_out :
  _guard19741 ? cond99_out :
  1'd0;
assign cond110_write_en = _guard19742;
assign cond110_clk = clk;
assign cond110_reset = reset;
assign cond110_in =
  _guard19743 ? idx_between_13_29_reg_out :
  1'd0;
assign cond113_write_en = _guard19744;
assign cond113_clk = clk;
assign cond113_reset = reset;
assign cond113_in =
  _guard19745 ? idx_between_10_26_reg_out :
  1'd0;
assign cond_wire113_in =
  _guard19748 ? cond113_out :
  _guard19749 ? idx_between_10_26_reg_out :
  1'd0;
assign cond_wire114_in =
  _guard19752 ? cond114_out :
  _guard19753 ? idx_between_14_30_reg_out :
  1'd0;
assign cond125_write_en = _guard19754;
assign cond125_clk = clk;
assign cond125_reset = reset;
assign cond125_in =
  _guard19755 ? idx_between_13_29_reg_out :
  1'd0;
assign cond130_write_en = _guard19756;
assign cond130_clk = clk;
assign cond130_reset = reset;
assign cond130_in =
  _guard19757 ? idx_between_18_34_reg_out :
  1'd0;
assign cond_wire133_in =
  _guard19760 ? cond133_out :
  _guard19761 ? idx_between_15_31_reg_out :
  1'd0;
assign cond144_write_en = _guard19762;
assign cond144_clk = clk;
assign cond144_reset = reset;
assign cond144_in =
  _guard19763 ? idx_between_2_18_reg_out :
  1'd0;
assign cond_wire155_in =
  _guard19766 ? cond155_out :
  _guard19767 ? idx_between_9_25_reg_out :
  1'd0;
assign cond160_write_en = _guard19768;
assign cond160_clk = clk;
assign cond160_reset = reset;
assign cond160_in =
  _guard19769 ? idx_between_26_27_reg_out :
  1'd0;
assign cond163_write_en = _guard19770;
assign cond163_clk = clk;
assign cond163_reset = reset;
assign cond163_in =
  _guard19771 ? idx_between_11_27_reg_out :
  1'd0;
assign cond165_write_en = _guard19772;
assign cond165_clk = clk;
assign cond165_reset = reset;
assign cond165_in =
  _guard19773 ? idx_between_8_12_reg_out :
  1'd0;
assign cond168_write_en = _guard19774;
assign cond168_clk = clk;
assign cond168_reset = reset;
assign cond168_in =
  _guard19775 ? idx_between_28_29_reg_out :
  1'd0;
assign cond_wire173_in =
  _guard19778 ? cond173_out :
  _guard19779 ? idx_between_10_14_reg_out :
  1'd0;
assign cond_wire179_in =
  _guard19782 ? cond179_out :
  _guard19783 ? idx_between_15_31_reg_out :
  1'd0;
assign cond184_write_en = _guard19784;
assign cond184_clk = clk;
assign cond184_reset = reset;
assign cond184_in =
  _guard19785 ? idx_between_32_33_reg_out :
  1'd0;
assign cond185_write_en = _guard19786;
assign cond185_clk = clk;
assign cond185_reset = reset;
assign cond185_in =
  _guard19787 ? idx_between_13_17_reg_out :
  1'd0;
assign cond195_write_en = _guard19788;
assign cond195_clk = clk;
assign cond195_reset = reset;
assign cond195_in =
  _guard19789 ? idx_between_19_35_reg_out :
  1'd0;
assign cond197_write_en = _guard19790;
assign cond197_clk = clk;
assign cond197_reset = reset;
assign cond197_in =
  _guard19791 ? idx_between_16_20_reg_out :
  1'd0;
assign cond207_write_en = _guard19792;
assign cond207_clk = clk;
assign cond207_reset = reset;
assign cond207_in =
  _guard19793 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire217_in =
  _guard19794 ? idx_between_25_26_reg_out :
  _guard19797 ? cond217_out :
  1'd0;
assign cond_wire219_in =
  _guard19798 ? idx_between_6_22_reg_out :
  _guard19801 ? cond219_out :
  1'd0;
assign cond_wire241_in =
  _guard19804 ? cond241_out :
  _guard19805 ? idx_between_31_32_reg_out :
  1'd0;
assign cond243_write_en = _guard19806;
assign cond243_clk = clk;
assign cond243_reset = reset;
assign cond243_in =
  _guard19807 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire244_in =
  _guard19808 ? idx_between_16_32_reg_out :
  _guard19811 ? cond244_out :
  1'd0;
assign cond267_write_en = _guard19812;
assign cond267_clk = clk;
assign cond267_reset = reset;
assign cond267_in =
  _guard19813 ? idx_between_18_34_reg_out :
  1'd0;
assign cond_wire271_in =
  _guard19816 ? cond271_out :
  _guard19817 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire275_in =
  _guard19818 ? idx_between_5_9_reg_out :
  _guard19821 ? cond275_out :
  1'd0;
assign cond278_write_en = _guard19822;
assign cond278_clk = clk;
assign cond278_reset = reset;
assign cond278_in =
  _guard19823 ? idx_between_25_26_reg_out :
  1'd0;
assign cond294_write_en = _guard19824;
assign cond294_clk = clk;
assign cond294_reset = reset;
assign cond294_in =
  _guard19825 ? idx_between_29_30_reg_out :
  1'd0;
assign cond296_write_en = _guard19826;
assign cond296_clk = clk;
assign cond296_reset = reset;
assign cond296_in =
  _guard19827 ? idx_between_10_26_reg_out :
  1'd0;
assign cond299_write_en = _guard19828;
assign cond299_clk = clk;
assign cond299_reset = reset;
assign cond299_in =
  _guard19829 ? idx_between_11_15_reg_out :
  1'd0;
assign cond_wire307_in =
  _guard19832 ? cond307_out :
  _guard19833 ? idx_between_13_17_reg_out :
  1'd0;
assign cond_wire313_in =
  _guard19836 ? cond313_out :
  _guard19837 ? idx_between_18_34_reg_out :
  1'd0;
assign cond318_write_en = _guard19838;
assign cond318_clk = clk;
assign cond318_reset = reset;
assign cond318_in =
  _guard19839 ? idx_between_35_36_reg_out :
  1'd0;
assign cond_wire343_in =
  _guard19840 ? idx_between_26_27_reg_out :
  _guard19843 ? cond343_out :
  1'd0;
assign cond_wire359_in =
  _guard19844 ? idx_between_30_31_reg_out :
  _guard19847 ? cond359_out :
  1'd0;
assign cond374_write_en = _guard19848;
assign cond374_clk = clk;
assign cond374_reset = reset;
assign cond374_in =
  _guard19849 ? idx_between_18_34_reg_out :
  1'd0;
assign cond_wire378_in =
  _guard19852 ? cond378_out :
  _guard19853 ? idx_between_19_35_reg_out :
  1'd0;
assign cond389_write_en = _guard19854;
assign cond389_clk = clk;
assign cond389_reset = reset;
assign cond389_in =
  _guard19855 ? idx_between_18_34_reg_out :
  1'd0;
assign cond_wire391_in =
  _guard19858 ? cond391_out :
  _guard19859 ? idx_between_38_39_reg_out :
  1'd0;
assign cond_wire392_in =
  _guard19860 ? idx_between_19_23_reg_out :
  _guard19863 ? cond392_out :
  1'd0;
assign cond398_write_en = _guard19864;
assign cond398_clk = clk;
assign cond398_reset = reset;
assign cond398_in =
  _guard19865 ? idx_between_24_40_reg_out :
  1'd0;
assign cond417_write_en = _guard19866;
assign cond417_clk = clk;
assign cond417_reset = reset;
assign cond417_in =
  _guard19867 ? idx_between_10_14_reg_out :
  1'd0;
assign cond425_write_en = _guard19868;
assign cond425_clk = clk;
assign cond425_reset = reset;
assign cond425_in =
  _guard19869 ? idx_between_12_16_reg_out :
  1'd0;
assign cond426_write_en = _guard19870;
assign cond426_clk = clk;
assign cond426_reset = reset;
assign cond426_in =
  _guard19871 ? idx_between_12_28_reg_out :
  1'd0;
assign cond427_write_en = _guard19872;
assign cond427_clk = clk;
assign cond427_reset = reset;
assign cond427_in =
  _guard19873 ? idx_between_16_32_reg_out :
  1'd0;
assign cond437_write_en = _guard19874;
assign cond437_clk = clk;
assign cond437_reset = reset;
assign cond437_in =
  _guard19875 ? idx_between_15_19_reg_out :
  1'd0;
assign cond_wire443_in =
  _guard19878 ? cond443_out :
  _guard19879 ? idx_between_20_36_reg_out :
  1'd0;
assign cond451_write_en = _guard19880;
assign cond451_clk = clk;
assign cond451_reset = reset;
assign cond451_in =
  _guard19881 ? idx_between_22_38_reg_out :
  1'd0;
assign cond468_write_en = _guard19882;
assign cond468_clk = clk;
assign cond468_reset = reset;
assign cond468_in =
  _guard19883 ? idx_between_42_43_reg_out :
  1'd0;
assign cond_wire470_in =
  _guard19884 ? idx_between_8_12_reg_out :
  _guard19887 ? cond470_out :
  1'd0;
assign cond_wire472_in =
  _guard19890 ? cond472_out :
  _guard19891 ? idx_between_12_28_reg_out :
  1'd0;
assign cond477_write_en = _guard19892;
assign cond477_clk = clk;
assign cond477_reset = reset;
assign cond477_in =
  _guard19893 ? idx_between_29_30_reg_out :
  1'd0;
assign cond_wire478_in =
  _guard19896 ? cond478_out :
  _guard19897 ? idx_between_10_14_reg_out :
  1'd0;
assign cond_wire482_in =
  _guard19900 ? cond482_out :
  _guard19901 ? idx_between_11_15_reg_out :
  1'd0;
assign cond_wire504_in =
  _guard19904 ? cond504_out :
  _guard19905 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire514_in =
  _guard19906 ? idx_between_19_23_reg_out :
  _guard19909 ? cond514_out :
  1'd0;
assign cond528_write_en = _guard19910;
assign cond528_clk = clk;
assign cond528_reset = reset;
assign cond528_in =
  _guard19911 ? idx_between_26_42_reg_out :
  1'd0;
assign cond_wire528_in =
  _guard19912 ? idx_between_26_42_reg_out :
  _guard19915 ? cond528_out :
  1'd0;
assign cond530_write_en = _guard19916;
assign cond530_clk = clk;
assign cond530_reset = reset;
assign cond530_in =
  _guard19917 ? idx_between_23_27_reg_out :
  1'd0;
assign cond536_write_en = _guard19918;
assign cond536_clk = clk;
assign cond536_reset = reset;
assign cond536_in =
  _guard19919 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire538_in =
  _guard19922 ? cond538_out :
  _guard19923 ? idx_between_29_30_reg_out :
  1'd0;
assign cond_wire540_in =
  _guard19924 ? idx_between_10_26_reg_out :
  _guard19927 ? cond540_out :
  1'd0;
assign cond550_write_en = _guard19928;
assign cond550_clk = clk;
assign cond550_reset = reset;
assign cond550_in =
  _guard19929 ? idx_between_32_33_reg_out :
  1'd0;
assign cond_wire555_in =
  _guard19930 ? idx_between_14_18_reg_out :
  _guard19933 ? cond555_out :
  1'd0;
assign cond571_write_en = _guard19934;
assign cond571_clk = clk;
assign cond571_reset = reset;
assign cond571_in =
  _guard19935 ? idx_between_18_22_reg_out :
  1'd0;
assign cond573_write_en = _guard19936;
assign cond573_clk = clk;
assign cond573_reset = reset;
assign cond573_in =
  _guard19937 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire593_in =
  _guard19938 ? idx_between_27_43_reg_out :
  _guard19941 ? cond593_out :
  1'd0;
assign cond_wire595_in =
  _guard19942 ? idx_between_24_28_reg_out :
  _guard19945 ? cond595_out :
  1'd0;
assign cond609_write_en = _guard19946;
assign cond609_clk = clk;
assign cond609_reset = reset;
assign cond609_in =
  _guard19947 ? idx_between_12_28_reg_out :
  1'd0;
assign cond613_write_en = _guard19948;
assign cond613_clk = clk;
assign cond613_reset = reset;
assign cond613_in =
  _guard19949 ? idx_between_13_29_reg_out :
  1'd0;
assign cond_wire619_in =
  _guard19950 ? idx_between_34_35_reg_out :
  _guard19953 ? cond619_out :
  1'd0;
assign cond627_write_en = _guard19954;
assign cond627_clk = clk;
assign cond627_reset = reset;
assign cond627_in =
  _guard19955 ? idx_between_36_37_reg_out :
  1'd0;
assign cond_wire627_in =
  _guard19956 ? idx_between_36_37_reg_out :
  _guard19959 ? cond627_out :
  1'd0;
assign cond_wire631_in =
  _guard19962 ? cond631_out :
  _guard19963 ? idx_between_37_38_reg_out :
  1'd0;
assign cond632_write_en = _guard19964;
assign cond632_clk = clk;
assign cond632_reset = reset;
assign cond632_in =
  _guard19965 ? idx_between_18_22_reg_out :
  1'd0;
assign cond_wire651_in =
  _guard19966 ? idx_between_42_43_reg_out :
  _guard19969 ? cond651_out :
  1'd0;
assign cond_wire673_in =
  _guard19970 ? idx_between_13_17_reg_out :
  _guard19973 ? cond673_out :
  1'd0;
assign cond678_write_en = _guard19974;
assign cond678_clk = clk;
assign cond678_reset = reset;
assign cond678_in =
  _guard19975 ? idx_between_14_30_reg_out :
  1'd0;
assign cond680_write_en = _guard19976;
assign cond680_clk = clk;
assign cond680_reset = reset;
assign cond680_in =
  _guard19977 ? idx_between_34_35_reg_out :
  1'd0;
assign cond_wire686_in =
  _guard19978 ? idx_between_16_32_reg_out :
  _guard19981 ? cond686_out :
  1'd0;
assign cond689_write_en = _guard19982;
assign cond689_clk = clk;
assign cond689_reset = reset;
assign cond689_in =
  _guard19983 ? idx_between_17_21_reg_out :
  1'd0;
assign cond_wire705_in =
  _guard19984 ? idx_between_21_25_reg_out :
  _guard19987 ? cond705_out :
  1'd0;
assign cond_wire716_in =
  _guard19988 ? idx_between_43_44_reg_out :
  _guard19991 ? cond716_out :
  1'd0;
assign cond726_write_en = _guard19992;
assign cond726_clk = clk;
assign cond726_reset = reset;
assign cond726_in =
  _guard19993 ? idx_between_26_42_reg_out :
  1'd0;
assign cond733_write_en = _guard19994;
assign cond733_clk = clk;
assign cond733_reset = reset;
assign cond733_in =
  _guard19995 ? idx_between_32_33_reg_out :
  1'd0;
assign cond735_write_en = _guard19996;
assign cond735_clk = clk;
assign cond735_reset = reset;
assign cond735_in =
  _guard19997 ? idx_between_13_29_reg_out :
  1'd0;
assign cond737_write_en = _guard19998;
assign cond737_clk = clk;
assign cond737_reset = reset;
assign cond737_in =
  _guard19999 ? idx_between_33_34_reg_out :
  1'd0;
assign cond_wire737_in =
  _guard20002 ? cond737_out :
  _guard20003 ? idx_between_33_34_reg_out :
  1'd0;
assign cond741_write_en = _guard20004;
assign cond741_clk = clk;
assign cond741_reset = reset;
assign cond741_in =
  _guard20005 ? idx_between_34_35_reg_out :
  1'd0;
assign cond_wire758_in =
  _guard20006 ? idx_between_19_23_reg_out :
  _guard20009 ? cond758_out :
  1'd0;
assign cond768_write_en = _guard20010;
assign cond768_clk = clk;
assign cond768_reset = reset;
assign cond768_in =
  _guard20011 ? idx_between_25_41_reg_out :
  1'd0;
assign cond805_write_en = _guard20012;
assign cond805_clk = clk;
assign cond805_reset = reset;
assign cond805_in =
  _guard20013 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire819_in =
  _guard20014 ? idx_between_19_23_reg_out :
  _guard20017 ? cond819_out :
  1'd0;
assign cond824_write_en = _guard20018;
assign cond824_clk = clk;
assign cond824_reset = reset;
assign cond824_in =
  _guard20019 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire825_in =
  _guard20020 ? idx_between_24_40_reg_out :
  _guard20023 ? cond825_out :
  1'd0;
assign cond826_write_en = _guard20024;
assign cond826_clk = clk;
assign cond826_reset = reset;
assign cond826_in =
  _guard20025 ? idx_between_40_41_reg_out :
  1'd0;
assign cond831_write_en = _guard20026;
assign cond831_clk = clk;
assign cond831_reset = reset;
assign cond831_in =
  _guard20027 ? idx_between_22_26_reg_out :
  1'd0;
assign cond_wire841_in =
  _guard20030 ? cond841_out :
  _guard20031 ? idx_between_28_44_reg_out :
  1'd0;
assign cond846_write_en = _guard20032;
assign cond846_clk = clk;
assign cond846_reset = reset;
assign cond846_in =
  _guard20033 ? idx_between_45_46_reg_out :
  1'd0;
assign cond_wire846_in =
  _guard20036 ? cond846_out :
  _guard20037 ? idx_between_45_46_reg_out :
  1'd0;
assign cond856_write_en = _guard20038;
assign cond856_clk = clk;
assign cond856_reset = reset;
assign cond856_in =
  _guard20039 ? idx_between_28_44_reg_out :
  1'd0;
assign cond_wire867_in =
  _guard20042 ? cond867_out :
  _guard20043 ? idx_between_35_36_reg_out :
  1'd0;
assign cond_wire873_in =
  _guard20044 ? idx_between_17_33_reg_out :
  _guard20047 ? cond873_out :
  1'd0;
assign cond879_write_en = _guard20048;
assign cond879_clk = clk;
assign cond879_reset = reset;
assign cond879_in =
  _guard20049 ? idx_between_38_39_reg_out :
  1'd0;
assign cond_wire896_in =
  _guard20052 ? cond896_out :
  _guard20053 ? idx_between_23_27_reg_out :
  1'd0;
assign cond898_write_en = _guard20054;
assign cond898_clk = clk;
assign cond898_reset = reset;
assign cond898_in =
  _guard20055 ? idx_between_27_43_reg_out :
  1'd0;
assign cond_wire898_in =
  _guard20056 ? idx_between_27_43_reg_out :
  _guard20059 ? cond898_out :
  1'd0;
assign cond902_write_en = _guard20060;
assign cond902_clk = clk;
assign cond902_reset = reset;
assign cond902_in =
  _guard20061 ? idx_between_28_44_reg_out :
  1'd0;
assign cond911_write_en = _guard20062;
assign cond911_clk = clk;
assign cond911_reset = reset;
assign cond911_in =
  _guard20063 ? idx_between_46_47_reg_out :
  1'd0;
assign cond_wire911_in =
  _guard20066 ? cond911_out :
  _guard20067 ? idx_between_46_47_reg_out :
  1'd0;
assign cond913_write_en = _guard20068;
assign cond913_clk = clk;
assign cond913_reset = reset;
assign cond913_in =
  _guard20069 ? idx_between_27_43_reg_out :
  1'd0;
assign cond952_write_en = _guard20070;
assign cond952_clk = clk;
assign cond952_reset = reset;
assign cond952_in =
  _guard20071 ? idx_between_41_42_reg_out :
  1'd0;
assign cond_wire960_in =
  _guard20072 ? idx_between_43_44_reg_out :
  _guard20075 ? cond960_out :
  1'd0;
assign cond963_write_en = _guard20076;
assign cond963_clk = clk;
assign cond963_reset = reset;
assign cond963_in =
  _guard20077 ? idx_between_28_44_reg_out :
  1'd0;
assign cond_wire973_in =
  _guard20080 ? cond973_out :
  _guard20081 ? idx_between_27_31_reg_out :
  1'd0;
assign cond975_write_en = _guard20082;
assign cond975_clk = clk;
assign cond975_reset = reset;
assign cond975_in =
  _guard20083 ? idx_between_31_47_reg_out :
  1'd0;
assign cond989_write_en = _guard20084;
assign cond989_clk = clk;
assign cond989_reset = reset;
assign cond989_in =
  _guard20085 ? idx_between_15_31_reg_out :
  1'd0;
assign cond995_write_en = _guard20086;
assign cond995_clk = clk;
assign cond995_reset = reset;
assign cond995_in =
  _guard20087 ? idx_between_17_33_reg_out :
  1'd0;
assign cond_wire1005_in =
  _guard20090 ? cond1005_out :
  _guard20091 ? idx_between_39_40_reg_out :
  1'd0;
assign cond_wire1009_in =
  _guard20094 ? cond1009_out :
  _guard20095 ? idx_between_40_41_reg_out :
  1'd0;
assign cond1042_write_en = _guard20096;
assign cond1042_clk = clk;
assign cond1042_reset = reset;
assign cond1042_in =
  _guard20097 ? idx_between_29_33_reg_out :
  1'd0;
assign cond1043_write_en = _guard20098;
assign cond1043_clk = clk;
assign cond1043_reset = reset;
assign cond1043_in =
  _guard20099 ? idx_between_29_45_reg_out :
  1'd0;
assign pe_0_0_mul_ready =
  _guard20102 ? 1'd1 :
  _guard20105 ? 1'd0 :
  1'd0;
assign pe_0_0_clk = clk;
assign pe_0_0_top =
  _guard20118 ? top_0_0_out :
  32'd0;
assign pe_0_0_left =
  _guard20131 ? left_0_0_out :
  32'd0;
assign pe_0_0_reset = reset;
assign pe_0_0_go = _guard20144;
assign left_0_13_write_en = _guard20147;
assign left_0_13_clk = clk;
assign left_0_13_reset = reset;
assign left_0_13_in = left_0_12_out;
assign left_1_6_write_en = _guard20153;
assign left_1_6_clk = clk;
assign left_1_6_reset = reset;
assign left_1_6_in = left_1_5_out;
assign left_1_8_write_en = _guard20159;
assign left_1_8_clk = clk;
assign left_1_8_reset = reset;
assign left_1_8_in = left_1_7_out;
assign top_1_14_write_en = _guard20165;
assign top_1_14_clk = clk;
assign top_1_14_reset = reset;
assign top_1_14_in = top_0_14_out;
assign top_2_8_write_en = _guard20171;
assign top_2_8_clk = clk;
assign top_2_8_reset = reset;
assign top_2_8_in = top_1_8_out;
assign left_2_10_write_en = _guard20177;
assign left_2_10_clk = clk;
assign left_2_10_reset = reset;
assign left_2_10_in = left_2_9_out;
assign pe_3_3_mul_ready =
  _guard20183 ? 1'd1 :
  _guard20186 ? 1'd0 :
  1'd0;
assign pe_3_3_clk = clk;
assign pe_3_3_top =
  _guard20199 ? top_3_3_out :
  32'd0;
assign pe_3_3_left =
  _guard20212 ? left_3_3_out :
  32'd0;
assign pe_3_3_reset = reset;
assign pe_3_3_go = _guard20225;
assign top_3_3_write_en = _guard20228;
assign top_3_3_clk = clk;
assign top_3_3_reset = reset;
assign top_3_3_in = top_2_3_out;
assign left_3_10_write_en = _guard20234;
assign left_3_10_clk = clk;
assign left_3_10_reset = reset;
assign left_3_10_in = left_3_9_out;
assign left_3_14_write_en = _guard20240;
assign left_3_14_clk = clk;
assign left_3_14_reset = reset;
assign left_3_14_in = left_3_13_out;
assign top_4_3_write_en = _guard20246;
assign top_4_3_clk = clk;
assign top_4_3_reset = reset;
assign top_4_3_in = top_3_3_out;
assign top_4_6_write_en = _guard20252;
assign top_4_6_clk = clk;
assign top_4_6_reset = reset;
assign top_4_6_in = top_3_6_out;
assign pe_5_6_mul_ready =
  _guard20258 ? 1'd1 :
  _guard20261 ? 1'd0 :
  1'd0;
assign pe_5_6_clk = clk;
assign pe_5_6_top =
  _guard20274 ? top_5_6_out :
  32'd0;
assign pe_5_6_left =
  _guard20287 ? left_5_6_out :
  32'd0;
assign pe_5_6_reset = reset;
assign pe_5_6_go = _guard20300;
assign top_5_6_write_en = _guard20303;
assign top_5_6_clk = clk;
assign top_5_6_reset = reset;
assign top_5_6_in = top_4_6_out;
assign top_6_2_write_en = _guard20309;
assign top_6_2_clk = clk;
assign top_6_2_reset = reset;
assign top_6_2_in = top_5_2_out;
assign left_6_9_write_en = _guard20315;
assign left_6_9_clk = clk;
assign left_6_9_reset = reset;
assign left_6_9_in = left_6_8_out;
assign top_6_15_write_en = _guard20321;
assign top_6_15_clk = clk;
assign top_6_15_reset = reset;
assign top_6_15_in = top_5_15_out;
assign pe_7_1_mul_ready =
  _guard20327 ? 1'd1 :
  _guard20330 ? 1'd0 :
  1'd0;
assign pe_7_1_clk = clk;
assign pe_7_1_top =
  _guard20343 ? top_7_1_out :
  32'd0;
assign pe_7_1_left =
  _guard20356 ? left_7_1_out :
  32'd0;
assign pe_7_1_reset = reset;
assign pe_7_1_go = _guard20369;
assign pe_7_12_mul_ready =
  _guard20372 ? 1'd1 :
  _guard20375 ? 1'd0 :
  1'd0;
assign pe_7_12_clk = clk;
assign pe_7_12_top =
  _guard20388 ? top_7_12_out :
  32'd0;
assign pe_7_12_left =
  _guard20401 ? left_7_12_out :
  32'd0;
assign pe_7_12_reset = reset;
assign pe_7_12_go = _guard20414;
assign left_7_13_write_en = _guard20417;
assign left_7_13_clk = clk;
assign left_7_13_reset = reset;
assign left_7_13_in = left_7_12_out;
assign pe_8_3_mul_ready =
  _guard20423 ? 1'd1 :
  _guard20426 ? 1'd0 :
  1'd0;
assign pe_8_3_clk = clk;
assign pe_8_3_top =
  _guard20439 ? top_8_3_out :
  32'd0;
assign pe_8_3_left =
  _guard20452 ? left_8_3_out :
  32'd0;
assign pe_8_3_reset = reset;
assign pe_8_3_go = _guard20465;
assign pe_8_12_mul_ready =
  _guard20468 ? 1'd1 :
  _guard20471 ? 1'd0 :
  1'd0;
assign pe_8_12_clk = clk;
assign pe_8_12_top =
  _guard20484 ? top_8_12_out :
  32'd0;
assign pe_8_12_left =
  _guard20497 ? left_8_12_out :
  32'd0;
assign pe_8_12_reset = reset;
assign pe_8_12_go = _guard20510;
assign left_9_0_write_en = _guard20513;
assign left_9_0_clk = clk;
assign left_9_0_reset = reset;
assign left_9_0_in = l9_read_data;
assign top_9_11_write_en = _guard20519;
assign top_9_11_clk = clk;
assign top_9_11_reset = reset;
assign top_9_11_in = top_8_11_out;
assign left_9_12_write_en = _guard20525;
assign left_9_12_clk = clk;
assign left_9_12_reset = reset;
assign left_9_12_in = left_9_11_out;
assign pe_9_14_mul_ready =
  _guard20531 ? 1'd1 :
  _guard20534 ? 1'd0 :
  1'd0;
assign pe_9_14_clk = clk;
assign pe_9_14_top =
  _guard20547 ? top_9_14_out :
  32'd0;
assign pe_9_14_left =
  _guard20560 ? left_9_14_out :
  32'd0;
assign pe_9_14_reset = reset;
assign pe_9_14_go = _guard20573;
assign left_10_2_write_en = _guard20576;
assign left_10_2_clk = clk;
assign left_10_2_reset = reset;
assign left_10_2_in = left_10_1_out;
assign pe_10_4_mul_ready =
  _guard20582 ? 1'd1 :
  _guard20585 ? 1'd0 :
  1'd0;
assign pe_10_4_clk = clk;
assign pe_10_4_top =
  _guard20598 ? top_10_4_out :
  32'd0;
assign pe_10_4_left =
  _guard20611 ? left_10_4_out :
  32'd0;
assign pe_10_4_reset = reset;
assign pe_10_4_go = _guard20624;
assign top_10_4_write_en = _guard20627;
assign top_10_4_clk = clk;
assign top_10_4_reset = reset;
assign top_10_4_in = top_9_4_out;
assign pe_10_15_mul_ready =
  _guard20633 ? 1'd1 :
  _guard20636 ? 1'd0 :
  1'd0;
assign pe_10_15_clk = clk;
assign pe_10_15_top =
  _guard20649 ? top_10_15_out :
  32'd0;
assign pe_10_15_left =
  _guard20662 ? left_10_15_out :
  32'd0;
assign pe_10_15_reset = reset;
assign pe_10_15_go = _guard20675;
assign top_10_15_write_en = _guard20678;
assign top_10_15_clk = clk;
assign top_10_15_reset = reset;
assign top_10_15_in = top_9_15_out;
assign top_11_4_write_en = _guard20684;
assign top_11_4_clk = clk;
assign top_11_4_reset = reset;
assign top_11_4_in = top_10_4_out;
assign left_11_6_write_en = _guard20690;
assign left_11_6_clk = clk;
assign left_11_6_reset = reset;
assign left_11_6_in = left_11_5_out;
assign top_11_9_write_en = _guard20696;
assign top_11_9_clk = clk;
assign top_11_9_reset = reset;
assign top_11_9_in = top_10_9_out;
assign top_11_10_write_en = _guard20702;
assign top_11_10_clk = clk;
assign top_11_10_reset = reset;
assign top_11_10_in = top_10_10_out;
assign pe_11_13_mul_ready =
  _guard20708 ? 1'd1 :
  _guard20711 ? 1'd0 :
  1'd0;
assign pe_11_13_clk = clk;
assign pe_11_13_top =
  _guard20724 ? top_11_13_out :
  32'd0;
assign pe_11_13_left =
  _guard20737 ? left_11_13_out :
  32'd0;
assign pe_11_13_reset = reset;
assign pe_11_13_go = _guard20750;
assign pe_11_14_mul_ready =
  _guard20753 ? 1'd1 :
  _guard20756 ? 1'd0 :
  1'd0;
assign pe_11_14_clk = clk;
assign pe_11_14_top =
  _guard20769 ? top_11_14_out :
  32'd0;
assign pe_11_14_left =
  _guard20782 ? left_11_14_out :
  32'd0;
assign pe_11_14_reset = reset;
assign pe_11_14_go = _guard20795;
assign left_12_2_write_en = _guard20798;
assign left_12_2_clk = clk;
assign left_12_2_reset = reset;
assign left_12_2_in = left_12_1_out;
assign pe_12_5_mul_ready =
  _guard20804 ? 1'd1 :
  _guard20807 ? 1'd0 :
  1'd0;
assign pe_12_5_clk = clk;
assign pe_12_5_top =
  _guard20820 ? top_12_5_out :
  32'd0;
assign pe_12_5_left =
  _guard20833 ? left_12_5_out :
  32'd0;
assign pe_12_5_reset = reset;
assign pe_12_5_go = _guard20846;
assign left_12_6_write_en = _guard20849;
assign left_12_6_clk = clk;
assign left_12_6_reset = reset;
assign left_12_6_in = left_12_5_out;
assign left_12_7_write_en = _guard20855;
assign left_12_7_clk = clk;
assign left_12_7_reset = reset;
assign left_12_7_in = left_12_6_out;
assign pe_12_13_mul_ready =
  _guard20861 ? 1'd1 :
  _guard20864 ? 1'd0 :
  1'd0;
assign pe_12_13_clk = clk;
assign pe_12_13_top =
  _guard20877 ? top_12_13_out :
  32'd0;
assign pe_12_13_left =
  _guard20890 ? left_12_13_out :
  32'd0;
assign pe_12_13_reset = reset;
assign pe_12_13_go = _guard20903;
assign pe_12_15_mul_ready =
  _guard20906 ? 1'd1 :
  _guard20909 ? 1'd0 :
  1'd0;
assign pe_12_15_clk = clk;
assign pe_12_15_top =
  _guard20922 ? top_12_15_out :
  32'd0;
assign pe_12_15_left =
  _guard20935 ? left_12_15_out :
  32'd0;
assign pe_12_15_reset = reset;
assign pe_12_15_go = _guard20948;
assign top_12_15_write_en = _guard20951;
assign top_12_15_clk = clk;
assign top_12_15_reset = reset;
assign top_12_15_in = top_11_15_out;
assign left_13_4_write_en = _guard20957;
assign left_13_4_clk = clk;
assign left_13_4_reset = reset;
assign left_13_4_in = left_13_3_out;
assign pe_13_9_mul_ready =
  _guard20963 ? 1'd1 :
  _guard20966 ? 1'd0 :
  1'd0;
assign pe_13_9_clk = clk;
assign pe_13_9_top =
  _guard20979 ? top_13_9_out :
  32'd0;
assign pe_13_9_left =
  _guard20992 ? left_13_9_out :
  32'd0;
assign pe_13_9_reset = reset;
assign pe_13_9_go = _guard21005;
assign pe_14_3_mul_ready =
  _guard21008 ? 1'd1 :
  _guard21011 ? 1'd0 :
  1'd0;
assign pe_14_3_clk = clk;
assign pe_14_3_top =
  _guard21024 ? top_14_3_out :
  32'd0;
assign pe_14_3_left =
  _guard21037 ? left_14_3_out :
  32'd0;
assign pe_14_3_reset = reset;
assign pe_14_3_go = _guard21050;
assign top_14_6_write_en = _guard21053;
assign top_14_6_clk = clk;
assign top_14_6_reset = reset;
assign top_14_6_in = top_13_6_out;
assign pe_14_10_mul_ready =
  _guard21059 ? 1'd1 :
  _guard21062 ? 1'd0 :
  1'd0;
assign pe_14_10_clk = clk;
assign pe_14_10_top =
  _guard21075 ? top_14_10_out :
  32'd0;
assign pe_14_10_left =
  _guard21088 ? left_14_10_out :
  32'd0;
assign pe_14_10_reset = reset;
assign pe_14_10_go = _guard21101;
assign left_14_14_write_en = _guard21104;
assign left_14_14_clk = clk;
assign left_14_14_reset = reset;
assign left_14_14_in = left_14_13_out;
assign left_15_1_write_en = _guard21110;
assign left_15_1_clk = clk;
assign left_15_1_reset = reset;
assign left_15_1_in = left_15_0_out;
assign top_15_2_write_en = _guard21116;
assign top_15_2_clk = clk;
assign top_15_2_reset = reset;
assign top_15_2_in = top_14_2_out;
assign pe_15_3_mul_ready =
  _guard21122 ? 1'd1 :
  _guard21125 ? 1'd0 :
  1'd0;
assign pe_15_3_clk = clk;
assign pe_15_3_top =
  _guard21138 ? top_15_3_out :
  32'd0;
assign pe_15_3_left =
  _guard21151 ? left_15_3_out :
  32'd0;
assign pe_15_3_reset = reset;
assign pe_15_3_go = _guard21164;
assign pe_15_6_mul_ready =
  _guard21167 ? 1'd1 :
  _guard21170 ? 1'd0 :
  1'd0;
assign pe_15_6_clk = clk;
assign pe_15_6_top =
  _guard21183 ? top_15_6_out :
  32'd0;
assign pe_15_6_left =
  _guard21196 ? left_15_6_out :
  32'd0;
assign pe_15_6_reset = reset;
assign pe_15_6_go = _guard21209;
assign pe_15_15_mul_ready =
  _guard21212 ? 1'd1 :
  _guard21215 ? 1'd0 :
  1'd0;
assign pe_15_15_clk = clk;
assign pe_15_15_top =
  _guard21228 ? top_15_15_out :
  32'd0;
assign pe_15_15_left =
  _guard21241 ? left_15_15_out :
  32'd0;
assign pe_15_15_reset = reset;
assign pe_15_15_go = _guard21254;
assign t2_add_left = 5'd1;
assign t2_add_right = t2_idx_out;
assign t5_add_left = 5'd1;
assign t5_add_right = t5_idx_out;
assign t9_add_left = 5'd1;
assign t9_add_right = t9_idx_out;
assign t13_idx_write_en = _guard21279;
assign t13_idx_clk = clk;
assign t13_idx_reset = reset;
assign t13_idx_in =
  _guard21282 ? 5'd0 :
  _guard21285 ? t13_add_out :
  'x;
assign l8_add_left = 5'd1;
assign l8_add_right = l8_idx_out;
assign idx_between_44_45_comb_left = index_ge_44_out;
assign idx_between_44_45_comb_right = index_lt_45_out;
assign index_lt_51_left = idx_add_out;
assign index_lt_51_right = 6'd51;
assign idx_between_40_41_comb_left = index_ge_40_out;
assign idx_between_40_41_comb_right = index_lt_41_out;
assign index_ge_5_left = idx_add_out;
assign index_ge_5_right = 6'd5;
assign idx_between_5_21_comb_left = index_ge_5_out;
assign idx_between_5_21_comb_right = index_lt_21_out;
assign idx_between_0_16_reg_write_en = _guard21306;
assign idx_between_0_16_reg_clk = clk;
assign idx_between_0_16_reg_reset = reset;
assign idx_between_0_16_reg_in =
  _guard21309 ? 1'd1 :
  _guard21310 ? index_lt_16_out :
  'x;
assign index_lt_48_left = idx_add_out;
assign index_lt_48_right = 6'd48;
assign idx_between_3_19_comb_left = index_ge_3_out;
assign idx_between_3_19_comb_right = index_lt_19_out;
assign idx_between_45_46_reg_write_en = _guard21319;
assign idx_between_45_46_reg_clk = clk;
assign idx_between_45_46_reg_reset = reset;
assign idx_between_45_46_reg_in =
  _guard21320 ? idx_between_45_46_comb_out :
  _guard21323 ? 1'd0 :
  'x;
assign idx_between_10_26_reg_write_en = _guard21328;
assign idx_between_10_26_reg_clk = clk;
assign idx_between_10_26_reg_reset = reset;
assign idx_between_10_26_reg_in =
  _guard21329 ? idx_between_10_26_comb_out :
  _guard21332 ? 1'd0 :
  'x;
assign index_ge_10_left = idx_add_out;
assign index_ge_10_right = 6'd10;
assign idx_between_7_11_comb_left = index_ge_7_out;
assign idx_between_7_11_comb_right = index_lt_11_out;
assign idx_between_12_28_comb_left = index_ge_12_out;
assign idx_between_12_28_comb_right = index_lt_28_out;
assign idx_between_27_28_comb_left = index_ge_27_out;
assign idx_between_27_28_comb_right = index_lt_28_out;
assign idx_between_19_35_reg_write_en = _guard21345;
assign idx_between_19_35_reg_clk = clk;
assign idx_between_19_35_reg_reset = reset;
assign idx_between_19_35_reg_in =
  _guard21346 ? idx_between_19_35_comb_out :
  _guard21349 ? 1'd0 :
  'x;
assign index_lt_12_left = idx_add_out;
assign index_lt_12_right = 6'd12;
assign idx_between_22_38_reg_write_en = _guard21356;
assign idx_between_22_38_reg_clk = clk;
assign idx_between_22_38_reg_reset = reset;
assign idx_between_22_38_reg_in =
  _guard21357 ? idx_between_22_38_comb_out :
  _guard21360 ? 1'd0 :
  'x;
assign index_lt_38_left = idx_add_out;
assign index_lt_38_right = 6'd38;
assign idx_between_18_22_reg_write_en = _guard21367;
assign idx_between_18_22_reg_clk = clk;
assign idx_between_18_22_reg_reset = reset;
assign idx_between_18_22_reg_in =
  _guard21368 ? idx_between_18_22_comb_out :
  _guard21371 ? 1'd0 :
  'x;
assign idx_between_33_34_reg_write_en = _guard21376;
assign idx_between_33_34_reg_clk = clk;
assign idx_between_33_34_reg_reset = reset;
assign idx_between_33_34_reg_in =
  _guard21377 ? idx_between_33_34_comb_out :
  _guard21380 ? 1'd0 :
  'x;
assign idx_between_24_40_reg_write_en = _guard21385;
assign idx_between_24_40_reg_clk = clk;
assign idx_between_24_40_reg_reset = reset;
assign idx_between_24_40_reg_in =
  _guard21388 ? 1'd0 :
  _guard21389 ? idx_between_24_40_comb_out :
  'x;
assign cond0_write_en = _guard21390;
assign cond0_clk = clk;
assign cond0_reset = reset;
assign cond0_in =
  _guard21391 ? idx_between_1_5_reg_out :
  1'd0;
assign cond_wire7_in =
  _guard21392 ? idx_between_6_22_reg_out :
  _guard21395 ? cond7_out :
  1'd0;
assign cond_wire10_in =
  _guard21396 ? idx_between_3_7_reg_out :
  _guard21399 ? cond10_out :
  1'd0;
assign cond_wire12_in =
  _guard21400 ? idx_between_7_23_reg_out :
  _guard21403 ? cond12_out :
  1'd0;
assign cond_wire17_in =
  _guard21406 ? cond17_out :
  _guard21407 ? idx_between_8_24_reg_out :
  1'd0;
assign cond_wire19_in =
  _guard21410 ? cond19_out :
  _guard21411 ? idx_between_4_20_reg_out :
  1'd0;
assign cond_wire23_in =
  _guard21412 ? idx_between_25_26_reg_out :
  _guard21415 ? cond23_out :
  1'd0;
assign cond_wire25_in =
  _guard21416 ? idx_between_6_10_reg_out :
  _guard21419 ? cond25_out :
  1'd0;
assign cond33_write_en = _guard21420;
assign cond33_clk = clk;
assign cond33_reset = reset;
assign cond33_in =
  _guard21421 ? idx_between_27_28_reg_out :
  1'd0;
assign cond_wire42_in =
  _guard21422 ? idx_between_13_29_reg_out :
  _guard21425 ? cond42_out :
  1'd0;
assign cond47_write_en = _guard21426;
assign cond47_clk = clk;
assign cond47_reset = reset;
assign cond47_in =
  _guard21427 ? idx_between_14_30_reg_out :
  1'd0;
assign cond48_write_en = _guard21428;
assign cond48_clk = clk;
assign cond48_reset = reset;
assign cond48_in =
  _guard21429 ? idx_between_30_31_reg_out :
  1'd0;
assign cond66_write_en = _guard21430;
assign cond66_clk = clk;
assign cond66_reset = reset;
assign cond66_in =
  _guard21431 ? idx_between_14_30_reg_out :
  1'd0;
assign cond_wire69_in =
  _guard21434 ? cond69_out :
  _guard21435 ? idx_between_14_30_reg_out :
  1'd0;
assign cond_wire71_in =
  _guard21438 ? cond71_out :
  _guard21439 ? idx_between_15_31_reg_out :
  1'd0;
assign cond82_write_en = _guard21440;
assign cond82_clk = clk;
assign cond82_reset = reset;
assign cond82_in =
  _guard21441 ? idx_between_6_22_reg_out :
  1'd0;
assign cond84_write_en = _guard21442;
assign cond84_clk = clk;
assign cond84_reset = reset;
assign cond84_in =
  _guard21443 ? idx_between_3_7_reg_out :
  1'd0;
assign cond_wire94_in =
  _guard21446 ? cond94_out :
  _guard21447 ? idx_between_9_25_reg_out :
  1'd0;
assign cond102_write_en = _guard21448;
assign cond102_clk = clk;
assign cond102_reset = reset;
assign cond102_in =
  _guard21449 ? idx_between_11_27_reg_out :
  1'd0;
assign cond_wire104_in =
  _guard21450 ? idx_between_8_12_reg_out :
  _guard21453 ? cond104_out :
  1'd0;
assign cond108_write_en = _guard21454;
assign cond108_clk = clk;
assign cond108_reset = reset;
assign cond108_in =
  _guard21455 ? idx_between_9_13_reg_out :
  1'd0;
assign cond_wire110_in =
  _guard21456 ? idx_between_13_29_reg_out :
  _guard21459 ? cond110_out :
  1'd0;
assign cond119_write_en = _guard21460;
assign cond119_clk = clk;
assign cond119_reset = reset;
assign cond119_in =
  _guard21461 ? idx_between_31_32_reg_out :
  1'd0;
assign cond120_write_en = _guard21462;
assign cond120_clk = clk;
assign cond120_reset = reset;
assign cond120_in =
  _guard21463 ? idx_between_12_16_reg_out :
  1'd0;
assign cond_wire130_in =
  _guard21464 ? idx_between_18_34_reg_out :
  _guard21467 ? cond130_out :
  1'd0;
assign cond_wire135_in =
  _guard21468 ? idx_between_35_36_reg_out :
  _guard21471 ? cond135_out :
  1'd0;
assign cond141_write_en = _guard21472;
assign cond141_clk = clk;
assign cond141_reset = reset;
assign cond141_in =
  _guard21473 ? idx_between_17_33_reg_out :
  1'd0;
assign cond_wire150_in =
  _guard21476 ? cond150_out :
  _guard21477 ? idx_between_4_20_reg_out :
  1'd0;
assign cond_wire152_in =
  _guard21478 ? idx_between_24_25_reg_out :
  _guard21481 ? cond152_out :
  1'd0;
assign cond_wire153_in =
  _guard21482 ? idx_between_5_9_reg_out :
  _guard21485 ? cond153_out :
  1'd0;
assign cond210_write_en = _guard21486;
assign cond210_clk = clk;
assign cond210_reset = reset;
assign cond210_in =
  _guard21487 ? idx_between_4_8_reg_out :
  1'd0;
assign cond218_write_en = _guard21488;
assign cond218_clk = clk;
assign cond218_reset = reset;
assign cond218_in =
  _guard21489 ? idx_between_6_10_reg_out :
  1'd0;
assign cond229_write_en = _guard21490;
assign cond229_clk = clk;
assign cond229_reset = reset;
assign cond229_in =
  _guard21491 ? idx_between_28_29_reg_out :
  1'd0;
assign cond_wire255_in =
  _guard21494 ? cond255_out :
  _guard21495 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire266_in =
  _guard21498 ? cond266_out :
  _guard21499 ? idx_between_18_22_reg_out :
  1'd0;
assign cond_wire272_in =
  _guard21500 ? idx_between_23_39_reg_out :
  _guard21503 ? cond272_out :
  1'd0;
assign cond_wire283_in =
  _guard21504 ? idx_between_7_11_reg_out :
  _guard21507 ? cond283_out :
  1'd0;
assign cond291_write_en = _guard21508;
assign cond291_clk = clk;
assign cond291_reset = reset;
assign cond291_in =
  _guard21509 ? idx_between_9_13_reg_out :
  1'd0;
assign cond295_write_en = _guard21510;
assign cond295_clk = clk;
assign cond295_reset = reset;
assign cond295_in =
  _guard21511 ? idx_between_10_14_reg_out :
  1'd0;
assign cond_wire297_in =
  _guard21512 ? idx_between_14_30_reg_out :
  _guard21515 ? cond297_out :
  1'd0;
assign cond_wire304_in =
  _guard21516 ? idx_between_12_28_reg_out :
  _guard21519 ? cond304_out :
  1'd0;
assign cond_wire320_in =
  _guard21520 ? idx_between_16_32_reg_out :
  _guard21523 ? cond320_out :
  1'd0;
assign cond327_write_en = _guard21524;
assign cond327_clk = clk;
assign cond327_reset = reset;
assign cond327_in =
  _guard21525 ? idx_between_18_22_reg_out :
  1'd0;
assign cond_wire331_in =
  _guard21526 ? idx_between_19_23_reg_out :
  _guard21529 ? cond331_out :
  1'd0;
assign cond345_write_en = _guard21530;
assign cond345_clk = clk;
assign cond345_reset = reset;
assign cond345_in =
  _guard21531 ? idx_between_7_23_reg_out :
  1'd0;
assign cond347_write_en = _guard21532;
assign cond347_clk = clk;
assign cond347_reset = reset;
assign cond347_in =
  _guard21533 ? idx_between_27_28_reg_out :
  1'd0;
assign cond_wire350_in =
  _guard21536 ? cond350_out :
  _guard21537 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire353_in =
  _guard21538 ? idx_between_9_25_reg_out :
  _guard21541 ? cond353_out :
  1'd0;
assign cond_wire369_in =
  _guard21542 ? idx_between_13_29_reg_out :
  _guard21545 ? cond369_out :
  1'd0;
assign cond_wire373_in =
  _guard21546 ? idx_between_14_30_reg_out :
  _guard21549 ? cond373_out :
  1'd0;
assign cond381_write_en = _guard21550;
assign cond381_clk = clk;
assign cond381_reset = reset;
assign cond381_in =
  _guard21551 ? idx_between_16_32_reg_out :
  1'd0;
assign cond_wire382_in =
  _guard21554 ? cond382_out :
  _guard21555 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire387_in =
  _guard21558 ? cond387_out :
  _guard21559 ? idx_between_37_38_reg_out :
  1'd0;
assign cond_wire397_in =
  _guard21562 ? cond397_out :
  _guard21563 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire400_in =
  _guard21564 ? idx_between_21_25_reg_out :
  _guard21567 ? cond400_out :
  1'd0;
assign cond403_write_en = _guard21568;
assign cond403_clk = clk;
assign cond403_reset = reset;
assign cond403_in =
  _guard21569 ? idx_between_41_42_reg_out :
  1'd0;
assign cond_wire406_in =
  _guard21570 ? idx_between_7_23_reg_out :
  _guard21573 ? cond406_out :
  1'd0;
assign cond409_write_en = _guard21574;
assign cond409_clk = clk;
assign cond409_reset = reset;
assign cond409_in =
  _guard21575 ? idx_between_8_12_reg_out :
  1'd0;
assign cond413_write_en = _guard21576;
assign cond413_clk = clk;
assign cond413_reset = reset;
assign cond413_in =
  _guard21577 ? idx_between_9_13_reg_out :
  1'd0;
assign cond422_write_en = _guard21578;
assign cond422_clk = clk;
assign cond422_reset = reset;
assign cond422_in =
  _guard21579 ? idx_between_11_27_reg_out :
  1'd0;
assign cond431_write_en = _guard21580;
assign cond431_clk = clk;
assign cond431_reset = reset;
assign cond431_in =
  _guard21581 ? idx_between_17_33_reg_out :
  1'd0;
assign cond456_write_en = _guard21582;
assign cond456_clk = clk;
assign cond456_reset = reset;
assign cond456_in =
  _guard21583 ? idx_between_39_40_reg_out :
  1'd0;
assign cond471_write_en = _guard21584;
assign cond471_clk = clk;
assign cond471_reset = reset;
assign cond471_in =
  _guard21585 ? idx_between_8_24_reg_out :
  1'd0;
assign cond_wire475_in =
  _guard21588 ? cond475_out :
  _guard21589 ? idx_between_9_25_reg_out :
  1'd0;
assign cond479_write_en = _guard21590;
assign cond479_clk = clk;
assign cond479_reset = reset;
assign cond479_in =
  _guard21591 ? idx_between_10_26_reg_out :
  1'd0;
assign cond_wire483_in =
  _guard21592 ? idx_between_11_27_reg_out :
  _guard21595 ? cond483_out :
  1'd0;
assign cond490_write_en = _guard21596;
assign cond490_clk = clk;
assign cond490_reset = reset;
assign cond490_in =
  _guard21597 ? idx_between_13_17_reg_out :
  1'd0;
assign cond493_write_en = _guard21598;
assign cond493_clk = clk;
assign cond493_reset = reset;
assign cond493_in =
  _guard21599 ? idx_between_33_34_reg_out :
  1'd0;
assign cond_wire499_in =
  _guard21602 ? cond499_out :
  _guard21603 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire507_in =
  _guard21604 ? idx_between_17_33_reg_out :
  _guard21607 ? cond507_out :
  1'd0;
assign cond512_write_en = _guard21608;
assign cond512_clk = clk;
assign cond512_reset = reset;
assign cond512_in =
  _guard21609 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire522_in =
  _guard21610 ? idx_between_21_25_reg_out :
  _guard21613 ? cond522_out :
  1'd0;
assign cond_wire539_in =
  _guard21616 ? cond539_out :
  _guard21617 ? idx_between_10_14_reg_out :
  1'd0;
assign cond564_write_en = _guard21618;
assign cond564_clk = clk;
assign cond564_reset = reset;
assign cond564_in =
  _guard21619 ? idx_between_16_32_reg_out :
  1'd0;
assign cond566_write_en = _guard21620;
assign cond566_clk = clk;
assign cond566_reset = reset;
assign cond566_in =
  _guard21621 ? idx_between_36_37_reg_out :
  1'd0;
assign cond_wire571_in =
  _guard21624 ? cond571_out :
  _guard21625 ? idx_between_18_22_reg_out :
  1'd0;
assign cond_wire590_in =
  _guard21626 ? idx_between_42_43_reg_out :
  _guard21629 ? cond590_out :
  1'd0;
assign cond593_write_en = _guard21630;
assign cond593_clk = clk;
assign cond593_reset = reset;
assign cond593_in =
  _guard21631 ? idx_between_27_43_reg_out :
  1'd0;
assign cond_wire601_in =
  _guard21634 ? cond601_out :
  _guard21635 ? idx_between_10_26_reg_out :
  1'd0;
assign cond623_write_en = _guard21636;
assign cond623_clk = clk;
assign cond623_reset = reset;
assign cond623_in =
  _guard21637 ? idx_between_35_36_reg_out :
  1'd0;
assign cond624_write_en = _guard21638;
assign cond624_clk = clk;
assign cond624_reset = reset;
assign cond624_in =
  _guard21639 ? idx_between_16_20_reg_out :
  1'd0;
assign cond_wire626_in =
  _guard21640 ? idx_between_20_36_reg_out :
  _guard21643 ? cond626_out :
  1'd0;
assign cond640_write_en = _guard21644;
assign cond640_clk = clk;
assign cond640_reset = reset;
assign cond640_in =
  _guard21645 ? idx_between_20_24_reg_out :
  1'd0;
assign cond641_write_en = _guard21646;
assign cond641_clk = clk;
assign cond641_reset = reset;
assign cond641_in =
  _guard21647 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire650_in =
  _guard21650 ? cond650_out :
  _guard21651 ? idx_between_26_42_reg_out :
  1'd0;
assign cond_wire664_in =
  _guard21654 ? cond664_out :
  _guard21655 ? idx_between_10_26_reg_out :
  1'd0;
assign cond671_write_en = _guard21656;
assign cond671_clk = clk;
assign cond671_reset = reset;
assign cond671_in =
  _guard21657 ? idx_between_16_32_reg_out :
  1'd0;
assign cond_wire676_in =
  _guard21658 ? idx_between_33_34_reg_out :
  _guard21661 ? cond676_out :
  1'd0;
assign cond_wire679_in =
  _guard21664 ? cond679_out :
  _guard21665 ? idx_between_18_34_reg_out :
  1'd0;
assign cond688_write_en = _guard21666;
assign cond688_clk = clk;
assign cond688_reset = reset;
assign cond688_in =
  _guard21667 ? idx_between_36_37_reg_out :
  1'd0;
assign cond_wire694_in =
  _guard21668 ? idx_between_18_34_reg_out :
  _guard21671 ? cond694_out :
  1'd0;
assign cond698_write_en = _guard21672;
assign cond698_clk = clk;
assign cond698_reset = reset;
assign cond698_in =
  _guard21673 ? idx_between_19_35_reg_out :
  1'd0;
assign cond700_write_en = _guard21674;
assign cond700_clk = clk;
assign cond700_reset = reset;
assign cond700_in =
  _guard21675 ? idx_between_39_40_reg_out :
  1'd0;
assign cond724_write_en = _guard21676;
assign cond724_clk = clk;
assign cond724_reset = reset;
assign cond724_in =
  _guard21677 ? idx_between_45_46_reg_out :
  1'd0;
assign cond_wire731_in =
  _guard21678 ? idx_between_12_28_reg_out :
  _guard21681 ? cond731_out :
  1'd0;
assign cond739_write_en = _guard21682;
assign cond739_clk = clk;
assign cond739_reset = reset;
assign cond739_in =
  _guard21683 ? idx_between_14_30_reg_out :
  1'd0;
assign cond749_write_en = _guard21684;
assign cond749_clk = clk;
assign cond749_reset = reset;
assign cond749_in =
  _guard21685 ? idx_between_36_37_reg_out :
  1'd0;
assign cond_wire754_in =
  _guard21688 ? cond754_out :
  _guard21689 ? idx_between_18_22_reg_out :
  1'd0;
assign cond_wire772_in =
  _guard21692 ? cond772_out :
  _guard21693 ? idx_between_26_42_reg_out :
  1'd0;
assign cond810_write_en = _guard21694;
assign cond810_clk = clk;
assign cond810_reset = reset;
assign cond810_in =
  _guard21695 ? idx_between_36_37_reg_out :
  1'd0;
assign cond_wire813_in =
  _guard21696 ? idx_between_21_37_reg_out :
  _guard21699 ? cond813_out :
  1'd0;
assign cond_wire816_in =
  _guard21700 ? idx_between_18_34_reg_out :
  _guard21703 ? cond816_out :
  1'd0;
assign cond_wire824_in =
  _guard21704 ? idx_between_20_36_reg_out :
  _guard21707 ? cond824_out :
  1'd0;
assign cond825_write_en = _guard21708;
assign cond825_clk = clk;
assign cond825_reset = reset;
assign cond825_in =
  _guard21709 ? idx_between_24_40_reg_out :
  1'd0;
assign cond_wire827_in =
  _guard21712 ? cond827_out :
  _guard21713 ? idx_between_21_25_reg_out :
  1'd0;
assign cond849_write_en = _guard21714;
assign cond849_clk = clk;
assign cond849_reset = reset;
assign cond849_in =
  _guard21715 ? idx_between_30_46_reg_out :
  1'd0;
assign cond873_write_en = _guard21716;
assign cond873_clk = clk;
assign cond873_reset = reset;
assign cond873_in =
  _guard21717 ? idx_between_17_33_reg_out :
  1'd0;
assign cond886_write_en = _guard21718;
assign cond886_clk = clk;
assign cond886_reset = reset;
assign cond886_in =
  _guard21719 ? idx_between_24_40_reg_out :
  1'd0;
assign cond_wire902_in =
  _guard21722 ? cond902_out :
  _guard21723 ? idx_between_28_44_reg_out :
  1'd0;
assign cond_wire921_in =
  _guard21726 ? cond921_out :
  _guard21727 ? idx_between_29_45_reg_out :
  1'd0;
assign cond_wire926_in =
  _guard21730 ? cond926_out :
  _guard21731 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire947_in =
  _guard21734 ? cond947_out :
  _guard21735 ? idx_between_24_40_reg_out :
  1'd0;
assign cond_wire950_in =
  _guard21738 ? cond950_out :
  _guard21739 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire953_in =
  _guard21742 ? cond953_out :
  _guard21743 ? idx_between_22_26_reg_out :
  1'd0;
assign cond_wire963_in =
  _guard21746 ? cond963_out :
  _guard21747 ? idx_between_28_44_reg_out :
  1'd0;
assign cond_wire971_in =
  _guard21748 ? idx_between_30_46_reg_out :
  _guard21751 ? cond971_out :
  1'd0;
assign cond_wire975_in =
  _guard21752 ? idx_between_31_47_reg_out :
  _guard21755 ? cond975_out :
  1'd0;
assign cond_wire988_in =
  _guard21756 ? idx_between_50_51_reg_out :
  _guard21759 ? cond988_out :
  1'd0;
assign cond990_write_en = _guard21760;
assign cond990_clk = clk;
assign cond990_reset = reset;
assign cond990_in =
  _guard21761 ? idx_between_16_20_reg_out :
  1'd0;
assign cond_wire997_in =
  _guard21764 ? cond997_out :
  _guard21765 ? idx_between_37_38_reg_out :
  1'd0;
assign cond_wire1000_in =
  _guard21768 ? cond1000_out :
  _guard21769 ? idx_between_22_38_reg_out :
  1'd0;
assign cond1009_write_en = _guard21770;
assign cond1009_clk = clk;
assign cond1009_reset = reset;
assign cond1009_in =
  _guard21771 ? idx_between_40_41_reg_out :
  1'd0;
assign cond_wire1012_in =
  _guard21774 ? cond1012_out :
  _guard21775 ? idx_between_25_41_reg_out :
  1'd0;
assign cond1014_write_en = _guard21776;
assign cond1014_clk = clk;
assign cond1014_reset = reset;
assign cond1014_in =
  _guard21777 ? idx_between_22_26_reg_out :
  1'd0;
assign cond_wire1025_in =
  _guard21778 ? idx_between_44_45_reg_out :
  _guard21781 ? cond1025_out :
  1'd0;
assign cond1027_write_en = _guard21782;
assign cond1027_clk = clk;
assign cond1027_reset = reset;
assign cond1027_in =
  _guard21783 ? idx_between_25_41_reg_out :
  1'd0;
assign cond1035_write_en = _guard21784;
assign cond1035_clk = clk;
assign cond1035_reset = reset;
assign cond1035_in =
  _guard21785 ? idx_between_27_43_reg_out :
  1'd0;
assign early_reset_static_seq_done_in = ud_out;
assign top_0_3_write_en = _guard21788;
assign top_0_3_clk = clk;
assign top_0_3_reset = reset;
assign top_0_3_in = t3_read_data;
assign pe_0_6_mul_ready =
  _guard21794 ? 1'd1 :
  _guard21797 ? 1'd0 :
  1'd0;
assign pe_0_6_clk = clk;
assign pe_0_6_top =
  _guard21810 ? top_0_6_out :
  32'd0;
assign pe_0_6_left =
  _guard21823 ? left_0_6_out :
  32'd0;
assign pe_0_6_reset = reset;
assign pe_0_6_go = _guard21836;
assign top_1_7_write_en = _guard21839;
assign top_1_7_clk = clk;
assign top_1_7_reset = reset;
assign top_1_7_in = top_0_7_out;
assign top_1_12_write_en = _guard21845;
assign top_1_12_clk = clk;
assign top_1_12_reset = reset;
assign top_1_12_in = top_0_12_out;
assign left_1_15_write_en = _guard21851;
assign left_1_15_clk = clk;
assign left_1_15_reset = reset;
assign left_1_15_in = left_1_14_out;
assign top_2_1_write_en = _guard21857;
assign top_2_1_clk = clk;
assign top_2_1_reset = reset;
assign top_2_1_in = top_1_1_out;
assign top_2_10_write_en = _guard21863;
assign top_2_10_clk = clk;
assign top_2_10_reset = reset;
assign top_2_10_in = top_1_10_out;
assign left_3_3_write_en = _guard21869;
assign left_3_3_clk = clk;
assign left_3_3_reset = reset;
assign left_3_3_in = left_3_2_out;
assign top_3_7_write_en = _guard21875;
assign top_3_7_clk = clk;
assign top_3_7_reset = reset;
assign top_3_7_in = top_2_7_out;
assign top_3_13_write_en = _guard21881;
assign top_3_13_clk = clk;
assign top_3_13_reset = reset;
assign top_3_13_in = top_2_13_out;
assign left_4_1_write_en = _guard21887;
assign left_4_1_clk = clk;
assign left_4_1_reset = reset;
assign left_4_1_in = left_4_0_out;
assign pe_4_3_mul_ready =
  _guard21893 ? 1'd1 :
  _guard21896 ? 1'd0 :
  1'd0;
assign pe_4_3_clk = clk;
assign pe_4_3_top =
  _guard21909 ? top_4_3_out :
  32'd0;
assign pe_4_3_left =
  _guard21922 ? left_4_3_out :
  32'd0;
assign pe_4_3_reset = reset;
assign pe_4_3_go = _guard21935;
assign top_4_8_write_en = _guard21938;
assign top_4_8_clk = clk;
assign top_4_8_reset = reset;
assign top_4_8_in = top_3_8_out;
assign pe_4_10_mul_ready =
  _guard21944 ? 1'd1 :
  _guard21947 ? 1'd0 :
  1'd0;
assign pe_4_10_clk = clk;
assign pe_4_10_top =
  _guard21960 ? top_4_10_out :
  32'd0;
assign pe_4_10_left =
  _guard21973 ? left_4_10_out :
  32'd0;
assign pe_4_10_reset = reset;
assign pe_4_10_go = _guard21986;
assign top_4_14_write_en = _guard21989;
assign top_4_14_clk = clk;
assign top_4_14_reset = reset;
assign top_4_14_in = top_3_14_out;
assign left_5_0_write_en = _guard21995;
assign left_5_0_clk = clk;
assign left_5_0_reset = reset;
assign left_5_0_in = l5_read_data;
assign pe_5_11_mul_ready =
  _guard22001 ? 1'd1 :
  _guard22004 ? 1'd0 :
  1'd0;
assign pe_5_11_clk = clk;
assign pe_5_11_top =
  _guard22017 ? top_5_11_out :
  32'd0;
assign pe_5_11_left =
  _guard22030 ? left_5_11_out :
  32'd0;
assign pe_5_11_reset = reset;
assign pe_5_11_go = _guard22043;
assign top_5_12_write_en = _guard22046;
assign top_5_12_clk = clk;
assign top_5_12_reset = reset;
assign top_5_12_in = top_4_12_out;
assign left_5_12_write_en = _guard22052;
assign left_5_12_clk = clk;
assign left_5_12_reset = reset;
assign left_5_12_in = left_5_11_out;
assign pe_5_15_mul_ready =
  _guard22058 ? 1'd1 :
  _guard22061 ? 1'd0 :
  1'd0;
assign pe_5_15_clk = clk;
assign pe_5_15_top =
  _guard22074 ? top_5_15_out :
  32'd0;
assign pe_5_15_left =
  _guard22087 ? left_5_15_out :
  32'd0;
assign pe_5_15_reset = reset;
assign pe_5_15_go = _guard22100;
assign pe_6_6_mul_ready =
  _guard22103 ? 1'd1 :
  _guard22106 ? 1'd0 :
  1'd0;
assign pe_6_6_clk = clk;
assign pe_6_6_top =
  _guard22119 ? top_6_6_out :
  32'd0;
assign pe_6_6_left =
  _guard22132 ? left_6_6_out :
  32'd0;
assign pe_6_6_reset = reset;
assign pe_6_6_go = _guard22145;
assign top_6_9_write_en = _guard22148;
assign top_6_9_clk = clk;
assign top_6_9_reset = reset;
assign top_6_9_in = top_5_9_out;
assign pe_7_2_mul_ready =
  _guard22154 ? 1'd1 :
  _guard22157 ? 1'd0 :
  1'd0;
assign pe_7_2_clk = clk;
assign pe_7_2_top =
  _guard22170 ? top_7_2_out :
  32'd0;
assign pe_7_2_left =
  _guard22183 ? left_7_2_out :
  32'd0;
assign pe_7_2_reset = reset;
assign pe_7_2_go = _guard22196;
assign pe_7_7_mul_ready =
  _guard22199 ? 1'd1 :
  _guard22202 ? 1'd0 :
  1'd0;
assign pe_7_7_clk = clk;
assign pe_7_7_top =
  _guard22215 ? top_7_7_out :
  32'd0;
assign pe_7_7_left =
  _guard22228 ? left_7_7_out :
  32'd0;
assign pe_7_7_reset = reset;
assign pe_7_7_go = _guard22241;
assign top_7_9_write_en = _guard22244;
assign top_7_9_clk = clk;
assign top_7_9_reset = reset;
assign top_7_9_in = top_6_9_out;
assign top_7_14_write_en = _guard22250;
assign top_7_14_clk = clk;
assign top_7_14_reset = reset;
assign top_7_14_in = top_6_14_out;
assign top_7_15_write_en = _guard22256;
assign top_7_15_clk = clk;
assign top_7_15_reset = reset;
assign top_7_15_in = top_6_15_out;
assign left_8_1_write_en = _guard22262;
assign left_8_1_clk = clk;
assign left_8_1_reset = reset;
assign left_8_1_in = left_8_0_out;
assign pe_8_10_mul_ready =
  _guard22268 ? 1'd1 :
  _guard22271 ? 1'd0 :
  1'd0;
assign pe_8_10_clk = clk;
assign pe_8_10_top =
  _guard22284 ? top_8_10_out :
  32'd0;
assign pe_8_10_left =
  _guard22297 ? left_8_10_out :
  32'd0;
assign pe_8_10_reset = reset;
assign pe_8_10_go = _guard22310;
assign left_8_13_write_en = _guard22313;
assign left_8_13_clk = clk;
assign left_8_13_reset = reset;
assign left_8_13_in = left_8_12_out;
assign pe_8_14_mul_ready =
  _guard22319 ? 1'd1 :
  _guard22322 ? 1'd0 :
  1'd0;
assign pe_8_14_clk = clk;
assign pe_8_14_top =
  _guard22335 ? top_8_14_out :
  32'd0;
assign pe_8_14_left =
  _guard22348 ? left_8_14_out :
  32'd0;
assign pe_8_14_reset = reset;
assign pe_8_14_go = _guard22361;
assign top_9_2_write_en = _guard22364;
assign top_9_2_clk = clk;
assign top_9_2_reset = reset;
assign top_9_2_in = top_8_2_out;
assign left_9_11_write_en = _guard22370;
assign left_9_11_clk = clk;
assign left_9_11_reset = reset;
assign left_9_11_in = left_9_10_out;
assign left_10_1_write_en = _guard22376;
assign left_10_1_clk = clk;
assign left_10_1_reset = reset;
assign left_10_1_in = left_10_0_out;
assign pe_10_11_mul_ready =
  _guard22382 ? 1'd1 :
  _guard22385 ? 1'd0 :
  1'd0;
assign pe_10_11_clk = clk;
assign pe_10_11_top =
  _guard22398 ? top_10_11_out :
  32'd0;
assign pe_10_11_left =
  _guard22411 ? left_10_11_out :
  32'd0;
assign pe_10_11_reset = reset;
assign pe_10_11_go = _guard22424;
assign top_10_11_write_en = _guard22427;
assign top_10_11_clk = clk;
assign top_10_11_reset = reset;
assign top_10_11_in = top_9_11_out;
assign left_10_12_write_en = _guard22433;
assign left_10_12_clk = clk;
assign left_10_12_reset = reset;
assign left_10_12_in = left_10_11_out;
assign top_11_0_write_en = _guard22439;
assign top_11_0_clk = clk;
assign top_11_0_reset = reset;
assign top_11_0_in = top_10_0_out;
assign left_11_1_write_en = _guard22445;
assign left_11_1_clk = clk;
assign left_11_1_reset = reset;
assign left_11_1_in = left_11_0_out;
assign pe_11_10_mul_ready =
  _guard22451 ? 1'd1 :
  _guard22454 ? 1'd0 :
  1'd0;
assign pe_11_10_clk = clk;
assign pe_11_10_top =
  _guard22467 ? top_11_10_out :
  32'd0;
assign pe_11_10_left =
  _guard22480 ? left_11_10_out :
  32'd0;
assign pe_11_10_reset = reset;
assign pe_11_10_go = _guard22493;
assign top_13_14_write_en = _guard22496;
assign top_13_14_clk = clk;
assign top_13_14_reset = reset;
assign top_13_14_in = top_12_14_out;
assign left_14_0_write_en = _guard22502;
assign left_14_0_clk = clk;
assign left_14_0_reset = reset;
assign left_14_0_in = l14_read_data;
assign top_14_2_write_en = _guard22508;
assign top_14_2_clk = clk;
assign top_14_2_reset = reset;
assign top_14_2_in = top_13_2_out;
assign top_14_3_write_en = _guard22514;
assign top_14_3_clk = clk;
assign top_14_3_reset = reset;
assign top_14_3_in = top_13_3_out;
assign left_15_4_write_en = _guard22520;
assign left_15_4_clk = clk;
assign left_15_4_reset = reset;
assign left_15_4_in = left_15_3_out;
assign pe_15_7_mul_ready =
  _guard22526 ? 1'd1 :
  _guard22529 ? 1'd0 :
  1'd0;
assign pe_15_7_clk = clk;
assign pe_15_7_top =
  _guard22542 ? top_15_7_out :
  32'd0;
assign pe_15_7_left =
  _guard22555 ? left_15_7_out :
  32'd0;
assign pe_15_7_reset = reset;
assign pe_15_7_go = _guard22568;
assign t2_idx_write_en = _guard22575;
assign t2_idx_clk = clk;
assign t2_idx_reset = reset;
assign t2_idx_in =
  _guard22578 ? 5'd0 :
  _guard22581 ? t2_add_out :
  'x;
assign t11_add_left = 5'd1;
assign t11_add_right = t11_idx_out;
assign l2_idx_write_en = _guard22594;
assign l2_idx_clk = clk;
assign l2_idx_reset = reset;
assign l2_idx_in =
  _guard22597 ? 5'd0 :
  _guard22600 ? l2_add_out :
  'x;
assign l6_idx_write_en = _guard22607;
assign l6_idx_clk = clk;
assign l6_idx_reset = reset;
assign l6_idx_in =
  _guard22610 ? 5'd0 :
  _guard22613 ? l6_add_out :
  'x;
assign l14_add_left = 5'd1;
assign l14_add_right = l14_idx_out;
assign index_ge_26_left = idx_add_out;
assign index_ge_26_right = 6'd26;
assign index_lt_41_left = idx_add_out;
assign index_lt_41_right = 6'd41;
assign idx_between_40_41_reg_write_en = _guard22628;
assign idx_between_40_41_reg_clk = clk;
assign idx_between_40_41_reg_reset = reset;
assign idx_between_40_41_reg_in =
  _guard22631 ? 1'd0 :
  _guard22632 ? idx_between_40_41_comb_out :
  'x;
assign index_ge_27_left = idx_add_out;
assign index_ge_27_right = 6'd27;
assign idx_between_24_28_reg_write_en = _guard22639;
assign idx_between_24_28_reg_clk = clk;
assign idx_between_24_28_reg_reset = reset;
assign idx_between_24_28_reg_in =
  _guard22642 ? 1'd0 :
  _guard22643 ? idx_between_24_28_comb_out :
  'x;
assign idx_between_24_28_comb_left = index_ge_24_out;
assign idx_between_24_28_comb_right = index_lt_28_out;
assign index_lt_29_left = idx_add_out;
assign index_lt_29_right = 6'd29;
assign index_ge_45_left = idx_add_out;
assign index_ge_45_right = 6'd45;
assign idx_between_46_47_reg_write_en = _guard22654;
assign idx_between_46_47_reg_clk = clk;
assign idx_between_46_47_reg_reset = reset;
assign idx_between_46_47_reg_in =
  _guard22655 ? idx_between_46_47_comb_out :
  _guard22658 ? 1'd0 :
  'x;
assign index_lt_32_left = idx_add_out;
assign index_lt_32_right = 6'd32;
assign index_ge_6_left = idx_add_out;
assign index_ge_6_right = 6'd6;
assign idx_between_30_31_reg_write_en = _guard22667;
assign idx_between_30_31_reg_clk = clk;
assign idx_between_30_31_reg_reset = reset;
assign idx_between_30_31_reg_in =
  _guard22668 ? idx_between_30_31_comb_out :
  _guard22671 ? 1'd0 :
  'x;
assign idx_between_25_26_comb_left = index_ge_25_out;
assign idx_between_25_26_comb_right = index_lt_26_out;
assign index_lt_7_left = idx_add_out;
assign index_lt_7_right = 6'd7;
assign idx_between_8_24_reg_write_en = _guard22680;
assign idx_between_8_24_reg_clk = clk;
assign idx_between_8_24_reg_reset = reset;
assign idx_between_8_24_reg_in =
  _guard22683 ? 1'd0 :
  _guard22684 ? idx_between_8_24_comb_out :
  'x;
assign idx_between_9_25_reg_write_en = _guard22689;
assign idx_between_9_25_reg_clk = clk;
assign idx_between_9_25_reg_reset = reset;
assign idx_between_9_25_reg_in =
  _guard22692 ? 1'd0 :
  _guard22693 ? idx_between_9_25_comb_out :
  'x;
assign idx_between_15_31_comb_left = index_ge_15_out;
assign idx_between_15_31_comb_right = index_lt_31_out;
assign idx_between_29_30_comb_left = index_ge_29_out;
assign idx_between_29_30_comb_right = index_lt_30_out;
assign index_ge_36_left = idx_add_out;
assign index_ge_36_right = 6'd36;
assign idx_between_39_40_reg_write_en = _guard22704;
assign idx_between_39_40_reg_clk = clk;
assign idx_between_39_40_reg_reset = reset;
assign idx_between_39_40_reg_in =
  _guard22705 ? idx_between_39_40_comb_out :
  _guard22708 ? 1'd0 :
  'x;
assign cond1_write_en = _guard22709;
assign cond1_clk = clk;
assign cond1_reset = reset;
assign cond1_in =
  _guard22710 ? idx_between_1_17_reg_out :
  1'd0;
assign cond2_write_en = _guard22711;
assign cond2_clk = clk;
assign cond2_reset = reset;
assign cond2_in =
  _guard22712 ? idx_between_5_21_reg_out :
  1'd0;
assign cond_wire5_in =
  _guard22715 ? cond5_out :
  _guard22716 ? idx_between_2_6_reg_out :
  1'd0;
assign cond22_write_en = _guard22717;
assign cond22_clk = clk;
assign cond22_reset = reset;
assign cond22_in =
  _guard22718 ? idx_between_9_25_reg_out :
  1'd0;
assign cond26_write_en = _guard22719;
assign cond26_clk = clk;
assign cond26_reset = reset;
assign cond26_in =
  _guard22720 ? idx_between_6_22_reg_out :
  1'd0;
assign cond_wire34_in =
  _guard22721 ? idx_between_7_23_reg_out :
  _guard22724 ? cond34_out :
  1'd0;
assign cond39_write_en = _guard22725;
assign cond39_clk = clk;
assign cond39_reset = reset;
assign cond39_in =
  _guard22726 ? idx_between_8_24_reg_out :
  1'd0;
assign cond49_write_en = _guard22727;
assign cond49_clk = clk;
assign cond49_reset = reset;
assign cond49_in =
  _guard22728 ? idx_between_10_26_reg_out :
  1'd0;
assign cond_wire52_in =
  _guard22731 ? cond52_out :
  _guard22732 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire68_in =
  _guard22733 ? idx_between_34_35_reg_out :
  _guard22736 ? cond68_out :
  1'd0;
assign cond_wire70_in =
  _guard22737 ? idx_between_15_19_reg_out :
  _guard22740 ? cond70_out :
  1'd0;
assign cond_wire83_in =
  _guard22741 ? idx_between_22_23_reg_out :
  _guard22744 ? cond83_out :
  1'd0;
assign cond87_write_en = _guard22745;
assign cond87_clk = clk;
assign cond87_reset = reset;
assign cond87_in =
  _guard22746 ? idx_between_23_24_reg_out :
  1'd0;
assign cond96_write_en = _guard22747;
assign cond96_clk = clk;
assign cond96_reset = reset;
assign cond96_in =
  _guard22748 ? idx_between_6_10_reg_out :
  1'd0;
assign cond_wire97_in =
  _guard22749 ? idx_between_6_22_reg_out :
  _guard22752 ? cond97_out :
  1'd0;
assign cond99_write_en = _guard22753;
assign cond99_clk = clk;
assign cond99_reset = reset;
assign cond99_in =
  _guard22754 ? idx_between_26_27_reg_out :
  1'd0;
assign cond104_write_en = _guard22755;
assign cond104_clk = clk;
assign cond104_reset = reset;
assign cond104_in =
  _guard22756 ? idx_between_8_12_reg_out :
  1'd0;
assign cond133_write_en = _guard22757;
assign cond133_clk = clk;
assign cond133_reset = reset;
assign cond133_in =
  _guard22758 ? idx_between_15_31_reg_out :
  1'd0;
assign cond138_write_en = _guard22759;
assign cond138_clk = clk;
assign cond138_reset = reset;
assign cond138_in =
  _guard22760 ? idx_between_20_36_reg_out :
  1'd0;
assign cond145_write_en = _guard22761;
assign cond145_clk = clk;
assign cond145_reset = reset;
assign cond145_in =
  _guard22762 ? idx_between_3_7_reg_out :
  1'd0;
assign cond147_write_en = _guard22763;
assign cond147_clk = clk;
assign cond147_reset = reset;
assign cond147_in =
  _guard22764 ? idx_between_7_23_reg_out :
  1'd0;
assign cond_wire147_in =
  _guard22765 ? idx_between_7_23_reg_out :
  _guard22768 ? cond147_out :
  1'd0;
assign cond154_write_en = _guard22769;
assign cond154_clk = clk;
assign cond154_reset = reset;
assign cond154_in =
  _guard22770 ? idx_between_5_21_reg_out :
  1'd0;
assign cond156_write_en = _guard22771;
assign cond156_clk = clk;
assign cond156_reset = reset;
assign cond156_in =
  _guard22772 ? idx_between_25_26_reg_out :
  1'd0;
assign cond_wire168_in =
  _guard22775 ? cond168_out :
  _guard22776 ? idx_between_28_29_reg_out :
  1'd0;
assign cond173_write_en = _guard22777;
assign cond173_clk = clk;
assign cond173_reset = reset;
assign cond173_in =
  _guard22778 ? idx_between_10_14_reg_out :
  1'd0;
assign cond175_write_en = _guard22779;
assign cond175_clk = clk;
assign cond175_reset = reset;
assign cond175_in =
  _guard22780 ? idx_between_14_30_reg_out :
  1'd0;
assign cond182_write_en = _guard22781;
assign cond182_clk = clk;
assign cond182_reset = reset;
assign cond182_in =
  _guard22782 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire199_in =
  _guard22783 ? idx_between_20_36_reg_out :
  _guard22786 ? cond199_out :
  1'd0;
assign cond_wire206_in =
  _guard22789 ? cond206_out :
  _guard22790 ? idx_between_18_34_reg_out :
  1'd0;
assign cond212_write_en = _guard22791;
assign cond212_clk = clk;
assign cond212_reset = reset;
assign cond212_in =
  _guard22792 ? idx_between_8_24_reg_out :
  1'd0;
assign cond_wire212_in =
  _guard22793 ? idx_between_8_24_reg_out :
  _guard22796 ? cond212_out :
  1'd0;
assign cond224_write_en = _guard22797;
assign cond224_clk = clk;
assign cond224_reset = reset;
assign cond224_in =
  _guard22798 ? idx_between_11_27_reg_out :
  1'd0;
assign cond_wire229_in =
  _guard22801 ? cond229_out :
  _guard22802 ? idx_between_28_29_reg_out :
  1'd0;
assign cond_wire232_in =
  _guard22803 ? idx_between_13_29_reg_out :
  _guard22806 ? cond232_out :
  1'd0;
assign cond_wire247_in =
  _guard22807 ? idx_between_13_29_reg_out :
  _guard22810 ? cond247_out :
  1'd0;
assign cond259_write_en = _guard22811;
assign cond259_clk = clk;
assign cond259_reset = reset;
assign cond259_in =
  _guard22812 ? idx_between_16_32_reg_out :
  1'd0;
assign cond_wire259_in =
  _guard22813 ? idx_between_16_32_reg_out :
  _guard22816 ? cond259_out :
  1'd0;
assign cond260_write_en = _guard22817;
assign cond260_clk = clk;
assign cond260_reset = reset;
assign cond260_in =
  _guard22818 ? idx_between_20_36_reg_out :
  1'd0;
assign cond273_write_en = _guard22819;
assign cond273_clk = clk;
assign cond273_reset = reset;
assign cond273_in =
  _guard22820 ? idx_between_39_40_reg_out :
  1'd0;
assign cond_wire277_in =
  _guard22823 ? cond277_out :
  _guard22824 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire280_in =
  _guard22825 ? idx_between_6_22_reg_out :
  _guard22828 ? cond280_out :
  1'd0;
assign cond303_write_en = _guard22829;
assign cond303_clk = clk;
assign cond303_reset = reset;
assign cond303_in =
  _guard22830 ? idx_between_12_16_reg_out :
  1'd0;
assign cond306_write_en = _guard22831;
assign cond306_clk = clk;
assign cond306_reset = reset;
assign cond306_in =
  _guard22832 ? idx_between_32_33_reg_out :
  1'd0;
assign cond310_write_en = _guard22833;
assign cond310_clk = clk;
assign cond310_reset = reset;
assign cond310_in =
  _guard22834 ? idx_between_33_34_reg_out :
  1'd0;
assign cond326_write_en = _guard22835;
assign cond326_clk = clk;
assign cond326_reset = reset;
assign cond326_in =
  _guard22836 ? idx_between_37_38_reg_out :
  1'd0;
assign cond328_write_en = _guard22837;
assign cond328_clk = clk;
assign cond328_reset = reset;
assign cond328_in =
  _guard22838 ? idx_between_18_34_reg_out :
  1'd0;
assign cond337_write_en = _guard22839;
assign cond337_clk = clk;
assign cond337_reset = reset;
assign cond337_in =
  _guard22840 ? idx_between_24_40_reg_out :
  1'd0;
assign cond339_write_en = _guard22841;
assign cond339_clk = clk;
assign cond339_reset = reset;
assign cond339_in =
  _guard22842 ? idx_between_5_21_reg_out :
  1'd0;
assign cond_wire360_in =
  _guard22845 ? cond360_out :
  _guard22846 ? idx_between_11_15_reg_out :
  1'd0;
assign cond361_write_en = _guard22847;
assign cond361_clk = clk;
assign cond361_reset = reset;
assign cond361_in =
  _guard22848 ? idx_between_11_27_reg_out :
  1'd0;
assign cond392_write_en = _guard22849;
assign cond392_clk = clk;
assign cond392_reset = reset;
assign cond392_in =
  _guard22850 ? idx_between_19_23_reg_out :
  1'd0;
assign cond399_write_en = _guard22851;
assign cond399_clk = clk;
assign cond399_reset = reset;
assign cond399_in =
  _guard22852 ? idx_between_40_41_reg_out :
  1'd0;
assign cond401_write_en = _guard22853;
assign cond401_clk = clk;
assign cond401_reset = reset;
assign cond401_in =
  _guard22854 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire407_in =
  _guard22855 ? idx_between_11_27_reg_out :
  _guard22858 ? cond407_out :
  1'd0;
assign cond_wire414_in =
  _guard22861 ? cond414_out :
  _guard22862 ? idx_between_9_25_reg_out :
  1'd0;
assign cond418_write_en = _guard22863;
assign cond418_clk = clk;
assign cond418_reset = reset;
assign cond418_in =
  _guard22864 ? idx_between_10_26_reg_out :
  1'd0;
assign cond423_write_en = _guard22865;
assign cond423_clk = clk;
assign cond423_reset = reset;
assign cond423_in =
  _guard22866 ? idx_between_15_31_reg_out :
  1'd0;
assign cond430_write_en = _guard22867;
assign cond430_clk = clk;
assign cond430_reset = reset;
assign cond430_in =
  _guard22868 ? idx_between_13_29_reg_out :
  1'd0;
assign cond_wire435_in =
  _guard22871 ? cond435_out :
  _guard22872 ? idx_between_18_34_reg_out :
  1'd0;
assign cond447_write_en = _guard22873;
assign cond447_clk = clk;
assign cond447_reset = reset;
assign cond447_in =
  _guard22874 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire448_in =
  _guard22877 ? cond448_out :
  _guard22878 ? idx_between_37_38_reg_out :
  1'd0;
assign cond_wire450_in =
  _guard22879 ? idx_between_18_34_reg_out :
  _guard22882 ? cond450_out :
  1'd0;
assign cond_wire454_in =
  _guard22885 ? cond454_out :
  _guard22886 ? idx_between_19_35_reg_out :
  1'd0;
assign cond469_write_en = _guard22887;
assign cond469_clk = clk;
assign cond469_reset = reset;
assign cond469_in =
  _guard22888 ? idx_between_7_23_reg_out :
  1'd0;
assign cond470_write_en = _guard22889;
assign cond470_clk = clk;
assign cond470_reset = reset;
assign cond470_in =
  _guard22890 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire480_in =
  _guard22891 ? idx_between_14_30_reg_out :
  _guard22894 ? cond480_out :
  1'd0;
assign cond483_write_en = _guard22895;
assign cond483_clk = clk;
assign cond483_reset = reset;
assign cond483_in =
  _guard22896 ? idx_between_11_27_reg_out :
  1'd0;
assign cond487_write_en = _guard22897;
assign cond487_clk = clk;
assign cond487_reset = reset;
assign cond487_in =
  _guard22898 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire488_in =
  _guard22899 ? idx_between_16_32_reg_out :
  _guard22902 ? cond488_out :
  1'd0;
assign cond491_write_en = _guard22903;
assign cond491_clk = clk;
assign cond491_reset = reset;
assign cond491_in =
  _guard22904 ? idx_between_13_29_reg_out :
  1'd0;
assign cond492_write_en = _guard22905;
assign cond492_clk = clk;
assign cond492_reset = reset;
assign cond492_in =
  _guard22906 ? idx_between_17_33_reg_out :
  1'd0;
assign cond505_write_en = _guard22907;
assign cond505_clk = clk;
assign cond505_reset = reset;
assign cond505_in =
  _guard22908 ? idx_between_36_37_reg_out :
  1'd0;
assign cond_wire513_in =
  _guard22911 ? cond513_out :
  _guard22912 ? idx_between_38_39_reg_out :
  1'd0;
assign cond_wire515_in =
  _guard22915 ? cond515_out :
  _guard22916 ? idx_between_19_35_reg_out :
  1'd0;
assign cond519_write_en = _guard22917;
assign cond519_clk = clk;
assign cond519_reset = reset;
assign cond519_in =
  _guard22918 ? idx_between_20_36_reg_out :
  1'd0;
assign cond_wire531_in =
  _guard22919 ? idx_between_23_39_reg_out :
  _guard22922 ? cond531_out :
  1'd0;
assign cond534_write_en = _guard22923;
assign cond534_clk = clk;
assign cond534_reset = reset;
assign cond534_in =
  _guard22924 ? idx_between_8_24_reg_out :
  1'd0;
assign cond_wire536_in =
  _guard22927 ? cond536_out :
  _guard22928 ? idx_between_9_25_reg_out :
  1'd0;
assign cond540_write_en = _guard22929;
assign cond540_clk = clk;
assign cond540_reset = reset;
assign cond540_in =
  _guard22930 ? idx_between_10_26_reg_out :
  1'd0;
assign cond_wire548_in =
  _guard22931 ? idx_between_12_28_reg_out :
  _guard22934 ? cond548_out :
  1'd0;
assign cond_wire551_in =
  _guard22937 ? cond551_out :
  _guard22938 ? idx_between_13_17_reg_out :
  1'd0;
assign cond555_write_en = _guard22939;
assign cond555_clk = clk;
assign cond555_reset = reset;
assign cond555_in =
  _guard22940 ? idx_between_14_18_reg_out :
  1'd0;
assign cond_wire557_in =
  _guard22941 ? idx_between_18_34_reg_out :
  _guard22944 ? cond557_out :
  1'd0;
assign cond562_write_en = _guard22945;
assign cond562_clk = clk;
assign cond562_reset = reset;
assign cond562_in =
  _guard22946 ? idx_between_35_36_reg_out :
  1'd0;
assign cond_wire576_in =
  _guard22949 ? cond576_out :
  _guard22950 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire584_in =
  _guard22953 ? cond584_out :
  _guard22954 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire602_in =
  _guard22955 ? idx_between_14_30_reg_out :
  _guard22958 ? cond602_out :
  1'd0;
assign cond605_write_en = _guard22959;
assign cond605_clk = clk;
assign cond605_reset = reset;
assign cond605_in =
  _guard22960 ? idx_between_11_27_reg_out :
  1'd0;
assign cond_wire605_in =
  _guard22961 ? idx_between_11_27_reg_out :
  _guard22964 ? cond605_out :
  1'd0;
assign cond620_write_en = _guard22965;
assign cond620_clk = clk;
assign cond620_reset = reset;
assign cond620_in =
  _guard22966 ? idx_between_15_19_reg_out :
  1'd0;
assign cond_wire633_in =
  _guard22967 ? idx_between_18_34_reg_out :
  _guard22970 ? cond633_out :
  1'd0;
assign cond635_write_en = _guard22971;
assign cond635_clk = clk;
assign cond635_reset = reset;
assign cond635_in =
  _guard22972 ? idx_between_38_39_reg_out :
  1'd0;
assign cond639_write_en = _guard22973;
assign cond639_clk = clk;
assign cond639_reset = reset;
assign cond639_in =
  _guard22974 ? idx_between_39_40_reg_out :
  1'd0;
assign cond646_write_en = _guard22975;
assign cond646_clk = clk;
assign cond646_reset = reset;
assign cond646_in =
  _guard22976 ? idx_between_25_41_reg_out :
  1'd0;
assign cond_wire647_in =
  _guard22979 ? cond647_out :
  _guard22980 ? idx_between_41_42_reg_out :
  1'd0;
assign cond649_write_en = _guard22981;
assign cond649_clk = clk;
assign cond649_reset = reset;
assign cond649_in =
  _guard22982 ? idx_between_22_38_reg_out :
  1'd0;
assign cond654_write_en = _guard22983;
assign cond654_clk = clk;
assign cond654_reset = reset;
assign cond654_in =
  _guard22984 ? idx_between_27_43_reg_out :
  1'd0;
assign cond658_write_en = _guard22985;
assign cond658_clk = clk;
assign cond658_reset = reset;
assign cond658_in =
  _guard22986 ? idx_between_28_44_reg_out :
  1'd0;
assign cond690_write_en = _guard22987;
assign cond690_clk = clk;
assign cond690_reset = reset;
assign cond690_in =
  _guard22988 ? idx_between_17_33_reg_out :
  1'd0;
assign cond_wire702_in =
  _guard22989 ? idx_between_20_36_reg_out :
  _guard22992 ? cond702_out :
  1'd0;
assign cond_wire704_in =
  _guard22995 ? cond704_out :
  _guard22996 ? idx_between_40_41_reg_out :
  1'd0;
assign cond_wire707_in =
  _guard22999 ? cond707_out :
  _guard23000 ? idx_between_25_41_reg_out :
  1'd0;
assign cond712_write_en = _guard23001;
assign cond712_clk = clk;
assign cond712_reset = reset;
assign cond712_in =
  _guard23002 ? idx_between_42_43_reg_out :
  1'd0;
assign cond_wire727_in =
  _guard23003 ? idx_between_30_46_reg_out :
  _guard23006 ? cond727_out :
  1'd0;
assign cond_wire728_in =
  _guard23009 ? cond728_out :
  _guard23010 ? idx_between_46_47_reg_out :
  1'd0;
assign cond730_write_en = _guard23011;
assign cond730_clk = clk;
assign cond730_reset = reset;
assign cond730_in =
  _guard23012 ? idx_between_12_16_reg_out :
  1'd0;
assign cond731_write_en = _guard23013;
assign cond731_clk = clk;
assign cond731_reset = reset;
assign cond731_in =
  _guard23014 ? idx_between_12_28_reg_out :
  1'd0;
assign cond732_write_en = _guard23015;
assign cond732_clk = clk;
assign cond732_reset = reset;
assign cond732_in =
  _guard23016 ? idx_between_16_32_reg_out :
  1'd0;
assign cond_wire736_in =
  _guard23017 ? idx_between_17_33_reg_out :
  _guard23020 ? cond736_out :
  1'd0;
assign cond_wire744_in =
  _guard23023 ? cond744_out :
  _guard23024 ? idx_between_19_35_reg_out :
  1'd0;
assign cond750_write_en = _guard23025;
assign cond750_clk = clk;
assign cond750_reset = reset;
assign cond750_in =
  _guard23026 ? idx_between_17_21_reg_out :
  1'd0;
assign cond756_write_en = _guard23027;
assign cond756_clk = clk;
assign cond756_reset = reset;
assign cond756_in =
  _guard23028 ? idx_between_22_38_reg_out :
  1'd0;
assign cond761_write_en = _guard23029;
assign cond761_clk = clk;
assign cond761_reset = reset;
assign cond761_in =
  _guard23030 ? idx_between_39_40_reg_out :
  1'd0;
assign cond_wire770_in =
  _guard23033 ? cond770_out :
  _guard23034 ? idx_between_22_26_reg_out :
  1'd0;
assign cond_wire777_in =
  _guard23035 ? idx_between_43_44_reg_out :
  _guard23038 ? cond777_out :
  1'd0;
assign cond_wire779_in =
  _guard23041 ? cond779_out :
  _guard23042 ? idx_between_24_40_reg_out :
  1'd0;
assign cond_wire789_in =
  _guard23045 ? cond789_out :
  _guard23046 ? idx_between_46_47_reg_out :
  1'd0;
assign cond_wire790_in =
  _guard23049 ? cond790_out :
  _guard23050 ? idx_between_27_31_reg_out :
  1'd0;
assign cond802_write_en = _guard23051;
assign cond802_clk = clk;
assign cond802_reset = reset;
assign cond802_in =
  _guard23052 ? idx_between_34_35_reg_out :
  1'd0;
assign cond807_write_en = _guard23053;
assign cond807_clk = clk;
assign cond807_reset = reset;
assign cond807_in =
  _guard23054 ? idx_between_16_20_reg_out :
  1'd0;
assign cond_wire809_in =
  _guard23055 ? idx_between_20_36_reg_out :
  _guard23058 ? cond809_out :
  1'd0;
assign cond818_write_en = _guard23059;
assign cond818_clk = clk;
assign cond818_reset = reset;
assign cond818_in =
  _guard23060 ? idx_between_38_39_reg_out :
  1'd0;
assign cond_wire828_in =
  _guard23063 ? cond828_out :
  _guard23064 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire835_in =
  _guard23067 ? cond835_out :
  _guard23068 ? idx_between_23_27_reg_out :
  1'd0;
assign cond_wire847_in =
  _guard23069 ? idx_between_26_30_reg_out :
  _guard23072 ? cond847_out :
  1'd0;
assign cond848_write_en = _guard23073;
assign cond848_clk = clk;
assign cond848_reset = reset;
assign cond848_in =
  _guard23074 ? idx_between_26_42_reg_out :
  1'd0;
assign cond_wire861_in =
  _guard23077 ? cond861_out :
  _guard23078 ? idx_between_14_30_reg_out :
  1'd0;
assign cond_wire913_in =
  _guard23079 ? idx_between_27_43_reg_out :
  _guard23082 ? cond913_out :
  1'd0;
assign cond914_write_en = _guard23083;
assign cond914_clk = clk;
assign cond914_reset = reset;
assign cond914_in =
  _guard23084 ? idx_between_31_47_reg_out :
  1'd0;
assign cond915_write_en = _guard23085;
assign cond915_clk = clk;
assign cond915_reset = reset;
assign cond915_in =
  _guard23086 ? idx_between_47_48_reg_out :
  1'd0;
assign cond928_write_en = _guard23087;
assign cond928_clk = clk;
assign cond928_reset = reset;
assign cond928_in =
  _guard23088 ? idx_between_35_36_reg_out :
  1'd0;
assign cond935_write_en = _guard23089;
assign cond935_clk = clk;
assign cond935_reset = reset;
assign cond935_in =
  _guard23090 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire938_in =
  _guard23091 ? idx_between_18_34_reg_out :
  _guard23094 ? cond938_out :
  1'd0;
assign cond_wire940_in =
  _guard23097 ? cond940_out :
  _guard23098 ? idx_between_38_39_reg_out :
  1'd0;
assign cond_wire942_in =
  _guard23101 ? cond942_out :
  _guard23102 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire944_in =
  _guard23105 ? cond944_out :
  _guard23106 ? idx_between_39_40_reg_out :
  1'd0;
assign cond951_write_en = _guard23107;
assign cond951_clk = clk;
assign cond951_reset = reset;
assign cond951_in =
  _guard23108 ? idx_between_25_41_reg_out :
  1'd0;
assign cond_wire957_in =
  _guard23111 ? cond957_out :
  _guard23112 ? idx_between_23_27_reg_out :
  1'd0;
assign cond959_write_en = _guard23113;
assign cond959_clk = clk;
assign cond959_reset = reset;
assign cond959_in =
  _guard23114 ? idx_between_27_43_reg_out :
  1'd0;
assign cond964_write_en = _guard23115;
assign cond964_clk = clk;
assign cond964_reset = reset;
assign cond964_in =
  _guard23116 ? idx_between_44_45_reg_out :
  1'd0;
assign cond965_write_en = _guard23117;
assign cond965_clk = clk;
assign cond965_reset = reset;
assign cond965_in =
  _guard23118 ? idx_between_25_29_reg_out :
  1'd0;
assign cond_wire966_in =
  _guard23121 ? cond966_out :
  _guard23122 ? idx_between_25_41_reg_out :
  1'd0;
assign cond978_write_en = _guard23123;
assign cond978_clk = clk;
assign cond978_reset = reset;
assign cond978_in =
  _guard23124 ? idx_between_28_44_reg_out :
  1'd0;
assign cond_wire981_in =
  _guard23127 ? cond981_out :
  _guard23128 ? idx_between_29_33_reg_out :
  1'd0;
assign cond_wire982_in =
  _guard23129 ? idx_between_29_45_reg_out :
  _guard23132 ? cond982_out :
  1'd0;
assign cond_wire986_in =
  _guard23133 ? idx_between_30_46_reg_out :
  _guard23136 ? cond986_out :
  1'd0;
assign cond988_write_en = _guard23137;
assign cond988_clk = clk;
assign cond988_reset = reset;
assign cond988_in =
  _guard23138 ? idx_between_50_51_reg_out :
  1'd0;
assign cond_wire991_in =
  _guard23139 ? idx_between_16_32_reg_out :
  _guard23142 ? cond991_out :
  1'd0;
assign cond1015_write_en = _guard23143;
assign cond1015_clk = clk;
assign cond1015_reset = reset;
assign cond1015_in =
  _guard23144 ? idx_between_22_38_reg_out :
  1'd0;
assign cond1028_write_en = _guard23145;
assign cond1028_clk = clk;
assign cond1028_reset = reset;
assign cond1028_in =
  _guard23146 ? idx_between_29_45_reg_out :
  1'd0;
assign cond1045_write_en = _guard23147;
assign cond1045_clk = clk;
assign cond1045_reset = reset;
assign cond1045_in =
  _guard23148 ? idx_between_49_50_reg_out :
  1'd0;
assign cond_wire1050_in =
  _guard23149 ? idx_between_31_35_reg_out :
  _guard23152 ? cond1050_out :
  1'd0;
assign top_0_0_write_en = _guard23155;
assign top_0_0_clk = clk;
assign top_0_0_reset = reset;
assign top_0_0_in = t0_read_data;
assign top_0_5_write_en = _guard23161;
assign top_0_5_clk = clk;
assign top_0_5_reset = reset;
assign top_0_5_in = t5_read_data;
assign top_0_8_write_en = _guard23167;
assign top_0_8_clk = clk;
assign top_0_8_reset = reset;
assign top_0_8_in = t8_read_data;
assign pe_1_1_mul_ready =
  _guard23173 ? 1'd1 :
  _guard23176 ? 1'd0 :
  1'd0;
assign pe_1_1_clk = clk;
assign pe_1_1_top =
  _guard23189 ? top_1_1_out :
  32'd0;
assign pe_1_1_left =
  _guard23202 ? left_1_1_out :
  32'd0;
assign pe_1_1_reset = reset;
assign pe_1_1_go = _guard23215;
assign top_1_9_write_en = _guard23218;
assign top_1_9_clk = clk;
assign top_1_9_reset = reset;
assign top_1_9_in = top_0_9_out;
assign pe_1_13_mul_ready =
  _guard23224 ? 1'd1 :
  _guard23227 ? 1'd0 :
  1'd0;
assign pe_1_13_clk = clk;
assign pe_1_13_top =
  _guard23240 ? top_1_13_out :
  32'd0;
assign pe_1_13_left =
  _guard23253 ? left_1_13_out :
  32'd0;
assign pe_1_13_reset = reset;
assign pe_1_13_go = _guard23266;
assign top_2_7_write_en = _guard23269;
assign top_2_7_clk = clk;
assign top_2_7_reset = reset;
assign top_2_7_in = top_1_7_out;
assign left_2_11_write_en = _guard23275;
assign left_2_11_clk = clk;
assign left_2_11_reset = reset;
assign left_2_11_in = left_2_10_out;
assign top_2_14_write_en = _guard23281;
assign top_2_14_clk = clk;
assign top_2_14_reset = reset;
assign top_2_14_in = top_1_14_out;
assign left_2_14_write_en = _guard23287;
assign left_2_14_clk = clk;
assign left_2_14_reset = reset;
assign left_2_14_in = left_2_13_out;
assign left_4_11_write_en = _guard23293;
assign left_4_11_clk = clk;
assign left_4_11_reset = reset;
assign left_4_11_in = left_4_10_out;
assign left_5_2_write_en = _guard23299;
assign left_5_2_clk = clk;
assign left_5_2_reset = reset;
assign left_5_2_in = left_5_1_out;
assign top_5_7_write_en = _guard23305;
assign top_5_7_clk = clk;
assign top_5_7_reset = reset;
assign top_5_7_in = top_4_7_out;
assign left_5_7_write_en = _guard23311;
assign left_5_7_clk = clk;
assign left_5_7_reset = reset;
assign left_5_7_in = left_5_6_out;
assign left_6_0_write_en = _guard23317;
assign left_6_0_clk = clk;
assign left_6_0_reset = reset;
assign left_6_0_in = l6_read_data;
assign pe_6_8_mul_ready =
  _guard23323 ? 1'd1 :
  _guard23326 ? 1'd0 :
  1'd0;
assign pe_6_8_clk = clk;
assign pe_6_8_top =
  _guard23339 ? top_6_8_out :
  32'd0;
assign pe_6_8_left =
  _guard23352 ? left_6_8_out :
  32'd0;
assign pe_6_8_reset = reset;
assign pe_6_8_go = _guard23365;
assign top_7_1_write_en = _guard23368;
assign top_7_1_clk = clk;
assign top_7_1_reset = reset;
assign top_7_1_in = top_6_1_out;
assign pe_7_8_mul_ready =
  _guard23374 ? 1'd1 :
  _guard23377 ? 1'd0 :
  1'd0;
assign pe_7_8_clk = clk;
assign pe_7_8_top =
  _guard23390 ? top_7_8_out :
  32'd0;
assign pe_7_8_left =
  _guard23403 ? left_7_8_out :
  32'd0;
assign pe_7_8_reset = reset;
assign pe_7_8_go = _guard23416;
assign pe_7_11_mul_ready =
  _guard23419 ? 1'd1 :
  _guard23422 ? 1'd0 :
  1'd0;
assign pe_7_11_clk = clk;
assign pe_7_11_top =
  _guard23435 ? top_7_11_out :
  32'd0;
assign pe_7_11_left =
  _guard23448 ? left_7_11_out :
  32'd0;
assign pe_7_11_reset = reset;
assign pe_7_11_go = _guard23461;
assign pe_7_13_mul_ready =
  _guard23464 ? 1'd1 :
  _guard23467 ? 1'd0 :
  1'd0;
assign pe_7_13_clk = clk;
assign pe_7_13_top =
  _guard23480 ? top_7_13_out :
  32'd0;
assign pe_7_13_left =
  _guard23493 ? left_7_13_out :
  32'd0;
assign pe_7_13_reset = reset;
assign pe_7_13_go = _guard23506;
assign top_7_13_write_en = _guard23509;
assign top_7_13_clk = clk;
assign top_7_13_reset = reset;
assign top_7_13_in = top_6_13_out;
assign left_7_15_write_en = _guard23515;
assign left_7_15_clk = clk;
assign left_7_15_reset = reset;
assign left_7_15_in = left_7_14_out;
assign top_8_5_write_en = _guard23521;
assign top_8_5_clk = clk;
assign top_8_5_reset = reset;
assign top_8_5_in = top_7_5_out;
assign top_8_9_write_en = _guard23527;
assign top_8_9_clk = clk;
assign top_8_9_reset = reset;
assign top_8_9_in = top_7_9_out;
assign pe_9_2_mul_ready =
  _guard23533 ? 1'd1 :
  _guard23536 ? 1'd0 :
  1'd0;
assign pe_9_2_clk = clk;
assign pe_9_2_top =
  _guard23549 ? top_9_2_out :
  32'd0;
assign pe_9_2_left =
  _guard23562 ? left_9_2_out :
  32'd0;
assign pe_9_2_reset = reset;
assign pe_9_2_go = _guard23575;
assign left_9_3_write_en = _guard23578;
assign left_9_3_clk = clk;
assign left_9_3_reset = reset;
assign left_9_3_in = left_9_2_out;
assign top_9_7_write_en = _guard23584;
assign top_9_7_clk = clk;
assign top_9_7_reset = reset;
assign top_9_7_in = top_8_7_out;
assign top_9_10_write_en = _guard23590;
assign top_9_10_clk = clk;
assign top_9_10_reset = reset;
assign top_9_10_in = top_8_10_out;
assign top_9_13_write_en = _guard23596;
assign top_9_13_clk = clk;
assign top_9_13_reset = reset;
assign top_9_13_in = top_8_13_out;
assign pe_10_1_mul_ready =
  _guard23602 ? 1'd1 :
  _guard23605 ? 1'd0 :
  1'd0;
assign pe_10_1_clk = clk;
assign pe_10_1_top =
  _guard23618 ? top_10_1_out :
  32'd0;
assign pe_10_1_left =
  _guard23631 ? left_10_1_out :
  32'd0;
assign pe_10_1_reset = reset;
assign pe_10_1_go = _guard23644;
assign top_10_3_write_en = _guard23647;
assign top_10_3_clk = clk;
assign top_10_3_reset = reset;
assign top_10_3_in = top_9_3_out;
assign pe_10_6_mul_ready =
  _guard23653 ? 1'd1 :
  _guard23656 ? 1'd0 :
  1'd0;
assign pe_10_6_clk = clk;
assign pe_10_6_top =
  _guard23669 ? top_10_6_out :
  32'd0;
assign pe_10_6_left =
  _guard23682 ? left_10_6_out :
  32'd0;
assign pe_10_6_reset = reset;
assign pe_10_6_go = _guard23695;
assign top_10_12_write_en = _guard23698;
assign top_10_12_clk = clk;
assign top_10_12_reset = reset;
assign top_10_12_in = top_9_12_out;
assign left_11_7_write_en = _guard23704;
assign left_11_7_clk = clk;
assign left_11_7_reset = reset;
assign left_11_7_in = left_11_6_out;
assign top_11_12_write_en = _guard23710;
assign top_11_12_clk = clk;
assign top_11_12_reset = reset;
assign top_11_12_in = top_10_12_out;
assign left_11_13_write_en = _guard23716;
assign left_11_13_clk = clk;
assign left_11_13_reset = reset;
assign left_11_13_in = left_11_12_out;
assign pe_12_0_mul_ready =
  _guard23722 ? 1'd1 :
  _guard23725 ? 1'd0 :
  1'd0;
assign pe_12_0_clk = clk;
assign pe_12_0_top =
  _guard23738 ? top_12_0_out :
  32'd0;
assign pe_12_0_left =
  _guard23751 ? left_12_0_out :
  32'd0;
assign pe_12_0_reset = reset;
assign pe_12_0_go = _guard23764;
assign top_12_4_write_en = _guard23767;
assign top_12_4_clk = clk;
assign top_12_4_reset = reset;
assign top_12_4_in = top_11_4_out;
assign left_12_12_write_en = _guard23773;
assign left_12_12_clk = clk;
assign left_12_12_reset = reset;
assign left_12_12_in = left_12_11_out;
assign left_13_5_write_en = _guard23779;
assign left_13_5_clk = clk;
assign left_13_5_reset = reset;
assign left_13_5_in = left_13_4_out;
assign pe_13_15_mul_ready =
  _guard23785 ? 1'd1 :
  _guard23788 ? 1'd0 :
  1'd0;
assign pe_13_15_clk = clk;
assign pe_13_15_top =
  _guard23801 ? top_13_15_out :
  32'd0;
assign pe_13_15_left =
  _guard23814 ? left_13_15_out :
  32'd0;
assign pe_13_15_reset = reset;
assign pe_13_15_go = _guard23827;
assign top_14_1_write_en = _guard23830;
assign top_14_1_clk = clk;
assign top_14_1_reset = reset;
assign top_14_1_in = top_13_1_out;
assign pe_14_2_mul_ready =
  _guard23836 ? 1'd1 :
  _guard23839 ? 1'd0 :
  1'd0;
assign pe_14_2_clk = clk;
assign pe_14_2_top =
  _guard23852 ? top_14_2_out :
  32'd0;
assign pe_14_2_left =
  _guard23865 ? left_14_2_out :
  32'd0;
assign pe_14_2_reset = reset;
assign pe_14_2_go = _guard23878;
assign left_14_2_write_en = _guard23881;
assign left_14_2_clk = clk;
assign left_14_2_reset = reset;
assign left_14_2_in = left_14_1_out;
assign left_14_5_write_en = _guard23887;
assign left_14_5_clk = clk;
assign left_14_5_reset = reset;
assign left_14_5_in = left_14_4_out;
assign left_14_10_write_en = _guard23893;
assign left_14_10_clk = clk;
assign left_14_10_reset = reset;
assign left_14_10_in = left_14_9_out;
assign pe_15_1_mul_ready =
  _guard23899 ? 1'd1 :
  _guard23902 ? 1'd0 :
  1'd0;
assign pe_15_1_clk = clk;
assign pe_15_1_top =
  _guard23915 ? top_15_1_out :
  32'd0;
assign pe_15_1_left =
  _guard23928 ? left_15_1_out :
  32'd0;
assign pe_15_1_reset = reset;
assign pe_15_1_go = _guard23941;
assign pe_15_5_mul_ready =
  _guard23944 ? 1'd1 :
  _guard23947 ? 1'd0 :
  1'd0;
assign pe_15_5_clk = clk;
assign pe_15_5_top =
  _guard23960 ? top_15_5_out :
  32'd0;
assign pe_15_5_left =
  _guard23973 ? left_15_5_out :
  32'd0;
assign pe_15_5_reset = reset;
assign pe_15_5_go = _guard23986;
assign pe_15_10_mul_ready =
  _guard23989 ? 1'd1 :
  _guard23992 ? 1'd0 :
  1'd0;
assign pe_15_10_clk = clk;
assign pe_15_10_top =
  _guard24005 ? top_15_10_out :
  32'd0;
assign pe_15_10_left =
  _guard24018 ? left_15_10_out :
  32'd0;
assign pe_15_10_reset = reset;
assign pe_15_10_go = _guard24031;
assign top_15_13_write_en = _guard24034;
assign top_15_13_clk = clk;
assign top_15_13_reset = reset;
assign top_15_13_in = top_14_13_out;
assign top_15_15_write_en = _guard24040;
assign top_15_15_clk = clk;
assign top_15_15_reset = reset;
assign top_15_15_in = top_14_15_out;
assign left_15_15_write_en = _guard24046;
assign left_15_15_clk = clk;
assign left_15_15_reset = reset;
assign left_15_15_in = left_15_14_out;
assign l9_add_left = 5'd1;
assign l9_add_right = l9_idx_out;
assign idx_between_26_30_reg_write_en = _guard24060;
assign idx_between_26_30_reg_clk = clk;
assign idx_between_26_30_reg_reset = reset;
assign idx_between_26_30_reg_in =
  _guard24061 ? idx_between_26_30_comb_out :
  _guard24064 ? 1'd0 :
  'x;
assign idx_between_25_41_reg_write_en = _guard24069;
assign idx_between_25_41_reg_clk = clk;
assign idx_between_25_41_reg_reset = reset;
assign idx_between_25_41_reg_in =
  _guard24070 ? idx_between_25_41_comb_out :
  _guard24073 ? 1'd0 :
  'x;
assign index_ge_35_left = idx_add_out;
assign index_ge_35_right = 6'd35;
assign index_ge_13_left = idx_add_out;
assign index_ge_13_right = 6'd13;
assign index_lt_28_left = idx_add_out;
assign index_lt_28_right = 6'd28;
assign idx_between_42_43_comb_left = index_ge_42_out;
assign idx_between_42_43_comb_right = index_lt_43_out;
assign idx_between_31_35_comb_left = index_ge_31_out;
assign idx_between_31_35_comb_right = index_lt_35_out;
assign idx_between_1_5_comb_left = index_ge_1_out;
assign idx_between_1_5_comb_right = index_lt_5_out;
assign idx_between_34_50_reg_write_en = _guard24090;
assign idx_between_34_50_reg_clk = clk;
assign idx_between_34_50_reg_reset = reset;
assign idx_between_34_50_reg_in =
  _guard24091 ? idx_between_34_50_comb_out :
  _guard24094 ? 1'd0 :
  'x;
assign idx_between_8_24_comb_left = index_ge_8_out;
assign idx_between_8_24_comb_right = index_lt_24_out;
assign index_lt_18_left = idx_add_out;
assign index_lt_18_right = 6'd18;
assign idx_between_10_14_reg_write_en = _guard24103;
assign idx_between_10_14_reg_clk = clk;
assign idx_between_10_14_reg_reset = reset;
assign idx_between_10_14_reg_in =
  _guard24104 ? idx_between_10_14_comb_out :
  _guard24107 ? 1'd0 :
  'x;
assign idx_between_28_29_reg_write_en = _guard24112;
assign idx_between_28_29_reg_clk = clk;
assign idx_between_28_29_reg_reset = reset;
assign idx_between_28_29_reg_in =
  _guard24113 ? idx_between_28_29_comb_out :
  _guard24116 ? 1'd0 :
  'x;
assign idx_between_15_31_reg_write_en = _guard24121;
assign idx_between_15_31_reg_clk = clk;
assign idx_between_15_31_reg_reset = reset;
assign idx_between_15_31_reg_in =
  _guard24124 ? 1'd0 :
  _guard24125 ? idx_between_15_31_comb_out :
  'x;
assign idx_between_11_15_reg_write_en = _guard24130;
assign idx_between_11_15_reg_clk = clk;
assign idx_between_11_15_reg_reset = reset;
assign idx_between_11_15_reg_in =
  _guard24133 ? 1'd0 :
  _guard24134 ? idx_between_11_15_comb_out :
  'x;
assign idx_between_35_36_comb_left = index_ge_35_out;
assign idx_between_35_36_comb_right = index_lt_36_out;
assign idx_between_8_12_comb_left = index_ge_8_out;
assign idx_between_8_12_comb_right = index_lt_12_out;
assign idx_between_36_37_comb_left = index_ge_36_out;
assign idx_between_36_37_comb_right = index_lt_37_out;
assign idx_between_9_13_reg_write_en = _guard24145;
assign idx_between_9_13_reg_clk = clk;
assign idx_between_9_13_reg_reset = reset;
assign idx_between_9_13_reg_in =
  _guard24146 ? idx_between_9_13_comb_out :
  _guard24149 ? 1'd0 :
  'x;
assign idx_between_28_44_reg_write_en = _guard24154;
assign idx_between_28_44_reg_clk = clk;
assign idx_between_28_44_reg_reset = reset;
assign idx_between_28_44_reg_in =
  _guard24155 ? idx_between_28_44_comb_out :
  _guard24158 ? 1'd0 :
  'x;
assign index_ge_43_left = idx_add_out;
assign index_ge_43_right = 6'd43;
assign idx_between_24_40_comb_left = index_ge_24_out;
assign idx_between_24_40_comb_right = index_lt_40_out;
assign cond_wire1_in =
  _guard24163 ? idx_between_1_17_reg_out :
  _guard24166 ? cond1_out :
  1'd0;
assign cond8_write_en = _guard24167;
assign cond8_clk = clk;
assign cond8_reset = reset;
assign cond8_in =
  _guard24168 ? idx_between_22_23_reg_out :
  1'd0;
assign cond12_write_en = _guard24169;
assign cond12_clk = clk;
assign cond12_reset = reset;
assign cond12_in =
  _guard24170 ? idx_between_7_23_reg_out :
  1'd0;
assign cond28_write_en = _guard24171;
assign cond28_clk = clk;
assign cond28_reset = reset;
assign cond28_in =
  _guard24172 ? idx_between_26_27_reg_out :
  1'd0;
assign cond_wire28_in =
  _guard24173 ? idx_between_26_27_reg_out :
  _guard24176 ? cond28_out :
  1'd0;
assign cond_wire53_in =
  _guard24179 ? cond53_out :
  _guard24180 ? idx_between_31_32_reg_out :
  1'd0;
assign cond55_write_en = _guard24181;
assign cond55_clk = clk;
assign cond55_reset = reset;
assign cond55_in =
  _guard24182 ? idx_between_12_16_reg_out :
  1'd0;
assign cond_wire65_in =
  _guard24185 ? cond65_out :
  _guard24186 ? idx_between_14_18_reg_out :
  1'd0;
assign cond79_write_en = _guard24187;
assign cond79_clk = clk;
assign cond79_reset = reset;
assign cond79_in =
  _guard24188 ? idx_between_1_17_reg_out :
  1'd0;
assign cond_wire84_in =
  _guard24189 ? idx_between_3_7_reg_out :
  _guard24192 ? cond84_out :
  1'd0;
assign cond_wire88_in =
  _guard24193 ? idx_between_4_8_reg_out :
  _guard24196 ? cond88_out :
  1'd0;
assign cond_wire91_in =
  _guard24199 ? cond91_out :
  _guard24200 ? idx_between_24_25_reg_out :
  1'd0;
assign cond_wire109_in =
  _guard24203 ? cond109_out :
  _guard24204 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire115_in =
  _guard24207 ? cond115_out :
  _guard24208 ? idx_between_30_31_reg_out :
  1'd0;
assign cond117_write_en = _guard24209;
assign cond117_clk = clk;
assign cond117_reset = reset;
assign cond117_in =
  _guard24210 ? idx_between_11_27_reg_out :
  1'd0;
assign cond_wire119_in =
  _guard24211 ? idx_between_31_32_reg_out :
  _guard24214 ? cond119_out :
  1'd0;
assign cond126_write_en = _guard24215;
assign cond126_clk = clk;
assign cond126_reset = reset;
assign cond126_in =
  _guard24216 ? idx_between_17_33_reg_out :
  1'd0;
assign cond135_write_en = _guard24217;
assign cond135_clk = clk;
assign cond135_reset = reset;
assign cond135_in =
  _guard24218 ? idx_between_35_36_reg_out :
  1'd0;
assign cond_wire141_in =
  _guard24219 ? idx_between_17_33_reg_out :
  _guard24222 ? cond141_out :
  1'd0;
assign cond153_write_en = _guard24223;
assign cond153_clk = clk;
assign cond153_reset = reset;
assign cond153_in =
  _guard24224 ? idx_between_5_9_reg_out :
  1'd0;
assign cond_wire158_in =
  _guard24225 ? idx_between_6_22_reg_out :
  _guard24228 ? cond158_out :
  1'd0;
assign cond_wire159_in =
  _guard24231 ? cond159_out :
  _guard24232 ? idx_between_10_26_reg_out :
  1'd0;
assign cond_wire169_in =
  _guard24235 ? cond169_out :
  _guard24236 ? idx_between_9_13_reg_out :
  1'd0;
assign cond171_write_en = _guard24237;
assign cond171_clk = clk;
assign cond171_reset = reset;
assign cond171_in =
  _guard24238 ? idx_between_13_29_reg_out :
  1'd0;
assign cond186_write_en = _guard24239;
assign cond186_clk = clk;
assign cond186_reset = reset;
assign cond186_in =
  _guard24240 ? idx_between_13_29_reg_out :
  1'd0;
assign cond_wire186_in =
  _guard24241 ? idx_between_13_29_reg_out :
  _guard24244 ? cond186_out :
  1'd0;
assign cond_wire196_in =
  _guard24247 ? cond196_out :
  _guard24248 ? idx_between_35_36_reg_out :
  1'd0;
assign cond213_write_en = _guard24249;
assign cond213_clk = clk;
assign cond213_reset = reset;
assign cond213_in =
  _guard24250 ? idx_between_24_25_reg_out :
  1'd0;
assign cond234_write_en = _guard24251;
assign cond234_clk = clk;
assign cond234_reset = reset;
assign cond234_in =
  _guard24252 ? idx_between_10_14_reg_out :
  1'd0;
assign cond_wire235_in =
  _guard24255 ? cond235_out :
  _guard24256 ? idx_between_10_26_reg_out :
  1'd0;
assign cond246_write_en = _guard24257;
assign cond246_clk = clk;
assign cond246_reset = reset;
assign cond246_in =
  _guard24258 ? idx_between_13_17_reg_out :
  1'd0;
assign cond_wire257_in =
  _guard24261 ? cond257_out :
  _guard24262 ? idx_between_35_36_reg_out :
  1'd0;
assign cond261_write_en = _guard24263;
assign cond261_clk = clk;
assign cond261_reset = reset;
assign cond261_in =
  _guard24264 ? idx_between_36_37_reg_out :
  1'd0;
assign cond_wire274_in =
  _guard24267 ? cond274_out :
  _guard24268 ? idx_between_4_20_reg_out :
  1'd0;
assign cond_wire306_in =
  _guard24269 ? idx_between_32_33_reg_out :
  _guard24272 ? cond306_out :
  1'd0;
assign cond308_write_en = _guard24273;
assign cond308_clk = clk;
assign cond308_reset = reset;
assign cond308_in =
  _guard24274 ? idx_between_13_29_reg_out :
  1'd0;
assign cond_wire309_in =
  _guard24275 ? idx_between_17_33_reg_out :
  _guard24278 ? cond309_out :
  1'd0;
assign cond312_write_en = _guard24279;
assign cond312_clk = clk;
assign cond312_reset = reset;
assign cond312_in =
  _guard24280 ? idx_between_14_30_reg_out :
  1'd0;
assign cond330_write_en = _guard24281;
assign cond330_clk = clk;
assign cond330_reset = reset;
assign cond330_in =
  _guard24282 ? idx_between_38_39_reg_out :
  1'd0;
assign cond338_write_en = _guard24283;
assign cond338_clk = clk;
assign cond338_reset = reset;
assign cond338_in =
  _guard24284 ? idx_between_40_41_reg_out :
  1'd0;
assign cond341_write_en = _guard24285;
assign cond341_clk = clk;
assign cond341_reset = reset;
assign cond341_in =
  _guard24286 ? idx_between_6_22_reg_out :
  1'd0;
assign cond348_write_en = _guard24287;
assign cond348_clk = clk;
assign cond348_reset = reset;
assign cond348_in =
  _guard24288 ? idx_between_8_12_reg_out :
  1'd0;
assign cond351_write_en = _guard24289;
assign cond351_clk = clk;
assign cond351_reset = reset;
assign cond351_in =
  _guard24290 ? idx_between_28_29_reg_out :
  1'd0;
assign cond353_write_en = _guard24291;
assign cond353_clk = clk;
assign cond353_reset = reset;
assign cond353_in =
  _guard24292 ? idx_between_9_25_reg_out :
  1'd0;
assign cond358_write_en = _guard24293;
assign cond358_clk = clk;
assign cond358_reset = reset;
assign cond358_in =
  _guard24294 ? idx_between_14_30_reg_out :
  1'd0;
assign cond359_write_en = _guard24295;
assign cond359_clk = clk;
assign cond359_reset = reset;
assign cond359_in =
  _guard24296 ? idx_between_30_31_reg_out :
  1'd0;
assign cond365_write_en = _guard24297;
assign cond365_clk = clk;
assign cond365_reset = reset;
assign cond365_in =
  _guard24298 ? idx_between_12_28_reg_out :
  1'd0;
assign cond384_write_en = _guard24299;
assign cond384_clk = clk;
assign cond384_reset = reset;
assign cond384_in =
  _guard24300 ? idx_between_17_21_reg_out :
  1'd0;
assign cond_wire389_in =
  _guard24301 ? idx_between_18_34_reg_out :
  _guard24304 ? cond389_out :
  1'd0;
assign cond393_write_en = _guard24305;
assign cond393_clk = clk;
assign cond393_reset = reset;
assign cond393_in =
  _guard24306 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire393_in =
  _guard24307 ? idx_between_19_35_reg_out :
  _guard24310 ? cond393_out :
  1'd0;
assign cond_wire396_in =
  _guard24311 ? idx_between_20_24_reg_out :
  _guard24314 ? cond396_out :
  1'd0;
assign cond_wire426_in =
  _guard24315 ? idx_between_12_28_reg_out :
  _guard24318 ? cond426_out :
  1'd0;
assign cond_wire429_in =
  _guard24321 ? cond429_out :
  _guard24322 ? idx_between_13_17_reg_out :
  1'd0;
assign cond_wire431_in =
  _guard24323 ? idx_between_17_33_reg_out :
  _guard24326 ? cond431_out :
  1'd0;
assign cond_wire437_in =
  _guard24327 ? idx_between_15_19_reg_out :
  _guard24330 ? cond437_out :
  1'd0;
assign cond_wire452_in =
  _guard24333 ? cond452_out :
  _guard24334 ? idx_between_38_39_reg_out :
  1'd0;
assign cond_wire492_in =
  _guard24335 ? idx_between_17_33_reg_out :
  _guard24338 ? cond492_out :
  1'd0;
assign cond_wire500_in =
  _guard24341 ? cond500_out :
  _guard24342 ? idx_between_19_35_reg_out :
  1'd0;
assign cond513_write_en = _guard24343;
assign cond513_clk = clk;
assign cond513_reset = reset;
assign cond513_in =
  _guard24344 ? idx_between_38_39_reg_out :
  1'd0;
assign cond_wire518_in =
  _guard24347 ? cond518_out :
  _guard24348 ? idx_between_20_24_reg_out :
  1'd0;
assign cond521_write_en = _guard24349;
assign cond521_clk = clk;
assign cond521_reset = reset;
assign cond521_in =
  _guard24350 ? idx_between_40_41_reg_out :
  1'd0;
assign cond_wire521_in =
  _guard24351 ? idx_between_40_41_reg_out :
  _guard24354 ? cond521_out :
  1'd0;
assign cond_wire529_in =
  _guard24355 ? idx_between_42_43_reg_out :
  _guard24358 ? cond529_out :
  1'd0;
assign cond535_write_en = _guard24359;
assign cond535_clk = clk;
assign cond535_reset = reset;
assign cond535_in =
  _guard24360 ? idx_between_9_13_reg_out :
  1'd0;
assign cond_wire564_in =
  _guard24361 ? idx_between_16_32_reg_out :
  _guard24364 ? cond564_out :
  1'd0;
assign cond_wire570_in =
  _guard24367 ? cond570_out :
  _guard24368 ? idx_between_37_38_reg_out :
  1'd0;
assign cond580_write_en = _guard24369;
assign cond580_clk = clk;
assign cond580_reset = reset;
assign cond580_in =
  _guard24370 ? idx_between_20_36_reg_out :
  1'd0;
assign cond591_write_en = _guard24371;
assign cond591_clk = clk;
assign cond591_reset = reset;
assign cond591_in =
  _guard24372 ? idx_between_23_27_reg_out :
  1'd0;
assign cond_wire608_in =
  _guard24375 ? cond608_out :
  _guard24376 ? idx_between_12_16_reg_out :
  1'd0;
assign cond611_write_en = _guard24377;
assign cond611_clk = clk;
assign cond611_reset = reset;
assign cond611_in =
  _guard24378 ? idx_between_32_33_reg_out :
  1'd0;
assign cond612_write_en = _guard24379;
assign cond612_clk = clk;
assign cond612_reset = reset;
assign cond612_in =
  _guard24380 ? idx_between_13_17_reg_out :
  1'd0;
assign cond_wire613_in =
  _guard24381 ? idx_between_13_29_reg_out :
  _guard24384 ? cond613_out :
  1'd0;
assign cond_wire624_in =
  _guard24385 ? idx_between_16_20_reg_out :
  _guard24388 ? cond624_out :
  1'd0;
assign cond_wire629_in =
  _guard24389 ? idx_between_17_33_reg_out :
  _guard24392 ? cond629_out :
  1'd0;
assign cond630_write_en = _guard24393;
assign cond630_clk = clk;
assign cond630_reset = reset;
assign cond630_in =
  _guard24394 ? idx_between_21_37_reg_out :
  1'd0;
assign cond645_write_en = _guard24395;
assign cond645_clk = clk;
assign cond645_reset = reset;
assign cond645_in =
  _guard24396 ? idx_between_21_37_reg_out :
  1'd0;
assign cond_wire658_in =
  _guard24399 ? cond658_out :
  _guard24400 ? idx_between_28_44_reg_out :
  1'd0;
assign cond_wire666_in =
  _guard24401 ? idx_between_11_27_reg_out :
  _guard24404 ? cond666_out :
  1'd0;
assign cond_wire675_in =
  _guard24405 ? idx_between_17_33_reg_out :
  _guard24408 ? cond675_out :
  1'd0;
assign cond676_write_en = _guard24409;
assign cond676_clk = clk;
assign cond676_reset = reset;
assign cond676_in =
  _guard24410 ? idx_between_33_34_reg_out :
  1'd0;
assign cond681_write_en = _guard24411;
assign cond681_clk = clk;
assign cond681_reset = reset;
assign cond681_in =
  _guard24412 ? idx_between_15_19_reg_out :
  1'd0;
assign cond_wire701_in =
  _guard24415 ? cond701_out :
  _guard24416 ? idx_between_20_24_reg_out :
  1'd0;
assign cond_wire708_in =
  _guard24419 ? cond708_out :
  _guard24420 ? idx_between_41_42_reg_out :
  1'd0;
assign cond_wire712_in =
  _guard24421 ? idx_between_42_43_reg_out :
  _guard24424 ? cond712_out :
  1'd0;
assign cond717_write_en = _guard24425;
assign cond717_clk = clk;
assign cond717_reset = reset;
assign cond717_in =
  _guard24426 ? idx_between_24_28_reg_out :
  1'd0;
assign cond_wire718_in =
  _guard24429 ? cond718_out :
  _guard24430 ? idx_between_24_40_reg_out :
  1'd0;
assign cond719_write_en = _guard24431;
assign cond719_clk = clk;
assign cond719_reset = reset;
assign cond719_in =
  _guard24432 ? idx_between_28_44_reg_out :
  1'd0;
assign cond721_write_en = _guard24433;
assign cond721_clk = clk;
assign cond721_reset = reset;
assign cond721_in =
  _guard24434 ? idx_between_25_29_reg_out :
  1'd0;
assign cond_wire724_in =
  _guard24435 ? idx_between_45_46_reg_out :
  _guard24438 ? cond724_out :
  1'd0;
assign cond_wire730_in =
  _guard24439 ? idx_between_12_16_reg_out :
  _guard24442 ? cond730_out :
  1'd0;
assign cond_wire732_in =
  _guard24443 ? idx_between_16_32_reg_out :
  _guard24446 ? cond732_out :
  1'd0;
assign cond738_write_en = _guard24447;
assign cond738_clk = clk;
assign cond738_reset = reset;
assign cond738_in =
  _guard24448 ? idx_between_14_18_reg_out :
  1'd0;
assign cond_wire740_in =
  _guard24449 ? idx_between_18_34_reg_out :
  _guard24452 ? cond740_out :
  1'd0;
assign cond_wire746_in =
  _guard24453 ? idx_between_16_20_reg_out :
  _guard24456 ? cond746_out :
  1'd0;
assign cond_wire753_in =
  _guard24459 ? cond753_out :
  _guard24460 ? idx_between_37_38_reg_out :
  1'd0;
assign cond_wire755_in =
  _guard24463 ? cond755_out :
  _guard24464 ? idx_between_18_34_reg_out :
  1'd0;
assign cond757_write_en = _guard24465;
assign cond757_clk = clk;
assign cond757_reset = reset;
assign cond757_in =
  _guard24466 ? idx_between_38_39_reg_out :
  1'd0;
assign cond_wire757_in =
  _guard24469 ? cond757_out :
  _guard24470 ? idx_between_38_39_reg_out :
  1'd0;
assign cond_wire759_in =
  _guard24473 ? cond759_out :
  _guard24474 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire766_in =
  _guard24477 ? cond766_out :
  _guard24478 ? idx_between_21_25_reg_out :
  1'd0;
assign cond_wire775_in =
  _guard24479 ? idx_between_23_39_reg_out :
  _guard24482 ? cond775_out :
  1'd0;
assign cond_wire778_in =
  _guard24485 ? cond778_out :
  _guard24486 ? idx_between_24_28_reg_out :
  1'd0;
assign cond_wire795_in =
  _guard24489 ? cond795_out :
  _guard24490 ? idx_between_13_17_reg_out :
  1'd0;
assign cond_wire804_in =
  _guard24493 ? cond804_out :
  _guard24494 ? idx_between_15_31_reg_out :
  1'd0;
assign cond_wire834_in =
  _guard24495 ? idx_between_42_43_reg_out :
  _guard24498 ? cond834_out :
  1'd0;
assign cond842_write_en = _guard24499;
assign cond842_clk = clk;
assign cond842_reset = reset;
assign cond842_in =
  _guard24500 ? idx_between_44_45_reg_out :
  1'd0;
assign cond843_write_en = _guard24501;
assign cond843_clk = clk;
assign cond843_reset = reset;
assign cond843_in =
  _guard24502 ? idx_between_25_29_reg_out :
  1'd0;
assign cond847_write_en = _guard24503;
assign cond847_clk = clk;
assign cond847_reset = reset;
assign cond847_in =
  _guard24504 ? idx_between_26_30_reg_out :
  1'd0;
assign cond_wire853_in =
  _guard24507 ? cond853_out :
  _guard24508 ? idx_between_31_47_reg_out :
  1'd0;
assign cond855_write_en = _guard24509;
assign cond855_clk = clk;
assign cond855_reset = reset;
assign cond855_in =
  _guard24510 ? idx_between_28_32_reg_out :
  1'd0;
assign cond_wire864_in =
  _guard24511 ? idx_between_15_19_reg_out :
  _guard24514 ? cond864_out :
  1'd0;
assign cond869_write_en = _guard24515;
assign cond869_clk = clk;
assign cond869_reset = reset;
assign cond869_in =
  _guard24516 ? idx_between_16_32_reg_out :
  1'd0;
assign cond875_write_en = _guard24517;
assign cond875_clk = clk;
assign cond875_reset = reset;
assign cond875_in =
  _guard24518 ? idx_between_37_38_reg_out :
  1'd0;
assign cond877_write_en = _guard24519;
assign cond877_clk = clk;
assign cond877_reset = reset;
assign cond877_in =
  _guard24520 ? idx_between_18_34_reg_out :
  1'd0;
assign cond_wire879_in =
  _guard24523 ? cond879_out :
  _guard24524 ? idx_between_38_39_reg_out :
  1'd0;
assign cond881_write_en = _guard24525;
assign cond881_clk = clk;
assign cond881_reset = reset;
assign cond881_in =
  _guard24526 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire882_in =
  _guard24527 ? idx_between_23_39_reg_out :
  _guard24530 ? cond882_out :
  1'd0;
assign cond883_write_en = _guard24531;
assign cond883_clk = clk;
assign cond883_reset = reset;
assign cond883_in =
  _guard24532 ? idx_between_39_40_reg_out :
  1'd0;
assign cond_wire894_in =
  _guard24535 ? cond894_out :
  _guard24536 ? idx_between_26_42_reg_out :
  1'd0;
assign cond900_write_en = _guard24537;
assign cond900_clk = clk;
assign cond900_reset = reset;
assign cond900_in =
  _guard24538 ? idx_between_24_28_reg_out :
  1'd0;
assign cond905_write_en = _guard24539;
assign cond905_clk = clk;
assign cond905_reset = reset;
assign cond905_in =
  _guard24540 ? idx_between_25_41_reg_out :
  1'd0;
assign cond_wire907_in =
  _guard24543 ? cond907_out :
  _guard24544 ? idx_between_45_46_reg_out :
  1'd0;
assign cond_wire914_in =
  _guard24545 ? idx_between_31_47_reg_out :
  _guard24548 ? cond914_out :
  1'd0;
assign cond_wire916_in =
  _guard24549 ? idx_between_28_32_reg_out :
  _guard24552 ? cond916_out :
  1'd0;
assign cond925_write_en = _guard24553;
assign cond925_clk = clk;
assign cond925_reset = reset;
assign cond925_in =
  _guard24554 ? idx_between_15_19_reg_out :
  1'd0;
assign cond_wire929_in =
  _guard24555 ? idx_between_16_20_reg_out :
  _guard24558 ? cond929_out :
  1'd0;
assign cond_wire930_in =
  _guard24559 ? idx_between_16_32_reg_out :
  _guard24562 ? cond930_out :
  1'd0;
assign cond933_write_en = _guard24563;
assign cond933_clk = clk;
assign cond933_reset = reset;
assign cond933_in =
  _guard24564 ? idx_between_17_21_reg_out :
  1'd0;
assign cond948_write_en = _guard24565;
assign cond948_clk = clk;
assign cond948_reset = reset;
assign cond948_in =
  _guard24566 ? idx_between_40_41_reg_out :
  1'd0;
assign cond956_write_en = _guard24567;
assign cond956_clk = clk;
assign cond956_reset = reset;
assign cond956_in =
  _guard24568 ? idx_between_42_43_reg_out :
  1'd0;
assign cond_wire978_in =
  _guard24571 ? cond978_out :
  _guard24572 ? idx_between_28_44_reg_out :
  1'd0;
assign cond983_write_en = _guard24573;
assign cond983_clk = clk;
assign cond983_reset = reset;
assign cond983_in =
  _guard24574 ? idx_between_33_49_reg_out :
  1'd0;
assign cond_wire994_in =
  _guard24575 ? idx_between_17_21_reg_out :
  _guard24578 ? cond994_out :
  1'd0;
assign cond_wire996_in =
  _guard24581 ? cond996_out :
  _guard24582 ? idx_between_21_37_reg_out :
  1'd0;
assign cond1004_write_en = _guard24583;
assign cond1004_clk = clk;
assign cond1004_reset = reset;
assign cond1004_in =
  _guard24584 ? idx_between_23_39_reg_out :
  1'd0;
assign cond1013_write_en = _guard24585;
assign cond1013_clk = clk;
assign cond1013_reset = reset;
assign cond1013_in =
  _guard24586 ? idx_between_41_42_reg_out :
  1'd0;
assign cond1020_write_en = _guard24587;
assign cond1020_clk = clk;
assign cond1020_reset = reset;
assign cond1020_in =
  _guard24588 ? idx_between_27_43_reg_out :
  1'd0;
assign cond1030_write_en = _guard24589;
assign cond1030_clk = clk;
assign cond1030_reset = reset;
assign cond1030_in =
  _guard24590 ? idx_between_26_30_reg_out :
  1'd0;
assign cond1046_write_en = _guard24591;
assign cond1046_clk = clk;
assign cond1046_reset = reset;
assign cond1046_in =
  _guard24592 ? idx_between_30_34_reg_out :
  1'd0;
assign cond1052_write_en = _guard24593;
assign cond1052_clk = clk;
assign cond1052_reset = reset;
assign cond1052_in =
  _guard24594 ? idx_between_51_52_reg_out :
  1'd0;
assign wrapper_early_reset_static_seq_go_in = go;
assign left_0_1_write_en = _guard24597;
assign left_0_1_clk = clk;
assign left_0_1_reset = reset;
assign left_0_1_in = left_0_0_out;
assign top_0_7_write_en = _guard24603;
assign top_0_7_clk = clk;
assign top_0_7_reset = reset;
assign top_0_7_in = t7_read_data;
assign left_0_11_write_en = _guard24609;
assign left_0_11_clk = clk;
assign left_0_11_reset = reset;
assign left_0_11_in = left_0_10_out;
assign pe_0_13_mul_ready =
  _guard24615 ? 1'd1 :
  _guard24618 ? 1'd0 :
  1'd0;
assign pe_0_13_clk = clk;
assign pe_0_13_top =
  _guard24631 ? top_0_13_out :
  32'd0;
assign pe_0_13_left =
  _guard24644 ? left_0_13_out :
  32'd0;
assign pe_0_13_reset = reset;
assign pe_0_13_go = _guard24657;
assign top_0_13_write_en = _guard24660;
assign top_0_13_clk = clk;
assign top_0_13_reset = reset;
assign top_0_13_in = t13_read_data;
assign left_0_15_write_en = _guard24666;
assign left_0_15_clk = clk;
assign left_0_15_reset = reset;
assign left_0_15_in = left_0_14_out;
assign left_1_7_write_en = _guard24672;
assign left_1_7_clk = clk;
assign left_1_7_reset = reset;
assign left_1_7_in = left_1_6_out;
assign pe_1_10_mul_ready =
  _guard24678 ? 1'd1 :
  _guard24681 ? 1'd0 :
  1'd0;
assign pe_1_10_clk = clk;
assign pe_1_10_top =
  _guard24694 ? top_1_10_out :
  32'd0;
assign pe_1_10_left =
  _guard24707 ? left_1_10_out :
  32'd0;
assign pe_1_10_reset = reset;
assign pe_1_10_go = _guard24720;
assign pe_1_14_mul_ready =
  _guard24723 ? 1'd1 :
  _guard24726 ? 1'd0 :
  1'd0;
assign pe_1_14_clk = clk;
assign pe_1_14_top =
  _guard24739 ? top_1_14_out :
  32'd0;
assign pe_1_14_left =
  _guard24752 ? left_1_14_out :
  32'd0;
assign pe_1_14_reset = reset;
assign pe_1_14_go = _guard24765;
assign pe_2_2_mul_ready =
  _guard24768 ? 1'd1 :
  _guard24771 ? 1'd0 :
  1'd0;
assign pe_2_2_clk = clk;
assign pe_2_2_top =
  _guard24784 ? top_2_2_out :
  32'd0;
assign pe_2_2_left =
  _guard24797 ? left_2_2_out :
  32'd0;
assign pe_2_2_reset = reset;
assign pe_2_2_go = _guard24810;
assign pe_2_9_mul_ready =
  _guard24813 ? 1'd1 :
  _guard24816 ? 1'd0 :
  1'd0;
assign pe_2_9_clk = clk;
assign pe_2_9_top =
  _guard24829 ? top_2_9_out :
  32'd0;
assign pe_2_9_left =
  _guard24842 ? left_2_9_out :
  32'd0;
assign pe_2_9_reset = reset;
assign pe_2_9_go = _guard24855;
assign top_2_9_write_en = _guard24858;
assign top_2_9_clk = clk;
assign top_2_9_reset = reset;
assign top_2_9_in = top_1_9_out;
assign pe_2_10_mul_ready =
  _guard24864 ? 1'd1 :
  _guard24867 ? 1'd0 :
  1'd0;
assign pe_2_10_clk = clk;
assign pe_2_10_top =
  _guard24880 ? top_2_10_out :
  32'd0;
assign pe_2_10_left =
  _guard24893 ? left_2_10_out :
  32'd0;
assign pe_2_10_reset = reset;
assign pe_2_10_go = _guard24906;
assign left_2_13_write_en = _guard24909;
assign left_2_13_clk = clk;
assign left_2_13_reset = reset;
assign left_2_13_in = left_2_12_out;
assign pe_4_1_mul_ready =
  _guard24915 ? 1'd1 :
  _guard24918 ? 1'd0 :
  1'd0;
assign pe_4_1_clk = clk;
assign pe_4_1_top =
  _guard24931 ? top_4_1_out :
  32'd0;
assign pe_4_1_left =
  _guard24944 ? left_4_1_out :
  32'd0;
assign pe_4_1_reset = reset;
assign pe_4_1_go = _guard24957;
assign left_4_3_write_en = _guard24960;
assign left_4_3_clk = clk;
assign left_4_3_reset = reset;
assign left_4_3_in = left_4_2_out;
assign top_4_10_write_en = _guard24966;
assign top_4_10_clk = clk;
assign top_4_10_reset = reset;
assign top_4_10_in = top_3_10_out;
assign left_4_12_write_en = _guard24972;
assign left_4_12_clk = clk;
assign left_4_12_reset = reset;
assign left_4_12_in = left_4_11_out;
assign left_4_13_write_en = _guard24978;
assign left_4_13_clk = clk;
assign left_4_13_reset = reset;
assign left_4_13_in = left_4_12_out;
assign top_4_15_write_en = _guard24984;
assign top_4_15_clk = clk;
assign top_4_15_reset = reset;
assign top_4_15_in = top_3_15_out;
assign pe_5_12_mul_ready =
  _guard24990 ? 1'd1 :
  _guard24993 ? 1'd0 :
  1'd0;
assign pe_5_12_clk = clk;
assign pe_5_12_top =
  _guard25006 ? top_5_12_out :
  32'd0;
assign pe_5_12_left =
  _guard25019 ? left_5_12_out :
  32'd0;
assign pe_5_12_reset = reset;
assign pe_5_12_go = _guard25032;
assign left_6_3_write_en = _guard25035;
assign left_6_3_clk = clk;
assign left_6_3_reset = reset;
assign left_6_3_in = left_6_2_out;
assign pe_6_9_mul_ready =
  _guard25041 ? 1'd1 :
  _guard25044 ? 1'd0 :
  1'd0;
assign pe_6_9_clk = clk;
assign pe_6_9_top =
  _guard25057 ? top_6_9_out :
  32'd0;
assign pe_6_9_left =
  _guard25070 ? left_6_9_out :
  32'd0;
assign pe_6_9_reset = reset;
assign pe_6_9_go = _guard25083;
assign top_6_10_write_en = _guard25086;
assign top_6_10_clk = clk;
assign top_6_10_reset = reset;
assign top_6_10_in = top_5_10_out;
assign left_7_11_write_en = _guard25092;
assign left_7_11_clk = clk;
assign left_7_11_reset = reset;
assign left_7_11_in = left_7_10_out;
assign top_7_12_write_en = _guard25098;
assign top_7_12_clk = clk;
assign top_7_12_reset = reset;
assign top_7_12_in = top_6_12_out;
assign top_8_1_write_en = _guard25104;
assign top_8_1_clk = clk;
assign top_8_1_reset = reset;
assign top_8_1_in = top_7_1_out;
assign pe_8_7_mul_ready =
  _guard25110 ? 1'd1 :
  _guard25113 ? 1'd0 :
  1'd0;
assign pe_8_7_clk = clk;
assign pe_8_7_top =
  _guard25126 ? top_8_7_out :
  32'd0;
assign pe_8_7_left =
  _guard25139 ? left_8_7_out :
  32'd0;
assign pe_8_7_reset = reset;
assign pe_8_7_go = _guard25152;
assign pe_8_8_mul_ready =
  _guard25155 ? 1'd1 :
  _guard25158 ? 1'd0 :
  1'd0;
assign pe_8_8_clk = clk;
assign pe_8_8_top =
  _guard25171 ? top_8_8_out :
  32'd0;
assign pe_8_8_left =
  _guard25184 ? left_8_8_out :
  32'd0;
assign pe_8_8_reset = reset;
assign pe_8_8_go = _guard25197;
assign top_9_0_write_en = _guard25200;
assign top_9_0_clk = clk;
assign top_9_0_reset = reset;
assign top_9_0_in = top_8_0_out;
assign left_9_6_write_en = _guard25206;
assign left_9_6_clk = clk;
assign left_9_6_reset = reset;
assign left_9_6_in = left_9_5_out;
assign top_9_8_write_en = _guard25212;
assign top_9_8_clk = clk;
assign top_9_8_reset = reset;
assign top_9_8_in = top_8_8_out;
assign left_10_8_write_en = _guard25218;
assign left_10_8_clk = clk;
assign left_10_8_reset = reset;
assign left_10_8_in = left_10_7_out;
assign left_11_0_write_en = _guard25224;
assign left_11_0_clk = clk;
assign left_11_0_reset = reset;
assign left_11_0_in = l11_read_data;
assign pe_12_2_mul_ready =
  _guard25230 ? 1'd1 :
  _guard25233 ? 1'd0 :
  1'd0;
assign pe_12_2_clk = clk;
assign pe_12_2_top =
  _guard25246 ? top_12_2_out :
  32'd0;
assign pe_12_2_left =
  _guard25259 ? left_12_2_out :
  32'd0;
assign pe_12_2_reset = reset;
assign pe_12_2_go = _guard25272;
assign pe_12_8_mul_ready =
  _guard25275 ? 1'd1 :
  _guard25278 ? 1'd0 :
  1'd0;
assign pe_12_8_clk = clk;
assign pe_12_8_top =
  _guard25291 ? top_12_8_out :
  32'd0;
assign pe_12_8_left =
  _guard25304 ? left_12_8_out :
  32'd0;
assign pe_12_8_reset = reset;
assign pe_12_8_go = _guard25317;
assign top_12_9_write_en = _guard25320;
assign top_12_9_clk = clk;
assign top_12_9_reset = reset;
assign top_12_9_in = top_11_9_out;
assign pe_12_14_mul_ready =
  _guard25326 ? 1'd1 :
  _guard25329 ? 1'd0 :
  1'd0;
assign pe_12_14_clk = clk;
assign pe_12_14_top =
  _guard25342 ? top_12_14_out :
  32'd0;
assign pe_12_14_left =
  _guard25355 ? left_12_14_out :
  32'd0;
assign pe_12_14_reset = reset;
assign pe_12_14_go = _guard25368;
assign pe_13_2_mul_ready =
  _guard25371 ? 1'd1 :
  _guard25374 ? 1'd0 :
  1'd0;
assign pe_13_2_clk = clk;
assign pe_13_2_top =
  _guard25387 ? top_13_2_out :
  32'd0;
assign pe_13_2_left =
  _guard25400 ? left_13_2_out :
  32'd0;
assign pe_13_2_reset = reset;
assign pe_13_2_go = _guard25413;
assign top_13_2_write_en = _guard25416;
assign top_13_2_clk = clk;
assign top_13_2_reset = reset;
assign top_13_2_in = top_12_2_out;
assign left_13_12_write_en = _guard25422;
assign left_13_12_clk = clk;
assign left_13_12_reset = reset;
assign left_13_12_in = left_13_11_out;
assign top_14_10_write_en = _guard25428;
assign top_14_10_clk = clk;
assign top_14_10_reset = reset;
assign top_14_10_in = top_13_10_out;
assign pe_14_11_mul_ready =
  _guard25434 ? 1'd1 :
  _guard25437 ? 1'd0 :
  1'd0;
assign pe_14_11_clk = clk;
assign pe_14_11_top =
  _guard25450 ? top_14_11_out :
  32'd0;
assign pe_14_11_left =
  _guard25463 ? left_14_11_out :
  32'd0;
assign pe_14_11_reset = reset;
assign pe_14_11_go = _guard25476;
assign top_14_13_write_en = _guard25479;
assign top_14_13_clk = clk;
assign top_14_13_reset = reset;
assign top_14_13_in = top_13_13_out;
assign left_15_3_write_en = _guard25485;
assign left_15_3_clk = clk;
assign left_15_3_reset = reset;
assign left_15_3_in = left_15_2_out;
assign pe_15_8_mul_ready =
  _guard25491 ? 1'd1 :
  _guard25494 ? 1'd0 :
  1'd0;
assign pe_15_8_clk = clk;
assign pe_15_8_top =
  _guard25507 ? top_15_8_out :
  32'd0;
assign pe_15_8_left =
  _guard25520 ? left_15_8_out :
  32'd0;
assign pe_15_8_reset = reset;
assign pe_15_8_go = _guard25533;
assign top_15_8_write_en = _guard25536;
assign top_15_8_clk = clk;
assign top_15_8_reset = reset;
assign top_15_8_in = top_14_8_out;
assign left_15_8_write_en = _guard25542;
assign left_15_8_clk = clk;
assign left_15_8_reset = reset;
assign left_15_8_in = left_15_7_out;
assign left_15_12_write_en = _guard25548;
assign left_15_12_clk = clk;
assign left_15_12_reset = reset;
assign left_15_12_in = left_15_11_out;
assign left_15_13_write_en = _guard25554;
assign left_15_13_clk = clk;
assign left_15_13_reset = reset;
assign left_15_13_in = left_15_12_out;
assign t8_add_left = 5'd1;
assign t8_add_right = t8_idx_out;
assign l2_add_left = 5'd1;
assign l2_add_right = l2_idx_out;
assign l5_idx_write_en = _guard25576;
assign l5_idx_clk = clk;
assign l5_idx_reset = reset;
assign l5_idx_in =
  _guard25579 ? 5'd0 :
  _guard25582 ? l5_add_out :
  'x;
assign l6_add_left = 5'd1;
assign l6_add_right = l6_idx_out;
assign l8_idx_write_en = _guard25595;
assign l8_idx_clk = clk;
assign l8_idx_reset = reset;
assign l8_idx_in =
  _guard25598 ? 5'd0 :
  _guard25601 ? l8_add_out :
  'x;
assign index_lt_45_left = idx_add_out;
assign index_lt_45_right = 6'd45;
assign index_lt_26_left = idx_add_out;
assign index_lt_26_right = 6'd26;
assign index_lt_43_left = idx_add_out;
assign index_lt_43_right = 6'd43;
assign index_lt_42_left = idx_add_out;
assign index_lt_42_right = 6'd42;
assign index_ge_41_left = idx_add_out;
assign index_ge_41_right = 6'd41;
assign idx_between_38_39_reg_write_en = _guard25616;
assign idx_between_38_39_reg_clk = clk;
assign idx_between_38_39_reg_reset = reset;
assign idx_between_38_39_reg_in =
  _guard25617 ? idx_between_38_39_comb_out :
  _guard25620 ? 1'd0 :
  'x;
assign index_lt_23_left = idx_add_out;
assign index_lt_23_right = 6'd23;
assign index_lt_25_left = idx_add_out;
assign index_lt_25_right = 6'd25;
assign idx_between_27_31_reg_write_en = _guard25629;
assign idx_between_27_31_reg_clk = clk;
assign idx_between_27_31_reg_reset = reset;
assign idx_between_27_31_reg_in =
  _guard25630 ? idx_between_27_31_comb_out :
  _guard25633 ? 1'd0 :
  'x;
assign index_lt_31_left = idx_add_out;
assign index_lt_31_right = 6'd31;
assign idx_between_4_20_reg_write_en = _guard25640;
assign idx_between_4_20_reg_clk = clk;
assign idx_between_4_20_reg_reset = reset;
assign idx_between_4_20_reg_in =
  _guard25643 ? 1'd0 :
  _guard25644 ? idx_between_4_20_comb_out :
  'x;
assign idx_between_2_6_reg_write_en = _guard25649;
assign idx_between_2_6_reg_clk = clk;
assign idx_between_2_6_reg_reset = reset;
assign idx_between_2_6_reg_in =
  _guard25652 ? 1'd0 :
  _guard25653 ? idx_between_2_6_comb_out :
  'x;
assign idx_between_2_6_comb_left = index_ge_2_out;
assign idx_between_2_6_comb_right = index_lt_6_out;
assign index_lt_14_left = idx_add_out;
assign index_lt_14_right = 6'd14;
assign idx_between_37_38_reg_write_en = _guard25662;
assign idx_between_37_38_reg_clk = clk;
assign idx_between_37_38_reg_reset = reset;
assign idx_between_37_38_reg_in =
  _guard25663 ? idx_between_37_38_comb_out :
  _guard25666 ? 1'd0 :
  'x;
assign cond_wire14_in =
  _guard25667 ? idx_between_3_19_reg_out :
  _guard25670 ? cond14_out :
  1'd0;
assign cond_wire21_in =
  _guard25671 ? idx_between_5_21_reg_out :
  _guard25674 ? cond21_out :
  1'd0;
assign cond38_write_en = _guard25675;
assign cond38_clk = clk;
assign cond38_reset = reset;
assign cond38_in =
  _guard25676 ? idx_between_28_29_reg_out :
  1'd0;
assign cond42_write_en = _guard25677;
assign cond42_clk = clk;
assign cond42_reset = reset;
assign cond42_in =
  _guard25678 ? idx_between_13_29_reg_out :
  1'd0;
assign cond_wire51_in =
  _guard25679 ? idx_between_11_27_reg_out :
  _guard25682 ? cond51_out :
  1'd0;
assign cond59_write_en = _guard25683;
assign cond59_clk = clk;
assign cond59_reset = reset;
assign cond59_in =
  _guard25684 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire78_in =
  _guard25685 ? idx_between_36_37_reg_out :
  _guard25688 ? cond78_out :
  1'd0;
assign cond_wire79_in =
  _guard25689 ? idx_between_1_17_reg_out :
  _guard25692 ? cond79_out :
  1'd0;
assign cond85_write_en = _guard25693;
assign cond85_clk = clk;
assign cond85_reset = reset;
assign cond85_in =
  _guard25694 ? idx_between_3_19_reg_out :
  1'd0;
assign cond_wire102_in =
  _guard25695 ? idx_between_11_27_reg_out :
  _guard25698 ? cond102_out :
  1'd0;
assign cond111_write_en = _guard25699;
assign cond111_clk = clk;
assign cond111_reset = reset;
assign cond111_in =
  _guard25700 ? idx_between_29_30_reg_out :
  1'd0;
assign cond_wire124_in =
  _guard25703 ? cond124_out :
  _guard25704 ? idx_between_13_17_reg_out :
  1'd0;
assign cond142_write_en = _guard25705;
assign cond142_clk = clk;
assign cond142_reset = reset;
assign cond142_in =
  _guard25706 ? idx_between_21_37_reg_out :
  1'd0;
assign cond157_write_en = _guard25707;
assign cond157_clk = clk;
assign cond157_reset = reset;
assign cond157_in =
  _guard25708 ? idx_between_6_10_reg_out :
  1'd0;
assign cond_wire166_in =
  _guard25711 ? cond166_out :
  _guard25712 ? idx_between_8_24_reg_out :
  1'd0;
assign cond_wire180_in =
  _guard25715 ? cond180_out :
  _guard25716 ? idx_between_31_32_reg_out :
  1'd0;
assign cond_wire183_in =
  _guard25717 ? idx_between_16_32_reg_out :
  _guard25720 ? cond183_out :
  1'd0;
assign cond_wire188_in =
  _guard25723 ? cond188_out :
  _guard25724 ? idx_between_33_34_reg_out :
  1'd0;
assign cond200_write_en = _guard25725;
assign cond200_clk = clk;
assign cond200_reset = reset;
assign cond200_in =
  _guard25726 ? idx_between_36_37_reg_out :
  1'd0;
assign cond_wire202_in =
  _guard25729 ? cond202_out :
  _guard25730 ? idx_between_17_33_reg_out :
  1'd0;
assign cond_wire211_in =
  _guard25733 ? cond211_out :
  _guard25734 ? idx_between_4_20_reg_out :
  1'd0;
assign cond_wire215_in =
  _guard25737 ? cond215_out :
  _guard25738 ? idx_between_5_21_reg_out :
  1'd0;
assign cond_wire226_in =
  _guard25741 ? cond226_out :
  _guard25742 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire227_in =
  _guard25745 ? cond227_out :
  _guard25746 ? idx_between_8_24_reg_out :
  1'd0;
assign cond253_write_en = _guard25747;
assign cond253_clk = clk;
assign cond253_reset = reset;
assign cond253_in =
  _guard25748 ? idx_between_34_35_reg_out :
  1'd0;
assign cond254_write_en = _guard25749;
assign cond254_clk = clk;
assign cond254_reset = reset;
assign cond254_in =
  _guard25750 ? idx_between_15_19_reg_out :
  1'd0;
assign cond_wire254_in =
  _guard25751 ? idx_between_15_19_reg_out :
  _guard25754 ? cond254_out :
  1'd0;
assign cond_wire269_in =
  _guard25757 ? cond269_out :
  _guard25758 ? idx_between_38_39_reg_out :
  1'd0;
assign cond282_write_en = _guard25759;
assign cond282_clk = clk;
assign cond282_reset = reset;
assign cond282_in =
  _guard25760 ? idx_between_26_27_reg_out :
  1'd0;
assign cond285_write_en = _guard25761;
assign cond285_clk = clk;
assign cond285_reset = reset;
assign cond285_in =
  _guard25762 ? idx_between_11_27_reg_out :
  1'd0;
assign cond_wire292_in =
  _guard25765 ? cond292_out :
  _guard25766 ? idx_between_9_25_reg_out :
  1'd0;
assign cond_wire293_in =
  _guard25767 ? idx_between_13_29_reg_out :
  _guard25770 ? cond293_out :
  1'd0;
assign cond_wire295_in =
  _guard25773 ? cond295_out :
  _guard25774 ? idx_between_10_14_reg_out :
  1'd0;
assign cond298_write_en = _guard25775;
assign cond298_clk = clk;
assign cond298_reset = reset;
assign cond298_in =
  _guard25776 ? idx_between_30_31_reg_out :
  1'd0;
assign cond_wire300_in =
  _guard25777 ? idx_between_11_27_reg_out :
  _guard25780 ? cond300_out :
  1'd0;
assign cond304_write_en = _guard25781;
assign cond304_clk = clk;
assign cond304_reset = reset;
assign cond304_in =
  _guard25782 ? idx_between_12_28_reg_out :
  1'd0;
assign cond_wire315_in =
  _guard25783 ? idx_between_15_19_reg_out :
  _guard25786 ? cond315_out :
  1'd0;
assign cond_wire318_in =
  _guard25787 ? idx_between_35_36_reg_out :
  _guard25790 ? cond318_out :
  1'd0;
assign cond_wire333_in =
  _guard25793 ? cond333_out :
  _guard25794 ? idx_between_23_39_reg_out :
  1'd0;
assign cond334_write_en = _guard25795;
assign cond334_clk = clk;
assign cond334_reset = reset;
assign cond334_in =
  _guard25796 ? idx_between_39_40_reg_out :
  1'd0;
assign cond_wire340_in =
  _guard25799 ? cond340_out :
  _guard25800 ? idx_between_6_10_reg_out :
  1'd0;
assign cond_wire352_in =
  _guard25803 ? cond352_out :
  _guard25804 ? idx_between_9_13_reg_out :
  1'd0;
assign cond_wire355_in =
  _guard25807 ? cond355_out :
  _guard25808 ? idx_between_29_30_reg_out :
  1'd0;
assign cond_wire361_in =
  _guard25809 ? idx_between_11_27_reg_out :
  _guard25812 ? cond361_out :
  1'd0;
assign cond364_write_en = _guard25813;
assign cond364_clk = clk;
assign cond364_reset = reset;
assign cond364_in =
  _guard25814 ? idx_between_12_16_reg_out :
  1'd0;
assign cond366_write_en = _guard25815;
assign cond366_clk = clk;
assign cond366_reset = reset;
assign cond366_in =
  _guard25816 ? idx_between_16_32_reg_out :
  1'd0;
assign cond_wire368_in =
  _guard25819 ? cond368_out :
  _guard25820 ? idx_between_13_17_reg_out :
  1'd0;
assign cond_wire370_in =
  _guard25821 ? idx_between_17_33_reg_out :
  _guard25824 ? cond370_out :
  1'd0;
assign cond_wire381_in =
  _guard25825 ? idx_between_16_32_reg_out :
  _guard25828 ? cond381_out :
  1'd0;
assign cond_wire401_in =
  _guard25829 ? idx_between_21_37_reg_out :
  _guard25832 ? cond401_out :
  1'd0;
assign cond_wire413_in =
  _guard25835 ? cond413_out :
  _guard25836 ? idx_between_9_13_reg_out :
  1'd0;
assign cond_wire417_in =
  _guard25839 ? cond417_out :
  _guard25840 ? idx_between_10_14_reg_out :
  1'd0;
assign cond_wire421_in =
  _guard25843 ? cond421_out :
  _guard25844 ? idx_between_11_15_reg_out :
  1'd0;
assign cond_wire439_in =
  _guard25847 ? cond439_out :
  _guard25848 ? idx_between_19_35_reg_out :
  1'd0;
assign cond_wire444_in =
  _guard25849 ? idx_between_36_37_reg_out :
  _guard25852 ? cond444_out :
  1'd0;
assign cond_wire455_in =
  _guard25855 ? cond455_out :
  _guard25856 ? idx_between_23_39_reg_out :
  1'd0;
assign cond480_write_en = _guard25857;
assign cond480_clk = clk;
assign cond480_reset = reset;
assign cond480_in =
  _guard25858 ? idx_between_14_30_reg_out :
  1'd0;
assign cond_wire485_in =
  _guard25861 ? cond485_out :
  _guard25862 ? idx_between_31_32_reg_out :
  1'd0;
assign cond509_write_en = _guard25863;
assign cond509_clk = clk;
assign cond509_reset = reset;
assign cond509_in =
  _guard25864 ? idx_between_37_38_reg_out :
  1'd0;
assign cond516_write_en = _guard25865;
assign cond516_clk = clk;
assign cond516_reset = reset;
assign cond516_in =
  _guard25866 ? idx_between_23_39_reg_out :
  1'd0;
assign cond517_write_en = _guard25867;
assign cond517_clk = clk;
assign cond517_reset = reset;
assign cond517_in =
  _guard25868 ? idx_between_39_40_reg_out :
  1'd0;
assign cond522_write_en = _guard25869;
assign cond522_clk = clk;
assign cond522_reset = reset;
assign cond522_in =
  _guard25870 ? idx_between_21_25_reg_out :
  1'd0;
assign cond_wire556_in =
  _guard25871 ? idx_between_14_30_reg_out :
  _guard25874 ? cond556_out :
  1'd0;
assign cond574_write_en = _guard25875;
assign cond574_clk = clk;
assign cond574_reset = reset;
assign cond574_in =
  _guard25876 ? idx_between_38_39_reg_out :
  1'd0;
assign cond575_write_en = _guard25877;
assign cond575_clk = clk;
assign cond575_reset = reset;
assign cond575_in =
  _guard25878 ? idx_between_19_23_reg_out :
  1'd0;
assign cond_wire575_in =
  _guard25879 ? idx_between_19_23_reg_out :
  _guard25882 ? cond575_out :
  1'd0;
assign cond577_write_en = _guard25883;
assign cond577_clk = clk;
assign cond577_reset = reset;
assign cond577_in =
  _guard25884 ? idx_between_23_39_reg_out :
  1'd0;
assign cond590_write_en = _guard25885;
assign cond590_clk = clk;
assign cond590_reset = reset;
assign cond590_in =
  _guard25886 ? idx_between_42_43_reg_out :
  1'd0;
assign cond_wire592_in =
  _guard25889 ? cond592_out :
  _guard25890 ? idx_between_23_39_reg_out :
  1'd0;
assign cond595_write_en = _guard25891;
assign cond595_clk = clk;
assign cond595_reset = reset;
assign cond595_in =
  _guard25892 ? idx_between_24_28_reg_out :
  1'd0;
assign cond598_write_en = _guard25893;
assign cond598_clk = clk;
assign cond598_reset = reset;
assign cond598_in =
  _guard25894 ? idx_between_44_45_reg_out :
  1'd0;
assign cond_wire603_in =
  _guard25897 ? cond603_out :
  _guard25898 ? idx_between_30_31_reg_out :
  1'd0;
assign cond616_write_en = _guard25899;
assign cond616_clk = clk;
assign cond616_reset = reset;
assign cond616_in =
  _guard25900 ? idx_between_14_18_reg_out :
  1'd0;
assign cond633_write_en = _guard25901;
assign cond633_clk = clk;
assign cond633_reset = reset;
assign cond633_in =
  _guard25902 ? idx_between_18_34_reg_out :
  1'd0;
assign cond_wire643_in =
  _guard25905 ? cond643_out :
  _guard25906 ? idx_between_40_41_reg_out :
  1'd0;
assign cond_wire665_in =
  _guard25909 ? cond665_out :
  _guard25910 ? idx_between_11_15_reg_out :
  1'd0;
assign cond_wire669_in =
  _guard25913 ? cond669_out :
  _guard25914 ? idx_between_12_16_reg_out :
  1'd0;
assign cond673_write_en = _guard25915;
assign cond673_clk = clk;
assign cond673_reset = reset;
assign cond673_in =
  _guard25916 ? idx_between_13_17_reg_out :
  1'd0;
assign cond_wire682_in =
  _guard25919 ? cond682_out :
  _guard25920 ? idx_between_15_31_reg_out :
  1'd0;
assign cond691_write_en = _guard25921;
assign cond691_clk = clk;
assign cond691_reset = reset;
assign cond691_in =
  _guard25922 ? idx_between_21_37_reg_out :
  1'd0;
assign cond703_write_en = _guard25923;
assign cond703_clk = clk;
assign cond703_reset = reset;
assign cond703_in =
  _guard25924 ? idx_between_24_40_reg_out :
  1'd0;
assign cond_wire706_in =
  _guard25925 ? idx_between_21_37_reg_out :
  _guard25928 ? cond706_out :
  1'd0;
assign cond711_write_en = _guard25929;
assign cond711_clk = clk;
assign cond711_reset = reset;
assign cond711_in =
  _guard25930 ? idx_between_26_42_reg_out :
  1'd0;
assign cond_wire721_in =
  _guard25931 ? idx_between_25_29_reg_out :
  _guard25934 ? cond721_out :
  1'd0;
assign cond_wire722_in =
  _guard25937 ? cond722_out :
  _guard25938 ? idx_between_25_41_reg_out :
  1'd0;
assign cond_wire771_in =
  _guard25941 ? cond771_out :
  _guard25942 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire782_in =
  _guard25945 ? cond782_out :
  _guard25946 ? idx_between_25_29_reg_out :
  1'd0;
assign cond_wire786_in =
  _guard25949 ? cond786_out :
  _guard25950 ? idx_between_26_30_reg_out :
  1'd0;
assign cond_wire793_in =
  _guard25953 ? cond793_out :
  _guard25954 ? idx_between_47_48_reg_out :
  1'd0;
assign cond796_write_en = _guard25955;
assign cond796_clk = clk;
assign cond796_reset = reset;
assign cond796_in =
  _guard25956 ? idx_between_13_29_reg_out :
  1'd0;
assign cond_wire796_in =
  _guard25957 ? idx_between_13_29_reg_out :
  _guard25960 ? cond796_out :
  1'd0;
assign cond801_write_en = _guard25961;
assign cond801_clk = clk;
assign cond801_reset = reset;
assign cond801_in =
  _guard25962 ? idx_between_18_34_reg_out :
  1'd0;
assign cond_wire836_in =
  _guard25963 ? idx_between_23_39_reg_out :
  _guard25966 ? cond836_out :
  1'd0;
assign cond_wire848_in =
  _guard25967 ? idx_between_26_42_reg_out :
  _guard25970 ? cond848_out :
  1'd0;
assign cond_wire849_in =
  _guard25971 ? idx_between_30_46_reg_out :
  _guard25974 ? cond849_out :
  1'd0;
assign cond_wire851_in =
  _guard25977 ? cond851_out :
  _guard25978 ? idx_between_27_31_reg_out :
  1'd0;
assign cond854_write_en = _guard25979;
assign cond854_clk = clk;
assign cond854_reset = reset;
assign cond854_in =
  _guard25980 ? idx_between_47_48_reg_out :
  1'd0;
assign cond_wire855_in =
  _guard25981 ? idx_between_28_32_reg_out :
  _guard25984 ? cond855_out :
  1'd0;
assign cond870_write_en = _guard25985;
assign cond870_clk = clk;
assign cond870_reset = reset;
assign cond870_in =
  _guard25986 ? idx_between_20_36_reg_out :
  1'd0;
assign cond872_write_en = _guard25987;
assign cond872_clk = clk;
assign cond872_reset = reset;
assign cond872_in =
  _guard25988 ? idx_between_17_21_reg_out :
  1'd0;
assign cond_wire887_in =
  _guard25991 ? cond887_out :
  _guard25992 ? idx_between_40_41_reg_out :
  1'd0;
assign cond_wire895_in =
  _guard25993 ? idx_between_42_43_reg_out :
  _guard25996 ? cond895_out :
  1'd0;
assign cond_wire899_in =
  _guard25999 ? cond899_out :
  _guard26000 ? idx_between_43_44_reg_out :
  1'd0;
assign cond920_write_en = _guard26001;
assign cond920_clk = clk;
assign cond920_reset = reset;
assign cond920_in =
  _guard26002 ? idx_between_29_33_reg_out :
  1'd0;
assign cond937_write_en = _guard26003;
assign cond937_clk = clk;
assign cond937_reset = reset;
assign cond937_in =
  _guard26004 ? idx_between_18_22_reg_out :
  1'd0;
assign cond954_write_en = _guard26005;
assign cond954_clk = clk;
assign cond954_reset = reset;
assign cond954_in =
  _guard26006 ? idx_between_22_38_reg_out :
  1'd0;
assign cond_wire967_in =
  _guard26009 ? cond967_out :
  _guard26010 ? idx_between_29_45_reg_out :
  1'd0;
assign cond969_write_en = _guard26011;
assign cond969_clk = clk;
assign cond969_reset = reset;
assign cond969_in =
  _guard26012 ? idx_between_26_30_reg_out :
  1'd0;
assign cond_wire972_in =
  _guard26015 ? cond972_out :
  _guard26016 ? idx_between_46_47_reg_out :
  1'd0;
assign cond_wire974_in =
  _guard26019 ? cond974_out :
  _guard26020 ? idx_between_27_43_reg_out :
  1'd0;
assign cond_wire976_in =
  _guard26023 ? cond976_out :
  _guard26024 ? idx_between_47_48_reg_out :
  1'd0;
assign cond980_write_en = _guard26025;
assign cond980_clk = clk;
assign cond980_reset = reset;
assign cond980_in =
  _guard26026 ? idx_between_48_49_reg_out :
  1'd0;
assign cond982_write_en = _guard26027;
assign cond982_clk = clk;
assign cond982_reset = reset;
assign cond982_in =
  _guard26028 ? idx_between_29_45_reg_out :
  1'd0;
assign cond999_write_en = _guard26029;
assign cond999_clk = clk;
assign cond999_reset = reset;
assign cond999_in =
  _guard26030 ? idx_between_18_34_reg_out :
  1'd0;
assign cond1002_write_en = _guard26031;
assign cond1002_clk = clk;
assign cond1002_reset = reset;
assign cond1002_in =
  _guard26032 ? idx_between_19_23_reg_out :
  1'd0;
assign cond1019_write_en = _guard26033;
assign cond1019_clk = clk;
assign cond1019_reset = reset;
assign cond1019_in =
  _guard26034 ? idx_between_23_39_reg_out :
  1'd0;
assign cond_wire1045_in =
  _guard26035 ? idx_between_49_50_reg_out :
  _guard26038 ? cond1045_out :
  1'd0;
assign cond1048_write_en = _guard26039;
assign cond1048_clk = clk;
assign cond1048_reset = reset;
assign cond1048_in =
  _guard26040 ? idx_between_34_50_reg_out :
  1'd0;
// COMPONENT END: main
endmodule

