
/// This is mostly used for testing the static guarantees currently.
/// A realistic implementation would probably take four cycles.
module pipelined_mult (
    input wire clk,
    input wire reset,
    // inputs
    input wire [31:0] left,
    input wire [31:0] right,
    // The input has been committed
    output wire [31:0] out
);

logic [31:0] lt, rt, buff0, buff1, buff2, tmp_prod;

assign out = buff2;
assign tmp_prod = lt * rt;

always_ff @(posedge clk) begin
    if (reset) begin
        lt <= 0;
        rt <= 0;
        buff0 <= 0;
        buff1 <= 0;
        buff2 <= 0;
    end else begin
        lt <= left;
        rt <= right;
        buff0 <= tmp_prod;
        buff1 <= buff0;
        buff2 <= buff1;
    end
end

endmodule

module bb_pipelined_mult(
	               input wire [31:0] left,
	               input wire [31:0] right,
	               output wire [31:0] out,
	               input wire clk
	               );
`ifdef __ICARUS__
   reg [31:0] reg0;
   reg [31:0] reg1;
   reg [31:0] reg2;
   reg [31:0] reg3;
   always @( posedge clk ) begin
      reg0 <= left * right;
      reg1 <= reg0;
      reg2 <= reg1;
      reg3 <= reg2;
   end
   assign out = reg3;
`elsif VERILATOR
   reg [31:0] reg0;
   reg [31:0] reg1;
   reg [31:0] reg2;
   reg [31:0] reg3;
   always @( posedge clk ) begin
      reg0 <= left * right;
      reg1 <= reg0;
      reg2 <= reg1;
      reg3 <= reg2;
   end
   assign out = reg3;
`else
   // mul_uint32 is a black box module generated by Xilinx's IP Core generator.
   // Generation commands are in the synth.tcl file.
   mul_uint32 mul_uint32 (
                   .A(left),
                   .B(right),
                   .P(out),
                   .CLK(clk)
                   );
`endif
endmodule
/* verilator lint_off MULTITOP */
/// =================== Unsigned, Fixed Point =========================
module std_fp_add #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  assign out = left + right;
endmodule

module std_fp_sub #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module std_fp_mult_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16,
    parameter SIGNED = 0
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    input  logic             go,
    input  logic             clk,
    input  logic             reset,
    output logic [WIDTH-1:0] out,
    output logic             done
);
  logic [WIDTH-1:0]          rtmp;
  logic [WIDTH-1:0]          ltmp;
  logic [(WIDTH << 1) - 1:0] out_tmp;
  // Buffer used to walk through the 3 cycles of the pipeline.
  logic done_buf[1:0];

  assign done = done_buf[1];

  assign out = out_tmp[(WIDTH << 1) - INT_WIDTH - 1 : WIDTH - INT_WIDTH];

  // If the done buffer is completely empty and go is high then execution
  // just started.
  logic start;
  assign start = go;

  // Start sending the done signal.
  always_ff @(posedge clk) begin
    if (start)
      done_buf[0] <= 1;
    else
      done_buf[0] <= 0;
  end

  // Push the done signal through the pipeline.
  always_ff @(posedge clk) begin
    if (go) begin
      done_buf[1] <= done_buf[0];
    end else begin
      done_buf[1] <= 0;
    end
  end

  // Register the inputs
  always_ff @(posedge clk) begin
    if (reset) begin
      rtmp <= 0;
      ltmp <= 0;
    end else if (go) begin
      if (SIGNED) begin
        rtmp <= $signed(right);
        ltmp <= $signed(left);
      end else begin
        rtmp <= right;
        ltmp <= left;
      end
    end else begin
      rtmp <= 0;
      ltmp <= 0;
    end

  end

  // Compute the output and save it into out_tmp
  always_ff @(posedge clk) begin
    if (reset) begin
      out_tmp <= 0;
    end else if (go) begin
      if (SIGNED) begin
        // In the first cycle, this performs an invalid computation because
        // ltmp and rtmp only get their actual values in cycle 1
        out_tmp <= $signed(
          { {WIDTH{ltmp[WIDTH-1]}}, ltmp} *
          { {WIDTH{rtmp[WIDTH-1]}}, rtmp}
        );
      end else begin
        out_tmp <= ltmp * rtmp;
      end
    end else begin
      out_tmp <= out_tmp;
    end
  end
endmodule

/* verilator lint_off WIDTH */
module std_fp_div_pipe #(
  parameter WIDTH = 32,
  parameter INT_WIDTH = 16,
  parameter FRAC_WIDTH = 16
) (
    input  logic             go,
    input  logic             clk,
    input  logic             reset,
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out_remainder,
    output logic [WIDTH-1:0] out_quotient,
    output logic             done
);
    localparam ITERATIONS = WIDTH + FRAC_WIDTH;

    logic [WIDTH-1:0] quotient, quotient_next;
    logic [WIDTH:0] acc, acc_next;
    logic [$clog2(ITERATIONS)-1:0] idx;
    logic start, running, finished, dividend_is_zero;

    assign start = go && !running;
    assign dividend_is_zero = start && left == 0;
    assign finished = idx == ITERATIONS - 1 && running;

    always_ff @(posedge clk) begin
      if (reset || finished || dividend_is_zero)
        running <= 0;
      else if (start)
        running <= 1;
      else
        running <= running;
    end

    always_comb begin
      if (acc >= {1'b0, right}) begin
        acc_next = acc - right;
        {acc_next, quotient_next} = {acc_next[WIDTH-1:0], quotient, 1'b1};
      end else begin
        {acc_next, quotient_next} = {acc, quotient} << 1;
      end
    end

    // `done` signaling
    always_ff @(posedge clk) begin
      if (dividend_is_zero || finished)
        done <= 1;
      else
        done <= 0;
    end

    always_ff @(posedge clk) begin
      if (running)
        idx <= idx + 1;
      else
        idx <= 0;
    end

    always_ff @(posedge clk) begin
      if (reset) begin
        out_quotient <= 0;
        out_remainder <= 0;
      end else if (start) begin
        out_quotient <= 0;
        out_remainder <= left;
      end else if (go == 0) begin
        out_quotient <= out_quotient;
        out_remainder <= out_remainder;
      end else if (dividend_is_zero) begin
        out_quotient <= 0;
        out_remainder <= 0;
      end else if (finished) begin
        out_quotient <= quotient_next;
        out_remainder <= out_remainder;
      end else begin
        out_quotient <= out_quotient;
        if (right <= out_remainder)
          out_remainder <= out_remainder - right;
        else
          out_remainder <= out_remainder;
      end
    end

    always_ff @(posedge clk) begin
      if (reset) begin
        acc <= 0;
        quotient <= 0;
      end else if (start) begin
        {acc, quotient} <= {{WIDTH{1'b0}}, left, 1'b0};
      end else begin
        acc <= acc_next;
        quotient <= quotient_next;
      end
    end
endmodule

module std_fp_gt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic             out
);
  assign out = left > right;
endmodule

/// =================== Signed, Fixed Point =========================
module std_fp_sadd #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left + right);
endmodule

module std_fp_ssub #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);

  assign out = $signed(left - right);
endmodule

module std_fp_smult_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  [WIDTH-1:0]              left,
    input  [WIDTH-1:0]              right,
    input  logic                    reset,
    input  logic                    go,
    input  logic                    clk,
    output logic [WIDTH-1:0]        out,
    output logic                    done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(INT_WIDTH),
    .FRAC_WIDTH(FRAC_WIDTH),
    .SIGNED(1)
  ) comp (
    .clk(clk),
    .done(done),
    .reset(reset),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

module std_fp_sdiv_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input                     clk,
    input                     go,
    input                     reset,
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out_quotient,
    output signed [WIDTH-1:0] out_remainder,
    output logic              done
);

  logic signed [WIDTH-1:0] left_abs, right_abs, comp_out_q, comp_out_r, right_save, out_rem_intermediate;

  // Registers to figure out how to transform outputs.
  logic different_signs, left_sign, right_sign;

  // Latch the value of control registers so that their available after
  // go signal becomes low.
  always_ff @(posedge clk) begin
    if (go) begin
      right_save <= right_abs;
      left_sign <= left[WIDTH-1];
      right_sign <= right[WIDTH-1];
    end else begin
      left_sign <= left_sign;
      right_save <= right_save;
      right_sign <= right_sign;
    end
  end

  assign right_abs = right[WIDTH-1] ? -right : right;
  assign left_abs = left[WIDTH-1] ? -left : left;

  assign different_signs = left_sign ^ right_sign;
  assign out_quotient = different_signs ? -comp_out_q : comp_out_q;

  // Remainder is computed as:
  //  t0 = |left| % |right|
  //  t1 = if left * right < 0 and t0 != 0 then |right| - t0 else t0
  //  rem = if right < 0 then -t1 else t1
  assign out_rem_intermediate = different_signs & |comp_out_r ? $signed(right_save - comp_out_r) : comp_out_r;
  assign out_remainder = right_sign ? -out_rem_intermediate : out_rem_intermediate;

  std_fp_div_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(INT_WIDTH),
    .FRAC_WIDTH(FRAC_WIDTH)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left_abs),
    .right(right_abs),
    .out_quotient(comp_out_q),
    .out_remainder(comp_out_r)
  );
endmodule

module std_fp_sgt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic signed [WIDTH-1:0] left,
    input  logic signed [WIDTH-1:0] right,
    output logic signed             out
);
  assign out = $signed(left > right);
endmodule

module std_fp_slt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
   input logic signed [WIDTH-1:0] left,
   input logic signed [WIDTH-1:0] right,
   output logic signed            out
);
  assign out = $signed(left < right);
endmodule

/// =================== Unsigned, Bitnum =========================
module std_mult_pipe #(
    parameter WIDTH = 32
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    input  logic             reset,
    input  logic             go,
    input  logic             clk,
    output logic [WIDTH-1:0] out,
    output logic             done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(WIDTH),
    .FRAC_WIDTH(0),
    .SIGNED(0)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

module std_div_pipe #(
    parameter WIDTH = 32
) (
    input                    reset,
    input                    clk,
    input                    go,
    input        [WIDTH-1:0] left,
    input        [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out_remainder,
    output logic [WIDTH-1:0] out_quotient,
    output logic             done
);

  logic [WIDTH-1:0] dividend;
  logic [(WIDTH-1)*2:0] divisor;
  logic [WIDTH-1:0] quotient;
  logic [WIDTH-1:0] quotient_msk;
  logic start, running, finished, dividend_is_zero;

  assign start = go && !running;
  assign finished = quotient_msk == 0 && running;
  assign dividend_is_zero = start && left == 0;

  always_ff @(posedge clk) begin
    // Early return if the divisor is zero.
    if (finished || dividend_is_zero)
      done <= 1;
    else
      done <= 0;
  end

  always_ff @(posedge clk) begin
    if (reset || finished || dividend_is_zero)
      running <= 0;
    else if (start)
      running <= 1;
    else
      running <= running;
  end

  // Outputs
  always_ff @(posedge clk) begin
    if (dividend_is_zero || start) begin
      out_quotient <= 0;
      out_remainder <= 0;
    end else if (finished) begin
      out_quotient <= quotient;
      out_remainder <= dividend;
    end else begin
      // Otherwise, explicitly latch the values.
      out_quotient <= out_quotient;
      out_remainder <= out_remainder;
    end
  end

  // Calculate the quotient mask.
  always_ff @(posedge clk) begin
    if (start)
      quotient_msk <= 1 << WIDTH - 1;
    else if (running)
      quotient_msk <= quotient_msk >> 1;
    else
      quotient_msk <= quotient_msk;
  end

  // Calculate the quotient.
  always_ff @(posedge clk) begin
    if (start)
      quotient <= 0;
    else if (divisor <= dividend)
      quotient <= quotient | quotient_msk;
    else
      quotient <= quotient;
  end

  // Calculate the dividend.
  always_ff @(posedge clk) begin
    if (start)
      dividend <= left;
    else if (divisor <= dividend)
      dividend <= dividend - divisor;
    else
      dividend <= dividend;
  end

  always_ff @(posedge clk) begin
    if (start) begin
      divisor <= right << WIDTH - 1;
    end else if (finished) begin
      divisor <= 0;
    end else begin
      divisor <= divisor >> 1;
    end
  end

  // Simulation self test against unsynthesizable implementation.
  `ifdef VERILATOR
    logic [WIDTH-1:0] l, r;
    always_ff @(posedge clk) begin
      if (go) begin
        l <= left;
        r <= right;
      end else begin
        l <= l;
        r <= r;
      end
    end

    always @(posedge clk) begin
      if (done && $unsigned(out_remainder) != $unsigned(l % r))
        $error(
          "\nstd_div_pipe (Remainder): Computed and golden outputs do not match!\n",
          "left: %0d", $unsigned(l),
          "  right: %0d\n", $unsigned(r),
          "expected: %0d", $unsigned(l % r),
          "  computed: %0d", $unsigned(out_remainder)
        );

      if (done && $unsigned(out_quotient) != $unsigned(l / r))
        $error(
          "\nstd_div_pipe (Quotient): Computed and golden outputs do not match!\n",
          "left: %0d", $unsigned(l),
          "  right: %0d\n", $unsigned(r),
          "expected: %0d", $unsigned(l / r),
          "  computed: %0d", $unsigned(out_quotient)
        );
    end
  `endif
endmodule

/// =================== Signed, Bitnum =========================
module std_sadd #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left + right);
endmodule

module std_ssub #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left - right);
endmodule

module std_smult_pipe #(
    parameter WIDTH = 32
) (
    input  logic                    reset,
    input  logic                    go,
    input  logic                    clk,
    input  signed       [WIDTH-1:0] left,
    input  signed       [WIDTH-1:0] right,
    output logic signed [WIDTH-1:0] out,
    output logic                    done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(WIDTH),
    .FRAC_WIDTH(0),
    .SIGNED(1)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

/* verilator lint_off WIDTH */
module std_sdiv_pipe #(
    parameter WIDTH = 32
) (
    input                           reset,
    input                           clk,
    input                           go,
    input  logic signed [WIDTH-1:0] left,
    input  logic signed [WIDTH-1:0] right,
    output logic signed [WIDTH-1:0] out_quotient,
    output logic signed [WIDTH-1:0] out_remainder,
    output logic                    done
);

  logic signed [WIDTH-1:0] left_abs, right_abs, comp_out_q, comp_out_r, right_save, out_rem_intermediate;

  // Registers to figure out how to transform outputs.
  logic different_signs, left_sign, right_sign;

  // Latch the value of control registers so that their available after
  // go signal becomes low.
  always_ff @(posedge clk) begin
    if (go) begin
      right_save <= right_abs;
      left_sign <= left[WIDTH-1];
      right_sign <= right[WIDTH-1];
    end else begin
      left_sign <= left_sign;
      right_save <= right_save;
      right_sign <= right_sign;
    end
  end

  assign right_abs = right[WIDTH-1] ? -right : right;
  assign left_abs = left[WIDTH-1] ? -left : left;

  assign different_signs = left_sign ^ right_sign;
  assign out_quotient = different_signs ? -comp_out_q : comp_out_q;

  // Remainder is computed as:
  //  t0 = |left| % |right|
  //  t1 = if left * right < 0 and t0 != 0 then |right| - t0 else t0
  //  rem = if right < 0 then -t1 else t1
  assign out_rem_intermediate = different_signs & |comp_out_r ? $signed(right_save - comp_out_r) : comp_out_r;
  assign out_remainder = right_sign ? -out_rem_intermediate : out_rem_intermediate;

  std_div_pipe #(
    .WIDTH(WIDTH)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left_abs),
    .right(right_abs),
    .out_quotient(comp_out_q),
    .out_remainder(comp_out_r)
  );

  // Simulation self test against unsynthesizable implementation.
  `ifdef VERILATOR
    logic signed [WIDTH-1:0] l, r;
    always_ff @(posedge clk) begin
      if (go) begin
        l <= left;
        r <= right;
      end else begin
        l <= l;
        r <= r;
      end
    end

    always @(posedge clk) begin
      if (done && out_quotient != $signed(l / r))
        $error(
          "\nstd_sdiv_pipe (Quotient): Computed and golden outputs do not match!\n",
          "left: %0d", l,
          "  right: %0d\n", r,
          "expected: %0d", $signed(l / r),
          "  computed: %0d", $signed(out_quotient),
        );
      if (done && out_remainder != $signed(((l % r) + r) % r))
        $error(
          "\nstd_sdiv_pipe (Remainder): Computed and golden outputs do not match!\n",
          "left: %0d", l,
          "  right: %0d\n", r,
          "expected: %0d", $signed(((l % r) + r) % r),
          "  computed: %0d", $signed(out_remainder),
        );
    end
  `endif
endmodule

module std_sgt #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left > right);
endmodule

module std_slt #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left < right);
endmodule

module std_seq #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left == right);
endmodule

module std_sneq #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left != right);
endmodule

module std_sge #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left >= right);
endmodule

module std_sle #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left <= right);
endmodule

module std_slsh #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = left <<< right;
endmodule

module std_srsh #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = left >>> right;
endmodule

/**
 * Core primitives for Calyx.
 * Implements core primitives used by the compiler.
 *
 * Conventions:
 * - All parameter names must be SNAKE_CASE and all caps.
 * - Port names must be snake_case, no caps.
 */
`default_nettype none

module std_slice #(
    parameter IN_WIDTH  = 32,
    parameter OUT_WIDTH = 32
) (
   input wire                   logic [ IN_WIDTH-1:0] in,
   output logic [OUT_WIDTH-1:0] out
);
  assign out = in[OUT_WIDTH-1:0];

  `ifdef VERILATOR
    always_comb begin
      if (IN_WIDTH < OUT_WIDTH)
        $error(
          "std_slice: Input width less than output width\n",
          "IN_WIDTH: %0d", IN_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_pad #(
    parameter IN_WIDTH  = 32,
    parameter OUT_WIDTH = 32
) (
   input wire logic [IN_WIDTH-1:0]  in,
   output logic     [OUT_WIDTH-1:0] out
);
  localparam EXTEND = OUT_WIDTH - IN_WIDTH;
  assign out = { {EXTEND {1'b0}}, in};

  `ifdef VERILATOR
    always_comb begin
      if (IN_WIDTH > OUT_WIDTH)
        $error(
          "std_pad: Output width less than input width\n",
          "IN_WIDTH: %0d", IN_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_cat #(
  parameter LEFT_WIDTH  = 32,
  parameter RIGHT_WIDTH = 32,
  parameter OUT_WIDTH = 64
) (
  input wire logic [LEFT_WIDTH-1:0] left,
  input wire logic [RIGHT_WIDTH-1:0] right,
  output logic [OUT_WIDTH-1:0] out
);
  assign out = {left, right};

  `ifdef VERILATOR
    always_comb begin
      if (LEFT_WIDTH + RIGHT_WIDTH != OUT_WIDTH)
        $error(
          "std_cat: Output width must equal sum of input widths\n",
          "LEFT_WIDTH: %0d", LEFT_WIDTH,
          "RIGHT_WIDTH: %0d", RIGHT_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_not #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] in,
   output logic [WIDTH-1:0] out
);
  assign out = ~in;
endmodule

module std_and #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left & right;
endmodule

module std_or #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left | right;
endmodule

module std_xor #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left ^ right;
endmodule

module std_sub #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module std_gt #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left > right;
endmodule

module std_lt #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left < right;
endmodule

module std_eq #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left == right;
endmodule

module std_neq #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left != right;
endmodule

module std_ge #(
    parameter WIDTH = 32
) (
    input wire   logic [WIDTH-1:0] left,
    input wire   logic [WIDTH-1:0] right,
    output logic out
);
  assign out = left >= right;
endmodule

module std_le #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left <= right;
endmodule

module std_lsh #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left << right;
endmodule

module std_rsh #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left >> right;
endmodule

/// this primitive is intended to be used
/// for lowering purposes (not in source programs)
module std_mux #(
    parameter WIDTH = 32
) (
   input wire               logic cond,
   input wire               logic [WIDTH-1:0] tru,
   input wire               logic [WIDTH-1:0] fal,
   output logic [WIDTH-1:0] out
);
  assign out = cond ? tru : fal;
endmodule

module std_mem_d1 #(
    parameter WIDTH = 32,
    parameter SIZE = 16,
    parameter IDX_SIZE = 4
) (
   input wire                logic [IDX_SIZE-1:0] addr0,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  logic [WIDTH-1:0] mem[SIZE-1:0];

  /* verilator lint_off WIDTH */
  assign read_data = mem[addr0];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= SIZE)
        $error(
          "std_mem_d1: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "SIZE: %0d", SIZE
        );
    end
  `endif
endmodule

module std_mem_d2 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0];

  assign read_data = mem[addr0][addr1];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d2: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d2: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
    end
  `endif
endmodule

module std_mem_d3 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D2_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4,
    parameter D2_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [D2_IDX_SIZE-1:0] addr2,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0][D2_SIZE-1:0];

  assign read_data = mem[addr0][addr1][addr2];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1][addr2] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
      if (addr2 >= D2_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr2: %0d\n", addr2,
          "D2_SIZE: %0d", D2_SIZE
        );
    end
  `endif
endmodule

module std_mem_d4 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D2_SIZE = 16,
    parameter D3_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4,
    parameter D2_IDX_SIZE = 4,
    parameter D3_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [D2_IDX_SIZE-1:0] addr2,
   input wire                logic [D3_IDX_SIZE-1:0] addr3,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0][D2_SIZE-1:0][D3_SIZE-1:0];

  assign read_data = mem[addr0][addr1][addr2][addr3];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1][addr2][addr3] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
      if (addr2 >= D2_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr2: %0d\n", addr2,
          "D2_SIZE: %0d", D2_SIZE
        );
      if (addr3 >= D3_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr3: %0d\n", addr3,
          "D3_SIZE: %0d", D3_SIZE
        );
    end
  `endif
endmodule

`default_nettype wire

module undef #(
    parameter WIDTH = 32
) (
   output logic [WIDTH-1:0] out
);
assign out = 'x;
endmodule

module std_const #(
    parameter WIDTH = 32,
    parameter VALUE = 32
) (
   output logic [WIDTH-1:0] out
);
assign out = VALUE;
endmodule

module std_wire #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] in,
   output logic [WIDTH-1:0] out
);
assign out = in;
endmodule

module std_add #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] left,
   input logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
assign out = left + right;
endmodule

module std_reg #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] in,
   input logic write_en,
   input logic clk,
   input logic reset,
   output logic [WIDTH-1:0] out,
   output logic done
);
always_ff @(posedge clk) begin
    if (reset) begin
       out <= 0;
       done <= 0;
    end else if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module mac_pe(
  input logic [31:0] top,
  input logic [31:0] left,
  input logic mul_ready,
  output logic [31:0] out,
  input logic go,
  input logic clk,
  input logic reset,
  output logic done
);
// COMPONENT START: mac_pe
logic [31:0] acc_in;
logic acc_write_en;
logic acc_clk;
logic acc_reset;
logic [31:0] acc_out;
logic acc_done;
logic [31:0] add_left;
logic [31:0] add_right;
logic [31:0] add_out;
logic mul_clk;
logic [31:0] mul_left;
logic [31:0] mul_right;
logic [31:0] mul_out;
logic fsm_in;
logic fsm_write_en;
logic fsm_clk;
logic fsm_reset;
logic fsm_out;
logic fsm_done;
logic ud_out;
logic adder_left;
logic adder_right;
logic adder_out;
logic signal_reg_in;
logic signal_reg_write_en;
logic signal_reg_clk;
logic signal_reg_reset;
logic signal_reg_out;
logic signal_reg_done;
logic early_reset_static_par_go_in;
logic early_reset_static_par_go_out;
logic early_reset_static_par_done_in;
logic early_reset_static_par_done_out;
logic wrapper_early_reset_static_par_go_in;
logic wrapper_early_reset_static_par_go_out;
logic wrapper_early_reset_static_par_done_in;
logic wrapper_early_reset_static_par_done_out;
std_reg # (
    .WIDTH(32)
) acc (
    .clk(acc_clk),
    .done(acc_done),
    .in(acc_in),
    .out(acc_out),
    .reset(acc_reset),
    .write_en(acc_write_en)
);
std_add # (
    .WIDTH(32)
) add (
    .left(add_left),
    .out(add_out),
    .right(add_right)
);
bb_pipelined_mult mul (
    .clk(mul_clk),
    .left(mul_left),
    .out(mul_out),
    .right(mul_right)
);
std_reg # (
    .WIDTH(1)
) fsm (
    .clk(fsm_clk),
    .done(fsm_done),
    .in(fsm_in),
    .out(fsm_out),
    .reset(fsm_reset),
    .write_en(fsm_write_en)
);
undef # (
    .WIDTH(1)
) ud (
    .out(ud_out)
);
std_add # (
    .WIDTH(1)
) adder (
    .left(adder_left),
    .out(adder_out),
    .right(adder_right)
);
std_reg # (
    .WIDTH(1)
) signal_reg (
    .clk(signal_reg_clk),
    .done(signal_reg_done),
    .in(signal_reg_in),
    .out(signal_reg_out),
    .reset(signal_reg_reset),
    .write_en(signal_reg_write_en)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_go (
    .in(early_reset_static_par_go_in),
    .out(early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_done (
    .in(early_reset_static_par_done_in),
    .out(early_reset_static_par_done_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_go (
    .in(wrapper_early_reset_static_par_go_in),
    .out(wrapper_early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_done (
    .in(wrapper_early_reset_static_par_done_in),
    .out(wrapper_early_reset_static_par_done_out)
);
wire _guard0 = 1;
wire _guard1 = early_reset_static_par_go_out;
wire _guard2 = early_reset_static_par_go_out;
wire _guard3 = wrapper_early_reset_static_par_done_out;
wire _guard4 = early_reset_static_par_go_out;
wire _guard5 = fsm_out != 1'd0;
wire _guard6 = early_reset_static_par_go_out;
wire _guard7 = _guard5 & _guard6;
wire _guard8 = fsm_out == 1'd0;
wire _guard9 = early_reset_static_par_go_out;
wire _guard10 = _guard8 & _guard9;
wire _guard11 = early_reset_static_par_go_out;
wire _guard12 = early_reset_static_par_go_out;
wire _guard13 = fsm_out == 1'd0;
wire _guard14 = signal_reg_out;
wire _guard15 = _guard13 & _guard14;
wire _guard16 = fsm_out == 1'd0;
wire _guard17 = signal_reg_out;
wire _guard18 = _guard16 & _guard17;
wire _guard19 = fsm_out == 1'd0;
wire _guard20 = signal_reg_out;
wire _guard21 = ~_guard20;
wire _guard22 = _guard19 & _guard21;
wire _guard23 = wrapper_early_reset_static_par_go_out;
wire _guard24 = _guard22 & _guard23;
wire _guard25 = _guard18 | _guard24;
wire _guard26 = fsm_out == 1'd0;
wire _guard27 = signal_reg_out;
wire _guard28 = ~_guard27;
wire _guard29 = _guard26 & _guard28;
wire _guard30 = wrapper_early_reset_static_par_go_out;
wire _guard31 = _guard29 & _guard30;
wire _guard32 = fsm_out == 1'd0;
wire _guard33 = signal_reg_out;
wire _guard34 = _guard32 & _guard33;
wire _guard35 = early_reset_static_par_go_out;
wire _guard36 = early_reset_static_par_go_out;
wire _guard37 = early_reset_static_par_go_out;
wire _guard38 = early_reset_static_par_go_out;
wire _guard39 = wrapper_early_reset_static_par_go_out;
assign acc_write_en =
  _guard1 ? mul_ready :
  1'd0;
assign acc_clk = clk;
assign acc_reset = reset;
assign acc_in = add_out;
assign done = _guard3;
assign out = acc_out;
assign fsm_write_en = _guard4;
assign fsm_clk = clk;
assign fsm_reset = reset;
assign fsm_in =
  _guard7 ? adder_out :
  _guard10 ? 1'd0 :
  1'd0;
assign adder_left =
  _guard11 ? fsm_out :
  1'd0;
assign adder_right = _guard12;
assign wrapper_early_reset_static_par_go_in = go;
assign wrapper_early_reset_static_par_done_in = _guard15;
assign early_reset_static_par_done_in = ud_out;
assign signal_reg_write_en = _guard25;
assign signal_reg_clk = clk;
assign signal_reg_reset = reset;
assign signal_reg_in =
  _guard31 ? 1'd1 :
  _guard34 ? 1'd0 :
  1'd0;
assign add_left = acc_out;
assign add_right = mul_out;
assign mul_clk = clk;
assign mul_left =
  _guard37 ? top :
  32'd0;
assign mul_right =
  _guard38 ? left :
  32'd0;
assign early_reset_static_par_go_in = _guard39;
// COMPONENT END: mac_pe
endmodule
module systolic_array_comp(
  input logic [31:0] depth,
  input logic [31:0] t0_read_data,
  input logic [31:0] t1_read_data,
  input logic [31:0] l0_read_data,
  input logic [31:0] l1_read_data,
  output logic [1:0] t0_addr0,
  output logic [1:0] t1_addr0,
  output logic [1:0] l0_addr0,
  output logic [1:0] l1_addr0,
  output logic [31:0] out_mem_0_addr0,
  output logic [31:0] out_mem_0_write_data,
  output logic out_mem_0_write_en,
  output logic [31:0] out_mem_1_addr0,
  output logic [31:0] out_mem_1_write_data,
  output logic out_mem_1_write_en,
  input logic go,
  input logic clk,
  input logic reset,
  output logic done
);
// COMPONENT START: systolic_array_comp
logic [31:0] min_depth_4_in;
logic min_depth_4_write_en;
logic min_depth_4_clk;
logic min_depth_4_reset;
logic [31:0] min_depth_4_out;
logic min_depth_4_done;
logic [31:0] iter_limit_in;
logic iter_limit_write_en;
logic iter_limit_clk;
logic iter_limit_reset;
logic [31:0] iter_limit_out;
logic iter_limit_done;
logic [31:0] depth_plus_5_left;
logic [31:0] depth_plus_5_right;
logic [31:0] depth_plus_5_out;
logic [31:0] depth_plus_2_left;
logic [31:0] depth_plus_2_right;
logic [31:0] depth_plus_2_out;
logic [31:0] depth_plus_7_left;
logic [31:0] depth_plus_7_right;
logic [31:0] depth_plus_7_out;
logic [31:0] depth_plus_0_left;
logic [31:0] depth_plus_0_right;
logic [31:0] depth_plus_0_out;
logic [31:0] min_depth_4_plus_1_left;
logic [31:0] min_depth_4_plus_1_right;
logic [31:0] min_depth_4_plus_1_out;
logic [31:0] depth_plus_1_left;
logic [31:0] depth_plus_1_right;
logic [31:0] depth_plus_1_out;
logic [31:0] depth_plus_6_left;
logic [31:0] depth_plus_6_right;
logic [31:0] depth_plus_6_out;
logic [31:0] min_depth_4_plus_3_left;
logic [31:0] min_depth_4_plus_3_right;
logic [31:0] min_depth_4_plus_3_out;
logic [31:0] min_depth_4_plus_2_left;
logic [31:0] min_depth_4_plus_2_right;
logic [31:0] min_depth_4_plus_2_out;
logic [31:0] depth_plus_8_left;
logic [31:0] depth_plus_8_right;
logic [31:0] depth_plus_8_out;
logic [31:0] pe_0_0_top;
logic [31:0] pe_0_0_left;
logic pe_0_0_mul_ready;
logic [31:0] pe_0_0_out;
logic pe_0_0_go;
logic pe_0_0_clk;
logic pe_0_0_reset;
logic pe_0_0_done;
logic [31:0] top_0_0_in;
logic top_0_0_write_en;
logic top_0_0_clk;
logic top_0_0_reset;
logic [31:0] top_0_0_out;
logic top_0_0_done;
logic [31:0] left_0_0_in;
logic left_0_0_write_en;
logic left_0_0_clk;
logic left_0_0_reset;
logic [31:0] left_0_0_out;
logic left_0_0_done;
logic [31:0] pe_0_1_top;
logic [31:0] pe_0_1_left;
logic pe_0_1_mul_ready;
logic [31:0] pe_0_1_out;
logic pe_0_1_go;
logic pe_0_1_clk;
logic pe_0_1_reset;
logic pe_0_1_done;
logic [31:0] top_0_1_in;
logic top_0_1_write_en;
logic top_0_1_clk;
logic top_0_1_reset;
logic [31:0] top_0_1_out;
logic top_0_1_done;
logic [31:0] left_0_1_in;
logic left_0_1_write_en;
logic left_0_1_clk;
logic left_0_1_reset;
logic [31:0] left_0_1_out;
logic left_0_1_done;
logic [31:0] pe_1_0_top;
logic [31:0] pe_1_0_left;
logic pe_1_0_mul_ready;
logic [31:0] pe_1_0_out;
logic pe_1_0_go;
logic pe_1_0_clk;
logic pe_1_0_reset;
logic pe_1_0_done;
logic [31:0] top_1_0_in;
logic top_1_0_write_en;
logic top_1_0_clk;
logic top_1_0_reset;
logic [31:0] top_1_0_out;
logic top_1_0_done;
logic [31:0] left_1_0_in;
logic left_1_0_write_en;
logic left_1_0_clk;
logic left_1_0_reset;
logic [31:0] left_1_0_out;
logic left_1_0_done;
logic [31:0] pe_1_1_top;
logic [31:0] pe_1_1_left;
logic pe_1_1_mul_ready;
logic [31:0] pe_1_1_out;
logic pe_1_1_go;
logic pe_1_1_clk;
logic pe_1_1_reset;
logic pe_1_1_done;
logic [31:0] top_1_1_in;
logic top_1_1_write_en;
logic top_1_1_clk;
logic top_1_1_reset;
logic [31:0] top_1_1_out;
logic top_1_1_done;
logic [31:0] left_1_1_in;
logic left_1_1_write_en;
logic left_1_1_clk;
logic left_1_1_reset;
logic [31:0] left_1_1_out;
logic left_1_1_done;
logic [1:0] t0_idx_in;
logic t0_idx_write_en;
logic t0_idx_clk;
logic t0_idx_reset;
logic [1:0] t0_idx_out;
logic t0_idx_done;
logic [1:0] t0_add_left;
logic [1:0] t0_add_right;
logic [1:0] t0_add_out;
logic [1:0] t1_idx_in;
logic t1_idx_write_en;
logic t1_idx_clk;
logic t1_idx_reset;
logic [1:0] t1_idx_out;
logic t1_idx_done;
logic [1:0] t1_add_left;
logic [1:0] t1_add_right;
logic [1:0] t1_add_out;
logic [1:0] l0_idx_in;
logic l0_idx_write_en;
logic l0_idx_clk;
logic l0_idx_reset;
logic [1:0] l0_idx_out;
logic l0_idx_done;
logic [1:0] l0_add_left;
logic [1:0] l0_add_right;
logic [1:0] l0_add_out;
logic [1:0] l1_idx_in;
logic l1_idx_write_en;
logic l1_idx_clk;
logic l1_idx_reset;
logic [1:0] l1_idx_out;
logic l1_idx_done;
logic [1:0] l1_add_left;
logic [1:0] l1_add_right;
logic [1:0] l1_add_out;
logic [31:0] idx_in;
logic idx_write_en;
logic idx_clk;
logic idx_reset;
logic [31:0] idx_out;
logic idx_done;
logic [31:0] idx_add_left;
logic [31:0] idx_add_right;
logic [31:0] idx_add_out;
logic [31:0] lt_iter_limit_left;
logic [31:0] lt_iter_limit_right;
logic lt_iter_limit_out;
logic cond_reg_in;
logic cond_reg_write_en;
logic cond_reg_clk;
logic cond_reg_reset;
logic cond_reg_out;
logic cond_reg_done;
logic idx_between_5_depth_plus_5_reg_in;
logic idx_between_5_depth_plus_5_reg_write_en;
logic idx_between_5_depth_plus_5_reg_clk;
logic idx_between_5_depth_plus_5_reg_reset;
logic idx_between_5_depth_plus_5_reg_out;
logic idx_between_5_depth_plus_5_reg_done;
logic [31:0] index_lt_depth_plus_5_left;
logic [31:0] index_lt_depth_plus_5_right;
logic index_lt_depth_plus_5_out;
logic [31:0] index_ge_5_left;
logic [31:0] index_ge_5_right;
logic index_ge_5_out;
logic idx_between_5_depth_plus_5_comb_left;
logic idx_between_5_depth_plus_5_comb_right;
logic idx_between_5_depth_plus_5_comb_out;
logic idx_between_2_depth_plus_2_reg_in;
logic idx_between_2_depth_plus_2_reg_write_en;
logic idx_between_2_depth_plus_2_reg_clk;
logic idx_between_2_depth_plus_2_reg_reset;
logic idx_between_2_depth_plus_2_reg_out;
logic idx_between_2_depth_plus_2_reg_done;
logic [31:0] index_lt_depth_plus_2_left;
logic [31:0] index_lt_depth_plus_2_right;
logic index_lt_depth_plus_2_out;
logic [31:0] index_ge_2_left;
logic [31:0] index_ge_2_right;
logic index_ge_2_out;
logic idx_between_2_depth_plus_2_comb_left;
logic idx_between_2_depth_plus_2_comb_right;
logic idx_between_2_depth_plus_2_comb_out;
logic idx_between_7_depth_plus_7_reg_in;
logic idx_between_7_depth_plus_7_reg_write_en;
logic idx_between_7_depth_plus_7_reg_clk;
logic idx_between_7_depth_plus_7_reg_reset;
logic idx_between_7_depth_plus_7_reg_out;
logic idx_between_7_depth_plus_7_reg_done;
logic [31:0] index_lt_depth_plus_7_left;
logic [31:0] index_lt_depth_plus_7_right;
logic index_lt_depth_plus_7_out;
logic [31:0] index_ge_7_left;
logic [31:0] index_ge_7_right;
logic index_ge_7_out;
logic idx_between_7_depth_plus_7_comb_left;
logic idx_between_7_depth_plus_7_comb_right;
logic idx_between_7_depth_plus_7_comb_out;
logic idx_between_0_depth_plus_0_reg_in;
logic idx_between_0_depth_plus_0_reg_write_en;
logic idx_between_0_depth_plus_0_reg_clk;
logic idx_between_0_depth_plus_0_reg_reset;
logic idx_between_0_depth_plus_0_reg_out;
logic idx_between_0_depth_plus_0_reg_done;
logic [31:0] index_lt_depth_plus_0_left;
logic [31:0] index_lt_depth_plus_0_right;
logic index_lt_depth_plus_0_out;
logic idx_between_1_min_depth_4_plus_1_reg_in;
logic idx_between_1_min_depth_4_plus_1_reg_write_en;
logic idx_between_1_min_depth_4_plus_1_reg_clk;
logic idx_between_1_min_depth_4_plus_1_reg_reset;
logic idx_between_1_min_depth_4_plus_1_reg_out;
logic idx_between_1_min_depth_4_plus_1_reg_done;
logic [31:0] index_lt_min_depth_4_plus_1_left;
logic [31:0] index_lt_min_depth_4_plus_1_right;
logic index_lt_min_depth_4_plus_1_out;
logic [31:0] index_ge_1_left;
logic [31:0] index_ge_1_right;
logic index_ge_1_out;
logic idx_between_1_min_depth_4_plus_1_comb_left;
logic idx_between_1_min_depth_4_plus_1_comb_right;
logic idx_between_1_min_depth_4_plus_1_comb_out;
logic idx_between_1_depth_plus_1_reg_in;
logic idx_between_1_depth_plus_1_reg_write_en;
logic idx_between_1_depth_plus_1_reg_clk;
logic idx_between_1_depth_plus_1_reg_reset;
logic idx_between_1_depth_plus_1_reg_out;
logic idx_between_1_depth_plus_1_reg_done;
logic [31:0] index_lt_depth_plus_1_left;
logic [31:0] index_lt_depth_plus_1_right;
logic index_lt_depth_plus_1_out;
logic idx_between_1_depth_plus_1_comb_left;
logic idx_between_1_depth_plus_1_comb_right;
logic idx_between_1_depth_plus_1_comb_out;
logic idx_between_depth_plus_6_depth_plus_7_reg_in;
logic idx_between_depth_plus_6_depth_plus_7_reg_write_en;
logic idx_between_depth_plus_6_depth_plus_7_reg_clk;
logic idx_between_depth_plus_6_depth_plus_7_reg_reset;
logic idx_between_depth_plus_6_depth_plus_7_reg_out;
logic idx_between_depth_plus_6_depth_plus_7_reg_done;
logic [31:0] index_ge_depth_plus_6_left;
logic [31:0] index_ge_depth_plus_6_right;
logic index_ge_depth_plus_6_out;
logic idx_between_depth_plus_6_depth_plus_7_comb_left;
logic idx_between_depth_plus_6_depth_plus_7_comb_right;
logic idx_between_depth_plus_6_depth_plus_7_comb_out;
logic idx_between_3_min_depth_4_plus_3_reg_in;
logic idx_between_3_min_depth_4_plus_3_reg_write_en;
logic idx_between_3_min_depth_4_plus_3_reg_clk;
logic idx_between_3_min_depth_4_plus_3_reg_reset;
logic idx_between_3_min_depth_4_plus_3_reg_out;
logic idx_between_3_min_depth_4_plus_3_reg_done;
logic [31:0] index_lt_min_depth_4_plus_3_left;
logic [31:0] index_lt_min_depth_4_plus_3_right;
logic index_lt_min_depth_4_plus_3_out;
logic [31:0] index_ge_3_left;
logic [31:0] index_ge_3_right;
logic index_ge_3_out;
logic idx_between_3_min_depth_4_plus_3_comb_left;
logic idx_between_3_min_depth_4_plus_3_comb_right;
logic idx_between_3_min_depth_4_plus_3_comb_out;
logic idx_between_depth_plus_5_depth_plus_6_reg_in;
logic idx_between_depth_plus_5_depth_plus_6_reg_write_en;
logic idx_between_depth_plus_5_depth_plus_6_reg_clk;
logic idx_between_depth_plus_5_depth_plus_6_reg_reset;
logic idx_between_depth_plus_5_depth_plus_6_reg_out;
logic idx_between_depth_plus_5_depth_plus_6_reg_done;
logic [31:0] index_lt_depth_plus_6_left;
logic [31:0] index_lt_depth_plus_6_right;
logic index_lt_depth_plus_6_out;
logic [31:0] index_ge_depth_plus_5_left;
logic [31:0] index_ge_depth_plus_5_right;
logic index_ge_depth_plus_5_out;
logic idx_between_depth_plus_5_depth_plus_6_comb_left;
logic idx_between_depth_plus_5_depth_plus_6_comb_right;
logic idx_between_depth_plus_5_depth_plus_6_comb_out;
logic idx_between_2_min_depth_4_plus_2_reg_in;
logic idx_between_2_min_depth_4_plus_2_reg_write_en;
logic idx_between_2_min_depth_4_plus_2_reg_clk;
logic idx_between_2_min_depth_4_plus_2_reg_reset;
logic idx_between_2_min_depth_4_plus_2_reg_out;
logic idx_between_2_min_depth_4_plus_2_reg_done;
logic [31:0] index_lt_min_depth_4_plus_2_left;
logic [31:0] index_lt_min_depth_4_plus_2_right;
logic index_lt_min_depth_4_plus_2_out;
logic idx_between_2_min_depth_4_plus_2_comb_left;
logic idx_between_2_min_depth_4_plus_2_comb_right;
logic idx_between_2_min_depth_4_plus_2_comb_out;
logic idx_between_6_depth_plus_6_reg_in;
logic idx_between_6_depth_plus_6_reg_write_en;
logic idx_between_6_depth_plus_6_reg_clk;
logic idx_between_6_depth_plus_6_reg_reset;
logic idx_between_6_depth_plus_6_reg_out;
logic idx_between_6_depth_plus_6_reg_done;
logic [31:0] index_ge_6_left;
logic [31:0] index_ge_6_right;
logic index_ge_6_out;
logic idx_between_6_depth_plus_6_comb_left;
logic idx_between_6_depth_plus_6_comb_right;
logic idx_between_6_depth_plus_6_comb_out;
logic idx_between_depth_plus_7_depth_plus_8_reg_in;
logic idx_between_depth_plus_7_depth_plus_8_reg_write_en;
logic idx_between_depth_plus_7_depth_plus_8_reg_clk;
logic idx_between_depth_plus_7_depth_plus_8_reg_reset;
logic idx_between_depth_plus_7_depth_plus_8_reg_out;
logic idx_between_depth_plus_7_depth_plus_8_reg_done;
logic [31:0] index_lt_depth_plus_8_left;
logic [31:0] index_lt_depth_plus_8_right;
logic index_lt_depth_plus_8_out;
logic [31:0] index_ge_depth_plus_7_left;
logic [31:0] index_ge_depth_plus_7_right;
logic index_ge_depth_plus_7_out;
logic idx_between_depth_plus_7_depth_plus_8_comb_left;
logic idx_between_depth_plus_7_depth_plus_8_comb_right;
logic idx_between_depth_plus_7_depth_plus_8_comb_out;
logic cond_in;
logic cond_write_en;
logic cond_clk;
logic cond_reset;
logic cond_out;
logic cond_done;
logic cond_wire_in;
logic cond_wire_out;
logic cond0_in;
logic cond0_write_en;
logic cond0_clk;
logic cond0_reset;
logic cond0_out;
logic cond0_done;
logic cond_wire0_in;
logic cond_wire0_out;
logic cond1_in;
logic cond1_write_en;
logic cond1_clk;
logic cond1_reset;
logic cond1_out;
logic cond1_done;
logic cond_wire1_in;
logic cond_wire1_out;
logic cond2_in;
logic cond2_write_en;
logic cond2_clk;
logic cond2_reset;
logic cond2_out;
logic cond2_done;
logic cond_wire2_in;
logic cond_wire2_out;
logic cond3_in;
logic cond3_write_en;
logic cond3_clk;
logic cond3_reset;
logic cond3_out;
logic cond3_done;
logic cond_wire3_in;
logic cond_wire3_out;
logic cond4_in;
logic cond4_write_en;
logic cond4_clk;
logic cond4_reset;
logic cond4_out;
logic cond4_done;
logic cond_wire4_in;
logic cond_wire4_out;
logic cond5_in;
logic cond5_write_en;
logic cond5_clk;
logic cond5_reset;
logic cond5_out;
logic cond5_done;
logic cond_wire5_in;
logic cond_wire5_out;
logic cond6_in;
logic cond6_write_en;
logic cond6_clk;
logic cond6_reset;
logic cond6_out;
logic cond6_done;
logic cond_wire6_in;
logic cond_wire6_out;
logic cond7_in;
logic cond7_write_en;
logic cond7_clk;
logic cond7_reset;
logic cond7_out;
logic cond7_done;
logic cond_wire7_in;
logic cond_wire7_out;
logic cond8_in;
logic cond8_write_en;
logic cond8_clk;
logic cond8_reset;
logic cond8_out;
logic cond8_done;
logic cond_wire8_in;
logic cond_wire8_out;
logic cond9_in;
logic cond9_write_en;
logic cond9_clk;
logic cond9_reset;
logic cond9_out;
logic cond9_done;
logic cond_wire9_in;
logic cond_wire9_out;
logic cond10_in;
logic cond10_write_en;
logic cond10_clk;
logic cond10_reset;
logic cond10_out;
logic cond10_done;
logic cond_wire10_in;
logic cond_wire10_out;
logic cond11_in;
logic cond11_write_en;
logic cond11_clk;
logic cond11_reset;
logic cond11_out;
logic cond11_done;
logic cond_wire11_in;
logic cond_wire11_out;
logic cond12_in;
logic cond12_write_en;
logic cond12_clk;
logic cond12_reset;
logic cond12_out;
logic cond12_done;
logic cond_wire12_in;
logic cond_wire12_out;
logic cond13_in;
logic cond13_write_en;
logic cond13_clk;
logic cond13_reset;
logic cond13_out;
logic cond13_done;
logic cond_wire13_in;
logic cond_wire13_out;
logic cond14_in;
logic cond14_write_en;
logic cond14_clk;
logic cond14_reset;
logic cond14_out;
logic cond14_done;
logic cond_wire14_in;
logic cond_wire14_out;
logic cond15_in;
logic cond15_write_en;
logic cond15_clk;
logic cond15_reset;
logic cond15_out;
logic cond15_done;
logic cond_wire15_in;
logic cond_wire15_out;
logic cond16_in;
logic cond16_write_en;
logic cond16_clk;
logic cond16_reset;
logic cond16_out;
logic cond16_done;
logic cond_wire16_in;
logic cond_wire16_out;
logic fsm_in;
logic fsm_write_en;
logic fsm_clk;
logic fsm_reset;
logic fsm_out;
logic fsm_done;
logic ud_out;
logic adder_left;
logic adder_right;
logic adder_out;
logic ud0_out;
logic adder0_left;
logic adder0_right;
logic adder0_out;
logic signal_reg_in;
logic signal_reg_write_en;
logic signal_reg_clk;
logic signal_reg_reset;
logic signal_reg_out;
logic signal_reg_done;
logic [1:0] fsm0_in;
logic fsm0_write_en;
logic fsm0_clk;
logic fsm0_reset;
logic [1:0] fsm0_out;
logic fsm0_done;
logic early_reset_static_par_go_in;
logic early_reset_static_par_go_out;
logic early_reset_static_par_done_in;
logic early_reset_static_par_done_out;
logic early_reset_static_par0_go_in;
logic early_reset_static_par0_go_out;
logic early_reset_static_par0_done_in;
logic early_reset_static_par0_done_out;
logic wrapper_early_reset_static_par_go_in;
logic wrapper_early_reset_static_par_go_out;
logic wrapper_early_reset_static_par_done_in;
logic wrapper_early_reset_static_par_done_out;
logic while_wrapper_early_reset_static_par0_go_in;
logic while_wrapper_early_reset_static_par0_go_out;
logic while_wrapper_early_reset_static_par0_done_in;
logic while_wrapper_early_reset_static_par0_done_out;
logic tdcc_go_in;
logic tdcc_go_out;
logic tdcc_done_in;
logic tdcc_done_out;
std_reg # (
    .WIDTH(32)
) min_depth_4 (
    .clk(min_depth_4_clk),
    .done(min_depth_4_done),
    .in(min_depth_4_in),
    .out(min_depth_4_out),
    .reset(min_depth_4_reset),
    .write_en(min_depth_4_write_en)
);
std_reg # (
    .WIDTH(32)
) iter_limit (
    .clk(iter_limit_clk),
    .done(iter_limit_done),
    .in(iter_limit_in),
    .out(iter_limit_out),
    .reset(iter_limit_reset),
    .write_en(iter_limit_write_en)
);
std_add # (
    .WIDTH(32)
) depth_plus_5 (
    .left(depth_plus_5_left),
    .out(depth_plus_5_out),
    .right(depth_plus_5_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_2 (
    .left(depth_plus_2_left),
    .out(depth_plus_2_out),
    .right(depth_plus_2_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_7 (
    .left(depth_plus_7_left),
    .out(depth_plus_7_out),
    .right(depth_plus_7_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_0 (
    .left(depth_plus_0_left),
    .out(depth_plus_0_out),
    .right(depth_plus_0_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_1 (
    .left(min_depth_4_plus_1_left),
    .out(min_depth_4_plus_1_out),
    .right(min_depth_4_plus_1_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_1 (
    .left(depth_plus_1_left),
    .out(depth_plus_1_out),
    .right(depth_plus_1_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_6 (
    .left(depth_plus_6_left),
    .out(depth_plus_6_out),
    .right(depth_plus_6_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_3 (
    .left(min_depth_4_plus_3_left),
    .out(min_depth_4_plus_3_out),
    .right(min_depth_4_plus_3_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_2 (
    .left(min_depth_4_plus_2_left),
    .out(min_depth_4_plus_2_out),
    .right(min_depth_4_plus_2_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_8 (
    .left(depth_plus_8_left),
    .out(depth_plus_8_out),
    .right(depth_plus_8_right)
);
mac_pe pe_0_0 (
    .clk(pe_0_0_clk),
    .done(pe_0_0_done),
    .go(pe_0_0_go),
    .left(pe_0_0_left),
    .mul_ready(pe_0_0_mul_ready),
    .out(pe_0_0_out),
    .reset(pe_0_0_reset),
    .top(pe_0_0_top)
);
std_reg # (
    .WIDTH(32)
) top_0_0 (
    .clk(top_0_0_clk),
    .done(top_0_0_done),
    .in(top_0_0_in),
    .out(top_0_0_out),
    .reset(top_0_0_reset),
    .write_en(top_0_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_0 (
    .clk(left_0_0_clk),
    .done(left_0_0_done),
    .in(left_0_0_in),
    .out(left_0_0_out),
    .reset(left_0_0_reset),
    .write_en(left_0_0_write_en)
);
mac_pe pe_0_1 (
    .clk(pe_0_1_clk),
    .done(pe_0_1_done),
    .go(pe_0_1_go),
    .left(pe_0_1_left),
    .mul_ready(pe_0_1_mul_ready),
    .out(pe_0_1_out),
    .reset(pe_0_1_reset),
    .top(pe_0_1_top)
);
std_reg # (
    .WIDTH(32)
) top_0_1 (
    .clk(top_0_1_clk),
    .done(top_0_1_done),
    .in(top_0_1_in),
    .out(top_0_1_out),
    .reset(top_0_1_reset),
    .write_en(top_0_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_1 (
    .clk(left_0_1_clk),
    .done(left_0_1_done),
    .in(left_0_1_in),
    .out(left_0_1_out),
    .reset(left_0_1_reset),
    .write_en(left_0_1_write_en)
);
mac_pe pe_1_0 (
    .clk(pe_1_0_clk),
    .done(pe_1_0_done),
    .go(pe_1_0_go),
    .left(pe_1_0_left),
    .mul_ready(pe_1_0_mul_ready),
    .out(pe_1_0_out),
    .reset(pe_1_0_reset),
    .top(pe_1_0_top)
);
std_reg # (
    .WIDTH(32)
) top_1_0 (
    .clk(top_1_0_clk),
    .done(top_1_0_done),
    .in(top_1_0_in),
    .out(top_1_0_out),
    .reset(top_1_0_reset),
    .write_en(top_1_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_0 (
    .clk(left_1_0_clk),
    .done(left_1_0_done),
    .in(left_1_0_in),
    .out(left_1_0_out),
    .reset(left_1_0_reset),
    .write_en(left_1_0_write_en)
);
mac_pe pe_1_1 (
    .clk(pe_1_1_clk),
    .done(pe_1_1_done),
    .go(pe_1_1_go),
    .left(pe_1_1_left),
    .mul_ready(pe_1_1_mul_ready),
    .out(pe_1_1_out),
    .reset(pe_1_1_reset),
    .top(pe_1_1_top)
);
std_reg # (
    .WIDTH(32)
) top_1_1 (
    .clk(top_1_1_clk),
    .done(top_1_1_done),
    .in(top_1_1_in),
    .out(top_1_1_out),
    .reset(top_1_1_reset),
    .write_en(top_1_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_1 (
    .clk(left_1_1_clk),
    .done(left_1_1_done),
    .in(left_1_1_in),
    .out(left_1_1_out),
    .reset(left_1_1_reset),
    .write_en(left_1_1_write_en)
);
std_reg # (
    .WIDTH(2)
) t0_idx (
    .clk(t0_idx_clk),
    .done(t0_idx_done),
    .in(t0_idx_in),
    .out(t0_idx_out),
    .reset(t0_idx_reset),
    .write_en(t0_idx_write_en)
);
std_add # (
    .WIDTH(2)
) t0_add (
    .left(t0_add_left),
    .out(t0_add_out),
    .right(t0_add_right)
);
std_reg # (
    .WIDTH(2)
) t1_idx (
    .clk(t1_idx_clk),
    .done(t1_idx_done),
    .in(t1_idx_in),
    .out(t1_idx_out),
    .reset(t1_idx_reset),
    .write_en(t1_idx_write_en)
);
std_add # (
    .WIDTH(2)
) t1_add (
    .left(t1_add_left),
    .out(t1_add_out),
    .right(t1_add_right)
);
std_reg # (
    .WIDTH(2)
) l0_idx (
    .clk(l0_idx_clk),
    .done(l0_idx_done),
    .in(l0_idx_in),
    .out(l0_idx_out),
    .reset(l0_idx_reset),
    .write_en(l0_idx_write_en)
);
std_add # (
    .WIDTH(2)
) l0_add (
    .left(l0_add_left),
    .out(l0_add_out),
    .right(l0_add_right)
);
std_reg # (
    .WIDTH(2)
) l1_idx (
    .clk(l1_idx_clk),
    .done(l1_idx_done),
    .in(l1_idx_in),
    .out(l1_idx_out),
    .reset(l1_idx_reset),
    .write_en(l1_idx_write_en)
);
std_add # (
    .WIDTH(2)
) l1_add (
    .left(l1_add_left),
    .out(l1_add_out),
    .right(l1_add_right)
);
std_reg # (
    .WIDTH(32)
) idx (
    .clk(idx_clk),
    .done(idx_done),
    .in(idx_in),
    .out(idx_out),
    .reset(idx_reset),
    .write_en(idx_write_en)
);
std_add # (
    .WIDTH(32)
) idx_add (
    .left(idx_add_left),
    .out(idx_add_out),
    .right(idx_add_right)
);
std_lt # (
    .WIDTH(32)
) lt_iter_limit (
    .left(lt_iter_limit_left),
    .out(lt_iter_limit_out),
    .right(lt_iter_limit_right)
);
std_reg # (
    .WIDTH(1)
) cond_reg (
    .clk(cond_reg_clk),
    .done(cond_reg_done),
    .in(cond_reg_in),
    .out(cond_reg_out),
    .reset(cond_reg_reset),
    .write_en(cond_reg_write_en)
);
std_reg # (
    .WIDTH(1)
) idx_between_5_depth_plus_5_reg (
    .clk(idx_between_5_depth_plus_5_reg_clk),
    .done(idx_between_5_depth_plus_5_reg_done),
    .in(idx_between_5_depth_plus_5_reg_in),
    .out(idx_between_5_depth_plus_5_reg_out),
    .reset(idx_between_5_depth_plus_5_reg_reset),
    .write_en(idx_between_5_depth_plus_5_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_5 (
    .left(index_lt_depth_plus_5_left),
    .out(index_lt_depth_plus_5_out),
    .right(index_lt_depth_plus_5_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_5 (
    .left(index_ge_5_left),
    .out(index_ge_5_out),
    .right(index_ge_5_right)
);
std_and # (
    .WIDTH(1)
) idx_between_5_depth_plus_5_comb (
    .left(idx_between_5_depth_plus_5_comb_left),
    .out(idx_between_5_depth_plus_5_comb_out),
    .right(idx_between_5_depth_plus_5_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_2_depth_plus_2_reg (
    .clk(idx_between_2_depth_plus_2_reg_clk),
    .done(idx_between_2_depth_plus_2_reg_done),
    .in(idx_between_2_depth_plus_2_reg_in),
    .out(idx_between_2_depth_plus_2_reg_out),
    .reset(idx_between_2_depth_plus_2_reg_reset),
    .write_en(idx_between_2_depth_plus_2_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_2 (
    .left(index_lt_depth_plus_2_left),
    .out(index_lt_depth_plus_2_out),
    .right(index_lt_depth_plus_2_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_2 (
    .left(index_ge_2_left),
    .out(index_ge_2_out),
    .right(index_ge_2_right)
);
std_and # (
    .WIDTH(1)
) idx_between_2_depth_plus_2_comb (
    .left(idx_between_2_depth_plus_2_comb_left),
    .out(idx_between_2_depth_plus_2_comb_out),
    .right(idx_between_2_depth_plus_2_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_7_depth_plus_7_reg (
    .clk(idx_between_7_depth_plus_7_reg_clk),
    .done(idx_between_7_depth_plus_7_reg_done),
    .in(idx_between_7_depth_plus_7_reg_in),
    .out(idx_between_7_depth_plus_7_reg_out),
    .reset(idx_between_7_depth_plus_7_reg_reset),
    .write_en(idx_between_7_depth_plus_7_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_7 (
    .left(index_lt_depth_plus_7_left),
    .out(index_lt_depth_plus_7_out),
    .right(index_lt_depth_plus_7_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_7 (
    .left(index_ge_7_left),
    .out(index_ge_7_out),
    .right(index_ge_7_right)
);
std_and # (
    .WIDTH(1)
) idx_between_7_depth_plus_7_comb (
    .left(idx_between_7_depth_plus_7_comb_left),
    .out(idx_between_7_depth_plus_7_comb_out),
    .right(idx_between_7_depth_plus_7_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_0_depth_plus_0_reg (
    .clk(idx_between_0_depth_plus_0_reg_clk),
    .done(idx_between_0_depth_plus_0_reg_done),
    .in(idx_between_0_depth_plus_0_reg_in),
    .out(idx_between_0_depth_plus_0_reg_out),
    .reset(idx_between_0_depth_plus_0_reg_reset),
    .write_en(idx_between_0_depth_plus_0_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_0 (
    .left(index_lt_depth_plus_0_left),
    .out(index_lt_depth_plus_0_out),
    .right(index_lt_depth_plus_0_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_1_min_depth_4_plus_1_reg (
    .clk(idx_between_1_min_depth_4_plus_1_reg_clk),
    .done(idx_between_1_min_depth_4_plus_1_reg_done),
    .in(idx_between_1_min_depth_4_plus_1_reg_in),
    .out(idx_between_1_min_depth_4_plus_1_reg_out),
    .reset(idx_between_1_min_depth_4_plus_1_reg_reset),
    .write_en(idx_between_1_min_depth_4_plus_1_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_1 (
    .left(index_lt_min_depth_4_plus_1_left),
    .out(index_lt_min_depth_4_plus_1_out),
    .right(index_lt_min_depth_4_plus_1_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_1 (
    .left(index_ge_1_left),
    .out(index_ge_1_out),
    .right(index_ge_1_right)
);
std_and # (
    .WIDTH(1)
) idx_between_1_min_depth_4_plus_1_comb (
    .left(idx_between_1_min_depth_4_plus_1_comb_left),
    .out(idx_between_1_min_depth_4_plus_1_comb_out),
    .right(idx_between_1_min_depth_4_plus_1_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_1_depth_plus_1_reg (
    .clk(idx_between_1_depth_plus_1_reg_clk),
    .done(idx_between_1_depth_plus_1_reg_done),
    .in(idx_between_1_depth_plus_1_reg_in),
    .out(idx_between_1_depth_plus_1_reg_out),
    .reset(idx_between_1_depth_plus_1_reg_reset),
    .write_en(idx_between_1_depth_plus_1_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_1 (
    .left(index_lt_depth_plus_1_left),
    .out(index_lt_depth_plus_1_out),
    .right(index_lt_depth_plus_1_right)
);
std_and # (
    .WIDTH(1)
) idx_between_1_depth_plus_1_comb (
    .left(idx_between_1_depth_plus_1_comb_left),
    .out(idx_between_1_depth_plus_1_comb_out),
    .right(idx_between_1_depth_plus_1_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_6_depth_plus_7_reg (
    .clk(idx_between_depth_plus_6_depth_plus_7_reg_clk),
    .done(idx_between_depth_plus_6_depth_plus_7_reg_done),
    .in(idx_between_depth_plus_6_depth_plus_7_reg_in),
    .out(idx_between_depth_plus_6_depth_plus_7_reg_out),
    .reset(idx_between_depth_plus_6_depth_plus_7_reg_reset),
    .write_en(idx_between_depth_plus_6_depth_plus_7_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_6 (
    .left(index_ge_depth_plus_6_left),
    .out(index_ge_depth_plus_6_out),
    .right(index_ge_depth_plus_6_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_6_depth_plus_7_comb (
    .left(idx_between_depth_plus_6_depth_plus_7_comb_left),
    .out(idx_between_depth_plus_6_depth_plus_7_comb_out),
    .right(idx_between_depth_plus_6_depth_plus_7_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_3_min_depth_4_plus_3_reg (
    .clk(idx_between_3_min_depth_4_plus_3_reg_clk),
    .done(idx_between_3_min_depth_4_plus_3_reg_done),
    .in(idx_between_3_min_depth_4_plus_3_reg_in),
    .out(idx_between_3_min_depth_4_plus_3_reg_out),
    .reset(idx_between_3_min_depth_4_plus_3_reg_reset),
    .write_en(idx_between_3_min_depth_4_plus_3_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_3 (
    .left(index_lt_min_depth_4_plus_3_left),
    .out(index_lt_min_depth_4_plus_3_out),
    .right(index_lt_min_depth_4_plus_3_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_3 (
    .left(index_ge_3_left),
    .out(index_ge_3_out),
    .right(index_ge_3_right)
);
std_and # (
    .WIDTH(1)
) idx_between_3_min_depth_4_plus_3_comb (
    .left(idx_between_3_min_depth_4_plus_3_comb_left),
    .out(idx_between_3_min_depth_4_plus_3_comb_out),
    .right(idx_between_3_min_depth_4_plus_3_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_5_depth_plus_6_reg (
    .clk(idx_between_depth_plus_5_depth_plus_6_reg_clk),
    .done(idx_between_depth_plus_5_depth_plus_6_reg_done),
    .in(idx_between_depth_plus_5_depth_plus_6_reg_in),
    .out(idx_between_depth_plus_5_depth_plus_6_reg_out),
    .reset(idx_between_depth_plus_5_depth_plus_6_reg_reset),
    .write_en(idx_between_depth_plus_5_depth_plus_6_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_6 (
    .left(index_lt_depth_plus_6_left),
    .out(index_lt_depth_plus_6_out),
    .right(index_lt_depth_plus_6_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_5 (
    .left(index_ge_depth_plus_5_left),
    .out(index_ge_depth_plus_5_out),
    .right(index_ge_depth_plus_5_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_5_depth_plus_6_comb (
    .left(idx_between_depth_plus_5_depth_plus_6_comb_left),
    .out(idx_between_depth_plus_5_depth_plus_6_comb_out),
    .right(idx_between_depth_plus_5_depth_plus_6_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_2_min_depth_4_plus_2_reg (
    .clk(idx_between_2_min_depth_4_plus_2_reg_clk),
    .done(idx_between_2_min_depth_4_plus_2_reg_done),
    .in(idx_between_2_min_depth_4_plus_2_reg_in),
    .out(idx_between_2_min_depth_4_plus_2_reg_out),
    .reset(idx_between_2_min_depth_4_plus_2_reg_reset),
    .write_en(idx_between_2_min_depth_4_plus_2_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_2 (
    .left(index_lt_min_depth_4_plus_2_left),
    .out(index_lt_min_depth_4_plus_2_out),
    .right(index_lt_min_depth_4_plus_2_right)
);
std_and # (
    .WIDTH(1)
) idx_between_2_min_depth_4_plus_2_comb (
    .left(idx_between_2_min_depth_4_plus_2_comb_left),
    .out(idx_between_2_min_depth_4_plus_2_comb_out),
    .right(idx_between_2_min_depth_4_plus_2_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_6_depth_plus_6_reg (
    .clk(idx_between_6_depth_plus_6_reg_clk),
    .done(idx_between_6_depth_plus_6_reg_done),
    .in(idx_between_6_depth_plus_6_reg_in),
    .out(idx_between_6_depth_plus_6_reg_out),
    .reset(idx_between_6_depth_plus_6_reg_reset),
    .write_en(idx_between_6_depth_plus_6_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_6 (
    .left(index_ge_6_left),
    .out(index_ge_6_out),
    .right(index_ge_6_right)
);
std_and # (
    .WIDTH(1)
) idx_between_6_depth_plus_6_comb (
    .left(idx_between_6_depth_plus_6_comb_left),
    .out(idx_between_6_depth_plus_6_comb_out),
    .right(idx_between_6_depth_plus_6_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_7_depth_plus_8_reg (
    .clk(idx_between_depth_plus_7_depth_plus_8_reg_clk),
    .done(idx_between_depth_plus_7_depth_plus_8_reg_done),
    .in(idx_between_depth_plus_7_depth_plus_8_reg_in),
    .out(idx_between_depth_plus_7_depth_plus_8_reg_out),
    .reset(idx_between_depth_plus_7_depth_plus_8_reg_reset),
    .write_en(idx_between_depth_plus_7_depth_plus_8_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_8 (
    .left(index_lt_depth_plus_8_left),
    .out(index_lt_depth_plus_8_out),
    .right(index_lt_depth_plus_8_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_7 (
    .left(index_ge_depth_plus_7_left),
    .out(index_ge_depth_plus_7_out),
    .right(index_ge_depth_plus_7_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_7_depth_plus_8_comb (
    .left(idx_between_depth_plus_7_depth_plus_8_comb_left),
    .out(idx_between_depth_plus_7_depth_plus_8_comb_out),
    .right(idx_between_depth_plus_7_depth_plus_8_comb_right)
);
std_reg # (
    .WIDTH(1)
) cond (
    .clk(cond_clk),
    .done(cond_done),
    .in(cond_in),
    .out(cond_out),
    .reset(cond_reset),
    .write_en(cond_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire (
    .in(cond_wire_in),
    .out(cond_wire_out)
);
std_reg # (
    .WIDTH(1)
) cond0 (
    .clk(cond0_clk),
    .done(cond0_done),
    .in(cond0_in),
    .out(cond0_out),
    .reset(cond0_reset),
    .write_en(cond0_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire0 (
    .in(cond_wire0_in),
    .out(cond_wire0_out)
);
std_reg # (
    .WIDTH(1)
) cond1 (
    .clk(cond1_clk),
    .done(cond1_done),
    .in(cond1_in),
    .out(cond1_out),
    .reset(cond1_reset),
    .write_en(cond1_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1 (
    .in(cond_wire1_in),
    .out(cond_wire1_out)
);
std_reg # (
    .WIDTH(1)
) cond2 (
    .clk(cond2_clk),
    .done(cond2_done),
    .in(cond2_in),
    .out(cond2_out),
    .reset(cond2_reset),
    .write_en(cond2_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire2 (
    .in(cond_wire2_in),
    .out(cond_wire2_out)
);
std_reg # (
    .WIDTH(1)
) cond3 (
    .clk(cond3_clk),
    .done(cond3_done),
    .in(cond3_in),
    .out(cond3_out),
    .reset(cond3_reset),
    .write_en(cond3_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire3 (
    .in(cond_wire3_in),
    .out(cond_wire3_out)
);
std_reg # (
    .WIDTH(1)
) cond4 (
    .clk(cond4_clk),
    .done(cond4_done),
    .in(cond4_in),
    .out(cond4_out),
    .reset(cond4_reset),
    .write_en(cond4_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire4 (
    .in(cond_wire4_in),
    .out(cond_wire4_out)
);
std_reg # (
    .WIDTH(1)
) cond5 (
    .clk(cond5_clk),
    .done(cond5_done),
    .in(cond5_in),
    .out(cond5_out),
    .reset(cond5_reset),
    .write_en(cond5_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire5 (
    .in(cond_wire5_in),
    .out(cond_wire5_out)
);
std_reg # (
    .WIDTH(1)
) cond6 (
    .clk(cond6_clk),
    .done(cond6_done),
    .in(cond6_in),
    .out(cond6_out),
    .reset(cond6_reset),
    .write_en(cond6_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire6 (
    .in(cond_wire6_in),
    .out(cond_wire6_out)
);
std_reg # (
    .WIDTH(1)
) cond7 (
    .clk(cond7_clk),
    .done(cond7_done),
    .in(cond7_in),
    .out(cond7_out),
    .reset(cond7_reset),
    .write_en(cond7_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire7 (
    .in(cond_wire7_in),
    .out(cond_wire7_out)
);
std_reg # (
    .WIDTH(1)
) cond8 (
    .clk(cond8_clk),
    .done(cond8_done),
    .in(cond8_in),
    .out(cond8_out),
    .reset(cond8_reset),
    .write_en(cond8_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire8 (
    .in(cond_wire8_in),
    .out(cond_wire8_out)
);
std_reg # (
    .WIDTH(1)
) cond9 (
    .clk(cond9_clk),
    .done(cond9_done),
    .in(cond9_in),
    .out(cond9_out),
    .reset(cond9_reset),
    .write_en(cond9_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire9 (
    .in(cond_wire9_in),
    .out(cond_wire9_out)
);
std_reg # (
    .WIDTH(1)
) cond10 (
    .clk(cond10_clk),
    .done(cond10_done),
    .in(cond10_in),
    .out(cond10_out),
    .reset(cond10_reset),
    .write_en(cond10_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire10 (
    .in(cond_wire10_in),
    .out(cond_wire10_out)
);
std_reg # (
    .WIDTH(1)
) cond11 (
    .clk(cond11_clk),
    .done(cond11_done),
    .in(cond11_in),
    .out(cond11_out),
    .reset(cond11_reset),
    .write_en(cond11_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire11 (
    .in(cond_wire11_in),
    .out(cond_wire11_out)
);
std_reg # (
    .WIDTH(1)
) cond12 (
    .clk(cond12_clk),
    .done(cond12_done),
    .in(cond12_in),
    .out(cond12_out),
    .reset(cond12_reset),
    .write_en(cond12_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire12 (
    .in(cond_wire12_in),
    .out(cond_wire12_out)
);
std_reg # (
    .WIDTH(1)
) cond13 (
    .clk(cond13_clk),
    .done(cond13_done),
    .in(cond13_in),
    .out(cond13_out),
    .reset(cond13_reset),
    .write_en(cond13_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire13 (
    .in(cond_wire13_in),
    .out(cond_wire13_out)
);
std_reg # (
    .WIDTH(1)
) cond14 (
    .clk(cond14_clk),
    .done(cond14_done),
    .in(cond14_in),
    .out(cond14_out),
    .reset(cond14_reset),
    .write_en(cond14_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire14 (
    .in(cond_wire14_in),
    .out(cond_wire14_out)
);
std_reg # (
    .WIDTH(1)
) cond15 (
    .clk(cond15_clk),
    .done(cond15_done),
    .in(cond15_in),
    .out(cond15_out),
    .reset(cond15_reset),
    .write_en(cond15_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire15 (
    .in(cond_wire15_in),
    .out(cond_wire15_out)
);
std_reg # (
    .WIDTH(1)
) cond16 (
    .clk(cond16_clk),
    .done(cond16_done),
    .in(cond16_in),
    .out(cond16_out),
    .reset(cond16_reset),
    .write_en(cond16_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire16 (
    .in(cond_wire16_in),
    .out(cond_wire16_out)
);
std_reg # (
    .WIDTH(1)
) fsm (
    .clk(fsm_clk),
    .done(fsm_done),
    .in(fsm_in),
    .out(fsm_out),
    .reset(fsm_reset),
    .write_en(fsm_write_en)
);
undef # (
    .WIDTH(1)
) ud (
    .out(ud_out)
);
std_add # (
    .WIDTH(1)
) adder (
    .left(adder_left),
    .out(adder_out),
    .right(adder_right)
);
undef # (
    .WIDTH(1)
) ud0 (
    .out(ud0_out)
);
std_add # (
    .WIDTH(1)
) adder0 (
    .left(adder0_left),
    .out(adder0_out),
    .right(adder0_right)
);
std_reg # (
    .WIDTH(1)
) signal_reg (
    .clk(signal_reg_clk),
    .done(signal_reg_done),
    .in(signal_reg_in),
    .out(signal_reg_out),
    .reset(signal_reg_reset),
    .write_en(signal_reg_write_en)
);
std_reg # (
    .WIDTH(2)
) fsm0 (
    .clk(fsm0_clk),
    .done(fsm0_done),
    .in(fsm0_in),
    .out(fsm0_out),
    .reset(fsm0_reset),
    .write_en(fsm0_write_en)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_go (
    .in(early_reset_static_par_go_in),
    .out(early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_done (
    .in(early_reset_static_par_done_in),
    .out(early_reset_static_par_done_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par0_go (
    .in(early_reset_static_par0_go_in),
    .out(early_reset_static_par0_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par0_done (
    .in(early_reset_static_par0_done_in),
    .out(early_reset_static_par0_done_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_go (
    .in(wrapper_early_reset_static_par_go_in),
    .out(wrapper_early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_done (
    .in(wrapper_early_reset_static_par_done_in),
    .out(wrapper_early_reset_static_par_done_out)
);
std_wire # (
    .WIDTH(1)
) while_wrapper_early_reset_static_par0_go (
    .in(while_wrapper_early_reset_static_par0_go_in),
    .out(while_wrapper_early_reset_static_par0_go_out)
);
std_wire # (
    .WIDTH(1)
) while_wrapper_early_reset_static_par0_done (
    .in(while_wrapper_early_reset_static_par0_done_in),
    .out(while_wrapper_early_reset_static_par0_done_out)
);
std_wire # (
    .WIDTH(1)
) tdcc_go (
    .in(tdcc_go_in),
    .out(tdcc_go_out)
);
std_wire # (
    .WIDTH(1)
) tdcc_done (
    .in(tdcc_done_in),
    .out(tdcc_done_out)
);
wire _guard0 = 1;
wire _guard1 = cond_wire9_out;
wire _guard2 = early_reset_static_par0_go_out;
wire _guard3 = _guard1 & _guard2;
wire _guard4 = cond_wire9_out;
wire _guard5 = early_reset_static_par0_go_out;
wire _guard6 = _guard4 & _guard5;
wire _guard7 = early_reset_static_par0_go_out;
wire _guard8 = ~_guard0;
wire _guard9 = early_reset_static_par0_go_out;
wire _guard10 = _guard8 & _guard9;
wire _guard11 = cond_wire1_out;
wire _guard12 = early_reset_static_par0_go_out;
wire _guard13 = _guard11 & _guard12;
wire _guard14 = cond_wire1_out;
wire _guard15 = early_reset_static_par0_go_out;
wire _guard16 = _guard14 & _guard15;
wire _guard17 = early_reset_static_par_go_out;
wire _guard18 = early_reset_static_par0_go_out;
wire _guard19 = _guard17 | _guard18;
wire _guard20 = early_reset_static_par0_go_out;
wire _guard21 = early_reset_static_par_go_out;
wire _guard22 = early_reset_static_par0_go_out;
wire _guard23 = early_reset_static_par0_go_out;
wire _guard24 = early_reset_static_par0_go_out;
wire _guard25 = early_reset_static_par0_go_out;
wire _guard26 = early_reset_static_par0_go_out;
wire _guard27 = early_reset_static_par0_go_out;
wire _guard28 = tdcc_done_out;
wire _guard29 = cond_wire_out;
wire _guard30 = early_reset_static_par0_go_out;
wire _guard31 = _guard29 & _guard30;
wire _guard32 = cond_wire13_out;
wire _guard33 = early_reset_static_par0_go_out;
wire _guard34 = _guard32 & _guard33;
wire _guard35 = cond_wire16_out;
wire _guard36 = early_reset_static_par0_go_out;
wire _guard37 = _guard35 & _guard36;
wire _guard38 = cond_wire8_out;
wire _guard39 = early_reset_static_par0_go_out;
wire _guard40 = _guard38 & _guard39;
wire _guard41 = cond_wire3_out;
wire _guard42 = early_reset_static_par0_go_out;
wire _guard43 = _guard41 & _guard42;
wire _guard44 = cond_wire9_out;
wire _guard45 = early_reset_static_par0_go_out;
wire _guard46 = _guard44 & _guard45;
wire _guard47 = cond_wire13_out;
wire _guard48 = early_reset_static_par0_go_out;
wire _guard49 = _guard47 & _guard48;
wire _guard50 = cond_wire16_out;
wire _guard51 = early_reset_static_par0_go_out;
wire _guard52 = _guard50 & _guard51;
wire _guard53 = fsm_out == 1'd0;
wire _guard54 = cond_wire13_out;
wire _guard55 = _guard53 & _guard54;
wire _guard56 = fsm_out == 1'd0;
wire _guard57 = _guard55 & _guard56;
wire _guard58 = fsm_out == 1'd0;
wire _guard59 = cond_wire16_out;
wire _guard60 = _guard58 & _guard59;
wire _guard61 = fsm_out == 1'd0;
wire _guard62 = _guard60 & _guard61;
wire _guard63 = _guard57 | _guard62;
wire _guard64 = early_reset_static_par0_go_out;
wire _guard65 = _guard63 & _guard64;
wire _guard66 = cond_wire_out;
wire _guard67 = early_reset_static_par0_go_out;
wire _guard68 = _guard66 & _guard67;
wire _guard69 = cond_wire4_out;
wire _guard70 = early_reset_static_par0_go_out;
wire _guard71 = _guard69 & _guard70;
wire _guard72 = fsm_out == 1'd0;
wire _guard73 = cond_wire3_out;
wire _guard74 = _guard72 & _guard73;
wire _guard75 = fsm_out == 1'd0;
wire _guard76 = _guard74 & _guard75;
wire _guard77 = fsm_out == 1'd0;
wire _guard78 = cond_wire8_out;
wire _guard79 = _guard77 & _guard78;
wire _guard80 = fsm_out == 1'd0;
wire _guard81 = _guard79 & _guard80;
wire _guard82 = _guard76 | _guard81;
wire _guard83 = early_reset_static_par0_go_out;
wire _guard84 = _guard82 & _guard83;
wire _guard85 = cond_wire3_out;
wire _guard86 = early_reset_static_par0_go_out;
wire _guard87 = _guard85 & _guard86;
wire _guard88 = cond_wire8_out;
wire _guard89 = early_reset_static_par0_go_out;
wire _guard90 = _guard88 & _guard89;
wire _guard91 = early_reset_static_par0_go_out;
wire _guard92 = ~_guard0;
wire _guard93 = early_reset_static_par0_go_out;
wire _guard94 = _guard92 & _guard93;
wire _guard95 = ~_guard0;
wire _guard96 = early_reset_static_par0_go_out;
wire _guard97 = _guard95 & _guard96;
wire _guard98 = early_reset_static_par0_go_out;
wire _guard99 = early_reset_static_par0_go_out;
wire _guard100 = early_reset_static_par0_go_out;
wire _guard101 = early_reset_static_par0_go_out;
wire _guard102 = ~_guard0;
wire _guard103 = early_reset_static_par0_go_out;
wire _guard104 = _guard102 & _guard103;
wire _guard105 = early_reset_static_par0_go_out;
wire _guard106 = ~_guard0;
wire _guard107 = early_reset_static_par0_go_out;
wire _guard108 = _guard106 & _guard107;
wire _guard109 = early_reset_static_par_go_out;
wire _guard110 = early_reset_static_par0_go_out;
wire _guard111 = _guard109 | _guard110;
wire _guard112 = fsm_out != 1'd0;
wire _guard113 = early_reset_static_par_go_out;
wire _guard114 = _guard112 & _guard113;
wire _guard115 = fsm_out == 1'd0;
wire _guard116 = early_reset_static_par_go_out;
wire _guard117 = _guard115 & _guard116;
wire _guard118 = fsm_out == 1'd0;
wire _guard119 = early_reset_static_par0_go_out;
wire _guard120 = _guard118 & _guard119;
wire _guard121 = _guard117 | _guard120;
wire _guard122 = fsm_out != 1'd0;
wire _guard123 = early_reset_static_par0_go_out;
wire _guard124 = _guard122 & _guard123;
wire _guard125 = early_reset_static_par_go_out;
wire _guard126 = early_reset_static_par_go_out;
wire _guard127 = while_wrapper_early_reset_static_par0_go_out;
wire _guard128 = early_reset_static_par_go_out;
wire _guard129 = cond_wire_out;
wire _guard130 = early_reset_static_par0_go_out;
wire _guard131 = _guard129 & _guard130;
wire _guard132 = _guard128 | _guard131;
wire _guard133 = early_reset_static_par_go_out;
wire _guard134 = cond_wire_out;
wire _guard135 = early_reset_static_par0_go_out;
wire _guard136 = _guard134 & _guard135;
wire _guard137 = early_reset_static_par_go_out;
wire _guard138 = early_reset_static_par0_go_out;
wire _guard139 = _guard137 | _guard138;
wire _guard140 = early_reset_static_par_go_out;
wire _guard141 = early_reset_static_par0_go_out;
wire _guard142 = early_reset_static_par0_go_out;
wire _guard143 = early_reset_static_par0_go_out;
wire _guard144 = early_reset_static_par0_go_out;
wire _guard145 = early_reset_static_par0_go_out;
wire _guard146 = early_reset_static_par0_go_out;
wire _guard147 = early_reset_static_par0_go_out;
wire _guard148 = cond_wire7_out;
wire _guard149 = early_reset_static_par0_go_out;
wire _guard150 = _guard148 & _guard149;
wire _guard151 = cond_wire5_out;
wire _guard152 = early_reset_static_par0_go_out;
wire _guard153 = _guard151 & _guard152;
wire _guard154 = fsm_out == 1'd0;
wire _guard155 = cond_wire5_out;
wire _guard156 = _guard154 & _guard155;
wire _guard157 = fsm_out == 1'd0;
wire _guard158 = _guard156 & _guard157;
wire _guard159 = fsm_out == 1'd0;
wire _guard160 = cond_wire7_out;
wire _guard161 = _guard159 & _guard160;
wire _guard162 = fsm_out == 1'd0;
wire _guard163 = _guard161 & _guard162;
wire _guard164 = _guard158 | _guard163;
wire _guard165 = early_reset_static_par0_go_out;
wire _guard166 = _guard164 & _guard165;
wire _guard167 = fsm_out == 1'd0;
wire _guard168 = cond_wire5_out;
wire _guard169 = _guard167 & _guard168;
wire _guard170 = fsm_out == 1'd0;
wire _guard171 = _guard169 & _guard170;
wire _guard172 = fsm_out == 1'd0;
wire _guard173 = cond_wire7_out;
wire _guard174 = _guard172 & _guard173;
wire _guard175 = fsm_out == 1'd0;
wire _guard176 = _guard174 & _guard175;
wire _guard177 = _guard171 | _guard176;
wire _guard178 = early_reset_static_par0_go_out;
wire _guard179 = _guard177 & _guard178;
wire _guard180 = fsm_out == 1'd0;
wire _guard181 = cond_wire5_out;
wire _guard182 = _guard180 & _guard181;
wire _guard183 = fsm_out == 1'd0;
wire _guard184 = _guard182 & _guard183;
wire _guard185 = fsm_out == 1'd0;
wire _guard186 = cond_wire7_out;
wire _guard187 = _guard185 & _guard186;
wire _guard188 = fsm_out == 1'd0;
wire _guard189 = _guard187 & _guard188;
wire _guard190 = _guard184 | _guard189;
wire _guard191 = early_reset_static_par0_go_out;
wire _guard192 = _guard190 & _guard191;
wire _guard193 = early_reset_static_par0_go_out;
wire _guard194 = early_reset_static_par0_go_out;
wire _guard195 = early_reset_static_par0_go_out;
wire _guard196 = early_reset_static_par0_go_out;
wire _guard197 = early_reset_static_par0_go_out;
wire _guard198 = early_reset_static_par0_go_out;
wire _guard199 = early_reset_static_par0_go_out;
wire _guard200 = early_reset_static_par_go_out;
wire _guard201 = early_reset_static_par0_go_out;
wire _guard202 = early_reset_static_par_go_out;
wire _guard203 = cond_wire12_out;
wire _guard204 = early_reset_static_par0_go_out;
wire _guard205 = _guard203 & _guard204;
wire _guard206 = cond_wire10_out;
wire _guard207 = early_reset_static_par0_go_out;
wire _guard208 = _guard206 & _guard207;
wire _guard209 = fsm_out == 1'd0;
wire _guard210 = cond_wire10_out;
wire _guard211 = _guard209 & _guard210;
wire _guard212 = fsm_out == 1'd0;
wire _guard213 = _guard211 & _guard212;
wire _guard214 = fsm_out == 1'd0;
wire _guard215 = cond_wire12_out;
wire _guard216 = _guard214 & _guard215;
wire _guard217 = fsm_out == 1'd0;
wire _guard218 = _guard216 & _guard217;
wire _guard219 = _guard213 | _guard218;
wire _guard220 = early_reset_static_par0_go_out;
wire _guard221 = _guard219 & _guard220;
wire _guard222 = fsm_out == 1'd0;
wire _guard223 = cond_wire10_out;
wire _guard224 = _guard222 & _guard223;
wire _guard225 = fsm_out == 1'd0;
wire _guard226 = _guard224 & _guard225;
wire _guard227 = fsm_out == 1'd0;
wire _guard228 = cond_wire12_out;
wire _guard229 = _guard227 & _guard228;
wire _guard230 = fsm_out == 1'd0;
wire _guard231 = _guard229 & _guard230;
wire _guard232 = _guard226 | _guard231;
wire _guard233 = early_reset_static_par0_go_out;
wire _guard234 = _guard232 & _guard233;
wire _guard235 = fsm_out == 1'd0;
wire _guard236 = cond_wire10_out;
wire _guard237 = _guard235 & _guard236;
wire _guard238 = fsm_out == 1'd0;
wire _guard239 = _guard237 & _guard238;
wire _guard240 = fsm_out == 1'd0;
wire _guard241 = cond_wire12_out;
wire _guard242 = _guard240 & _guard241;
wire _guard243 = fsm_out == 1'd0;
wire _guard244 = _guard242 & _guard243;
wire _guard245 = _guard239 | _guard244;
wire _guard246 = early_reset_static_par0_go_out;
wire _guard247 = _guard245 & _guard246;
wire _guard248 = cond_wire9_out;
wire _guard249 = early_reset_static_par0_go_out;
wire _guard250 = _guard248 & _guard249;
wire _guard251 = cond_wire9_out;
wire _guard252 = early_reset_static_par0_go_out;
wire _guard253 = _guard251 & _guard252;
wire _guard254 = cond_wire11_out;
wire _guard255 = early_reset_static_par0_go_out;
wire _guard256 = _guard254 & _guard255;
wire _guard257 = cond_wire11_out;
wire _guard258 = early_reset_static_par0_go_out;
wire _guard259 = _guard257 & _guard258;
wire _guard260 = early_reset_static_par_go_out;
wire _guard261 = cond_wire4_out;
wire _guard262 = early_reset_static_par0_go_out;
wire _guard263 = _guard261 & _guard262;
wire _guard264 = _guard260 | _guard263;
wire _guard265 = early_reset_static_par_go_out;
wire _guard266 = cond_wire4_out;
wire _guard267 = early_reset_static_par0_go_out;
wire _guard268 = _guard266 & _guard267;
wire _guard269 = early_reset_static_par0_go_out;
wire _guard270 = early_reset_static_par0_go_out;
wire _guard271 = early_reset_static_par0_go_out;
wire _guard272 = early_reset_static_par0_go_out;
wire _guard273 = early_reset_static_par0_go_out;
wire _guard274 = early_reset_static_par0_go_out;
wire _guard275 = cond_wire_out;
wire _guard276 = early_reset_static_par0_go_out;
wire _guard277 = _guard275 & _guard276;
wire _guard278 = cond_wire_out;
wire _guard279 = early_reset_static_par0_go_out;
wire _guard280 = _guard278 & _guard279;
wire _guard281 = early_reset_static_par_go_out;
wire _guard282 = early_reset_static_par0_go_out;
wire _guard283 = _guard281 | _guard282;
wire _guard284 = early_reset_static_par_go_out;
wire _guard285 = early_reset_static_par0_go_out;
wire _guard286 = early_reset_static_par0_go_out;
wire _guard287 = early_reset_static_par0_go_out;
wire _guard288 = wrapper_early_reset_static_par_done_out;
wire _guard289 = ~_guard288;
wire _guard290 = fsm0_out == 2'd0;
wire _guard291 = _guard289 & _guard290;
wire _guard292 = tdcc_go_out;
wire _guard293 = _guard291 & _guard292;
wire _guard294 = early_reset_static_par0_go_out;
wire _guard295 = early_reset_static_par0_go_out;
wire _guard296 = early_reset_static_par_go_out;
wire _guard297 = cond_wire_out;
wire _guard298 = early_reset_static_par0_go_out;
wire _guard299 = _guard297 & _guard298;
wire _guard300 = _guard296 | _guard299;
wire _guard301 = early_reset_static_par_go_out;
wire _guard302 = cond_wire_out;
wire _guard303 = early_reset_static_par0_go_out;
wire _guard304 = _guard302 & _guard303;
wire _guard305 = early_reset_static_par_go_out;
wire _guard306 = cond_wire9_out;
wire _guard307 = early_reset_static_par0_go_out;
wire _guard308 = _guard306 & _guard307;
wire _guard309 = _guard305 | _guard308;
wire _guard310 = cond_wire9_out;
wire _guard311 = early_reset_static_par0_go_out;
wire _guard312 = _guard310 & _guard311;
wire _guard313 = early_reset_static_par_go_out;
wire _guard314 = early_reset_static_par0_go_out;
wire _guard315 = early_reset_static_par0_go_out;
wire _guard316 = early_reset_static_par0_go_out;
wire _guard317 = early_reset_static_par0_go_out;
wire _guard318 = early_reset_static_par0_go_out;
wire _guard319 = early_reset_static_par0_go_out;
wire _guard320 = early_reset_static_par0_go_out;
wire _guard321 = early_reset_static_par0_go_out;
wire _guard322 = early_reset_static_par0_go_out;
wire _guard323 = early_reset_static_par0_go_out;
wire _guard324 = fsm_out == 1'd0;
wire _guard325 = signal_reg_out;
wire _guard326 = _guard324 & _guard325;
wire _guard327 = early_reset_static_par_go_out;
wire _guard328 = early_reset_static_par0_go_out;
wire _guard329 = early_reset_static_par_go_out;
wire _guard330 = early_reset_static_par0_go_out;
wire _guard331 = early_reset_static_par0_go_out;
wire _guard332 = early_reset_static_par0_go_out;
wire _guard333 = early_reset_static_par0_go_out;
wire _guard334 = early_reset_static_par0_go_out;
wire _guard335 = early_reset_static_par0_go_out;
wire _guard336 = early_reset_static_par0_go_out;
wire _guard337 = fsm0_out == 2'd2;
wire _guard338 = fsm0_out == 2'd0;
wire _guard339 = wrapper_early_reset_static_par_done_out;
wire _guard340 = _guard338 & _guard339;
wire _guard341 = tdcc_go_out;
wire _guard342 = _guard340 & _guard341;
wire _guard343 = _guard337 | _guard342;
wire _guard344 = fsm0_out == 2'd1;
wire _guard345 = while_wrapper_early_reset_static_par0_done_out;
wire _guard346 = _guard344 & _guard345;
wire _guard347 = tdcc_go_out;
wire _guard348 = _guard346 & _guard347;
wire _guard349 = _guard343 | _guard348;
wire _guard350 = fsm0_out == 2'd0;
wire _guard351 = wrapper_early_reset_static_par_done_out;
wire _guard352 = _guard350 & _guard351;
wire _guard353 = tdcc_go_out;
wire _guard354 = _guard352 & _guard353;
wire _guard355 = fsm0_out == 2'd2;
wire _guard356 = fsm0_out == 2'd1;
wire _guard357 = while_wrapper_early_reset_static_par0_done_out;
wire _guard358 = _guard356 & _guard357;
wire _guard359 = tdcc_go_out;
wire _guard360 = _guard358 & _guard359;
wire _guard361 = early_reset_static_par0_go_out;
wire _guard362 = early_reset_static_par0_go_out;
wire _guard363 = early_reset_static_par0_go_out;
wire _guard364 = early_reset_static_par0_go_out;
wire _guard365 = early_reset_static_par_go_out;
wire _guard366 = early_reset_static_par0_go_out;
wire _guard367 = _guard365 | _guard366;
wire _guard368 = early_reset_static_par_go_out;
wire _guard369 = early_reset_static_par0_go_out;
wire _guard370 = early_reset_static_par_go_out;
wire _guard371 = early_reset_static_par0_go_out;
wire _guard372 = _guard370 | _guard371;
wire _guard373 = early_reset_static_par0_go_out;
wire _guard374 = early_reset_static_par_go_out;
wire _guard375 = early_reset_static_par0_go_out;
wire _guard376 = early_reset_static_par0_go_out;
wire _guard377 = early_reset_static_par0_go_out;
wire _guard378 = early_reset_static_par0_go_out;
wire _guard379 = early_reset_static_par0_go_out;
wire _guard380 = early_reset_static_par0_go_out;
wire _guard381 = early_reset_static_par0_go_out;
wire _guard382 = ~_guard0;
wire _guard383 = early_reset_static_par0_go_out;
wire _guard384 = _guard382 & _guard383;
wire _guard385 = early_reset_static_par0_go_out;
wire _guard386 = early_reset_static_par0_go_out;
wire _guard387 = early_reset_static_par0_go_out;
wire _guard388 = early_reset_static_par0_go_out;
wire _guard389 = early_reset_static_par_go_out;
wire _guard390 = lt_iter_limit_out;
wire _guard391 = early_reset_static_par_go_out;
wire _guard392 = _guard390 & _guard391;
wire _guard393 = lt_iter_limit_out;
wire _guard394 = ~_guard393;
wire _guard395 = early_reset_static_par_go_out;
wire _guard396 = _guard394 & _guard395;
wire _guard397 = cond_wire4_out;
wire _guard398 = early_reset_static_par0_go_out;
wire _guard399 = _guard397 & _guard398;
wire _guard400 = cond_wire4_out;
wire _guard401 = early_reset_static_par0_go_out;
wire _guard402 = _guard400 & _guard401;
wire _guard403 = early_reset_static_par0_go_out;
wire _guard404 = early_reset_static_par0_go_out;
wire _guard405 = early_reset_static_par_go_out;
wire _guard406 = early_reset_static_par0_go_out;
wire _guard407 = _guard405 | _guard406;
wire _guard408 = early_reset_static_par0_go_out;
wire _guard409 = early_reset_static_par_go_out;
wire _guard410 = early_reset_static_par0_go_out;
wire _guard411 = early_reset_static_par0_go_out;
wire _guard412 = early_reset_static_par0_go_out;
wire _guard413 = early_reset_static_par0_go_out;
wire _guard414 = ~_guard0;
wire _guard415 = early_reset_static_par0_go_out;
wire _guard416 = _guard414 & _guard415;
wire _guard417 = early_reset_static_par0_go_out;
wire _guard418 = early_reset_static_par0_go_out;
wire _guard419 = early_reset_static_par0_go_out;
wire _guard420 = cond_wire6_out;
wire _guard421 = early_reset_static_par0_go_out;
wire _guard422 = _guard420 & _guard421;
wire _guard423 = cond_wire6_out;
wire _guard424 = early_reset_static_par0_go_out;
wire _guard425 = _guard423 & _guard424;
wire _guard426 = cond_wire_out;
wire _guard427 = early_reset_static_par0_go_out;
wire _guard428 = _guard426 & _guard427;
wire _guard429 = cond_wire_out;
wire _guard430 = early_reset_static_par0_go_out;
wire _guard431 = _guard429 & _guard430;
wire _guard432 = cond_wire_out;
wire _guard433 = early_reset_static_par0_go_out;
wire _guard434 = _guard432 & _guard433;
wire _guard435 = cond_wire_out;
wire _guard436 = early_reset_static_par0_go_out;
wire _guard437 = _guard435 & _guard436;
wire _guard438 = early_reset_static_par0_go_out;
wire _guard439 = early_reset_static_par0_go_out;
wire _guard440 = early_reset_static_par0_go_out;
wire _guard441 = early_reset_static_par0_go_out;
wire _guard442 = ~_guard0;
wire _guard443 = early_reset_static_par0_go_out;
wire _guard444 = _guard442 & _guard443;
wire _guard445 = early_reset_static_par0_go_out;
wire _guard446 = ~_guard0;
wire _guard447 = early_reset_static_par0_go_out;
wire _guard448 = _guard446 & _guard447;
wire _guard449 = early_reset_static_par0_go_out;
wire _guard450 = early_reset_static_par0_go_out;
wire _guard451 = early_reset_static_par0_go_out;
wire _guard452 = ~_guard0;
wire _guard453 = early_reset_static_par0_go_out;
wire _guard454 = _guard452 & _guard453;
wire _guard455 = early_reset_static_par0_go_out;
wire _guard456 = fsm_out == 1'd0;
wire _guard457 = signal_reg_out;
wire _guard458 = _guard456 & _guard457;
wire _guard459 = fsm_out == 1'd0;
wire _guard460 = signal_reg_out;
wire _guard461 = ~_guard460;
wire _guard462 = _guard459 & _guard461;
wire _guard463 = wrapper_early_reset_static_par_go_out;
wire _guard464 = _guard462 & _guard463;
wire _guard465 = _guard458 | _guard464;
wire _guard466 = fsm_out == 1'd0;
wire _guard467 = signal_reg_out;
wire _guard468 = ~_guard467;
wire _guard469 = _guard466 & _guard468;
wire _guard470 = wrapper_early_reset_static_par_go_out;
wire _guard471 = _guard469 & _guard470;
wire _guard472 = fsm_out == 1'd0;
wire _guard473 = signal_reg_out;
wire _guard474 = _guard472 & _guard473;
wire _guard475 = early_reset_static_par0_go_out;
wire _guard476 = early_reset_static_par0_go_out;
wire _guard477 = cond_wire4_out;
wire _guard478 = early_reset_static_par0_go_out;
wire _guard479 = _guard477 & _guard478;
wire _guard480 = cond_wire4_out;
wire _guard481 = early_reset_static_par0_go_out;
wire _guard482 = _guard480 & _guard481;
wire _guard483 = early_reset_static_par0_go_out;
wire _guard484 = early_reset_static_par0_go_out;
wire _guard485 = early_reset_static_par0_go_out;
wire _guard486 = early_reset_static_par0_go_out;
wire _guard487 = early_reset_static_par_go_out;
wire _guard488 = early_reset_static_par0_go_out;
wire _guard489 = _guard487 | _guard488;
wire _guard490 = early_reset_static_par_go_out;
wire _guard491 = early_reset_static_par0_go_out;
wire _guard492 = early_reset_static_par_go_out;
wire _guard493 = early_reset_static_par0_go_out;
wire _guard494 = _guard492 | _guard493;
wire _guard495 = early_reset_static_par0_go_out;
wire _guard496 = early_reset_static_par_go_out;
wire _guard497 = early_reset_static_par_go_out;
wire _guard498 = early_reset_static_par0_go_out;
wire _guard499 = _guard497 | _guard498;
wire _guard500 = early_reset_static_par_go_out;
wire _guard501 = early_reset_static_par0_go_out;
wire _guard502 = ~_guard0;
wire _guard503 = early_reset_static_par0_go_out;
wire _guard504 = _guard502 & _guard503;
wire _guard505 = early_reset_static_par0_go_out;
wire _guard506 = ~_guard0;
wire _guard507 = early_reset_static_par0_go_out;
wire _guard508 = _guard506 & _guard507;
wire _guard509 = early_reset_static_par0_go_out;
wire _guard510 = early_reset_static_par0_go_out;
wire _guard511 = early_reset_static_par0_go_out;
wire _guard512 = early_reset_static_par0_go_out;
wire _guard513 = early_reset_static_par0_go_out;
wire _guard514 = cond_wire2_out;
wire _guard515 = early_reset_static_par0_go_out;
wire _guard516 = _guard514 & _guard515;
wire _guard517 = cond_wire0_out;
wire _guard518 = early_reset_static_par0_go_out;
wire _guard519 = _guard517 & _guard518;
wire _guard520 = fsm_out == 1'd0;
wire _guard521 = cond_wire0_out;
wire _guard522 = _guard520 & _guard521;
wire _guard523 = fsm_out == 1'd0;
wire _guard524 = _guard522 & _guard523;
wire _guard525 = fsm_out == 1'd0;
wire _guard526 = cond_wire2_out;
wire _guard527 = _guard525 & _guard526;
wire _guard528 = fsm_out == 1'd0;
wire _guard529 = _guard527 & _guard528;
wire _guard530 = _guard524 | _guard529;
wire _guard531 = early_reset_static_par0_go_out;
wire _guard532 = _guard530 & _guard531;
wire _guard533 = fsm_out == 1'd0;
wire _guard534 = cond_wire0_out;
wire _guard535 = _guard533 & _guard534;
wire _guard536 = fsm_out == 1'd0;
wire _guard537 = _guard535 & _guard536;
wire _guard538 = fsm_out == 1'd0;
wire _guard539 = cond_wire2_out;
wire _guard540 = _guard538 & _guard539;
wire _guard541 = fsm_out == 1'd0;
wire _guard542 = _guard540 & _guard541;
wire _guard543 = _guard537 | _guard542;
wire _guard544 = early_reset_static_par0_go_out;
wire _guard545 = _guard543 & _guard544;
wire _guard546 = fsm_out == 1'd0;
wire _guard547 = cond_wire0_out;
wire _guard548 = _guard546 & _guard547;
wire _guard549 = fsm_out == 1'd0;
wire _guard550 = _guard548 & _guard549;
wire _guard551 = fsm_out == 1'd0;
wire _guard552 = cond_wire2_out;
wire _guard553 = _guard551 & _guard552;
wire _guard554 = fsm_out == 1'd0;
wire _guard555 = _guard553 & _guard554;
wire _guard556 = _guard550 | _guard555;
wire _guard557 = early_reset_static_par0_go_out;
wire _guard558 = _guard556 & _guard557;
wire _guard559 = early_reset_static_par0_go_out;
wire _guard560 = early_reset_static_par0_go_out;
wire _guard561 = early_reset_static_par_go_out;
wire _guard562 = early_reset_static_par0_go_out;
wire _guard563 = _guard561 | _guard562;
wire _guard564 = early_reset_static_par_go_out;
wire _guard565 = early_reset_static_par0_go_out;
wire _guard566 = early_reset_static_par0_go_out;
wire _guard567 = early_reset_static_par0_go_out;
wire _guard568 = early_reset_static_par0_go_out;
wire _guard569 = early_reset_static_par0_go_out;
wire _guard570 = early_reset_static_par_go_out;
wire _guard571 = early_reset_static_par0_go_out;
wire _guard572 = _guard570 | _guard571;
wire _guard573 = early_reset_static_par0_go_out;
wire _guard574 = early_reset_static_par_go_out;
wire _guard575 = early_reset_static_par0_go_out;
wire _guard576 = early_reset_static_par0_go_out;
wire _guard577 = ~_guard0;
wire _guard578 = early_reset_static_par0_go_out;
wire _guard579 = _guard577 & _guard578;
wire _guard580 = early_reset_static_par0_go_out;
wire _guard581 = ~_guard0;
wire _guard582 = early_reset_static_par0_go_out;
wire _guard583 = _guard581 & _guard582;
wire _guard584 = early_reset_static_par0_go_out;
wire _guard585 = early_reset_static_par0_go_out;
wire _guard586 = ~_guard0;
wire _guard587 = early_reset_static_par0_go_out;
wire _guard588 = _guard586 & _guard587;
wire _guard589 = fsm0_out == 2'd2;
wire _guard590 = early_reset_static_par0_go_out;
wire _guard591 = early_reset_static_par0_go_out;
wire _guard592 = early_reset_static_par_go_out;
wire _guard593 = early_reset_static_par0_go_out;
wire _guard594 = _guard592 | _guard593;
wire _guard595 = early_reset_static_par0_go_out;
wire _guard596 = early_reset_static_par_go_out;
wire _guard597 = early_reset_static_par0_go_out;
wire _guard598 = early_reset_static_par0_go_out;
wire _guard599 = early_reset_static_par0_go_out;
wire _guard600 = early_reset_static_par0_go_out;
wire _guard601 = early_reset_static_par0_go_out;
wire _guard602 = early_reset_static_par0_go_out;
wire _guard603 = early_reset_static_par0_go_out;
wire _guard604 = early_reset_static_par0_go_out;
wire _guard605 = ~_guard0;
wire _guard606 = early_reset_static_par0_go_out;
wire _guard607 = _guard605 & _guard606;
wire _guard608 = early_reset_static_par0_go_out;
wire _guard609 = wrapper_early_reset_static_par_go_out;
wire _guard610 = early_reset_static_par_go_out;
wire _guard611 = early_reset_static_par_go_out;
wire _guard612 = early_reset_static_par0_go_out;
wire _guard613 = early_reset_static_par0_go_out;
wire _guard614 = early_reset_static_par0_go_out;
wire _guard615 = early_reset_static_par0_go_out;
wire _guard616 = cond_wire_out;
wire _guard617 = early_reset_static_par0_go_out;
wire _guard618 = _guard616 & _guard617;
wire _guard619 = cond_wire_out;
wire _guard620 = early_reset_static_par0_go_out;
wire _guard621 = _guard619 & _guard620;
wire _guard622 = cond_wire15_out;
wire _guard623 = early_reset_static_par0_go_out;
wire _guard624 = _guard622 & _guard623;
wire _guard625 = cond_wire14_out;
wire _guard626 = early_reset_static_par0_go_out;
wire _guard627 = _guard625 & _guard626;
wire _guard628 = fsm_out == 1'd0;
wire _guard629 = cond_wire14_out;
wire _guard630 = _guard628 & _guard629;
wire _guard631 = fsm_out == 1'd0;
wire _guard632 = _guard630 & _guard631;
wire _guard633 = fsm_out == 1'd0;
wire _guard634 = cond_wire15_out;
wire _guard635 = _guard633 & _guard634;
wire _guard636 = fsm_out == 1'd0;
wire _guard637 = _guard635 & _guard636;
wire _guard638 = _guard632 | _guard637;
wire _guard639 = early_reset_static_par0_go_out;
wire _guard640 = _guard638 & _guard639;
wire _guard641 = fsm_out == 1'd0;
wire _guard642 = cond_wire14_out;
wire _guard643 = _guard641 & _guard642;
wire _guard644 = fsm_out == 1'd0;
wire _guard645 = _guard643 & _guard644;
wire _guard646 = fsm_out == 1'd0;
wire _guard647 = cond_wire15_out;
wire _guard648 = _guard646 & _guard647;
wire _guard649 = fsm_out == 1'd0;
wire _guard650 = _guard648 & _guard649;
wire _guard651 = _guard645 | _guard650;
wire _guard652 = early_reset_static_par0_go_out;
wire _guard653 = _guard651 & _guard652;
wire _guard654 = fsm_out == 1'd0;
wire _guard655 = cond_wire14_out;
wire _guard656 = _guard654 & _guard655;
wire _guard657 = fsm_out == 1'd0;
wire _guard658 = _guard656 & _guard657;
wire _guard659 = fsm_out == 1'd0;
wire _guard660 = cond_wire15_out;
wire _guard661 = _guard659 & _guard660;
wire _guard662 = fsm_out == 1'd0;
wire _guard663 = _guard661 & _guard662;
wire _guard664 = _guard658 | _guard663;
wire _guard665 = early_reset_static_par0_go_out;
wire _guard666 = _guard664 & _guard665;
wire _guard667 = early_reset_static_par0_go_out;
wire _guard668 = early_reset_static_par0_go_out;
wire _guard669 = early_reset_static_par0_go_out;
wire _guard670 = early_reset_static_par0_go_out;
wire _guard671 = early_reset_static_par0_go_out;
wire _guard672 = early_reset_static_par0_go_out;
wire _guard673 = early_reset_static_par0_go_out;
wire _guard674 = ~_guard0;
wire _guard675 = early_reset_static_par0_go_out;
wire _guard676 = _guard674 & _guard675;
wire _guard677 = early_reset_static_par0_go_out;
wire _guard678 = early_reset_static_par0_go_out;
wire _guard679 = early_reset_static_par0_go_out;
wire _guard680 = early_reset_static_par0_go_out;
wire _guard681 = cond_wire1_out;
wire _guard682 = early_reset_static_par0_go_out;
wire _guard683 = _guard681 & _guard682;
wire _guard684 = cond_wire1_out;
wire _guard685 = early_reset_static_par0_go_out;
wire _guard686 = _guard684 & _guard685;
wire _guard687 = early_reset_static_par_go_out;
wire _guard688 = early_reset_static_par0_go_out;
wire _guard689 = _guard687 | _guard688;
wire _guard690 = early_reset_static_par_go_out;
wire _guard691 = early_reset_static_par0_go_out;
wire _guard692 = early_reset_static_par_go_out;
wire _guard693 = early_reset_static_par0_go_out;
wire _guard694 = _guard692 | _guard693;
wire _guard695 = early_reset_static_par0_go_out;
wire _guard696 = early_reset_static_par_go_out;
wire _guard697 = early_reset_static_par0_go_out;
wire _guard698 = early_reset_static_par0_go_out;
wire _guard699 = ~_guard0;
wire _guard700 = early_reset_static_par0_go_out;
wire _guard701 = _guard699 & _guard700;
wire _guard702 = early_reset_static_par0_go_out;
wire _guard703 = while_wrapper_early_reset_static_par0_done_out;
wire _guard704 = ~_guard703;
wire _guard705 = fsm0_out == 2'd1;
wire _guard706 = _guard704 & _guard705;
wire _guard707 = tdcc_go_out;
wire _guard708 = _guard706 & _guard707;
wire _guard709 = cond_reg_out;
wire _guard710 = ~_guard709;
wire _guard711 = fsm_out == 1'd0;
wire _guard712 = _guard710 & _guard711;
assign l1_add_left = 2'd1;
assign l1_add_right = l1_idx_out;
assign cond_wire3_in =
  _guard7 ? idx_between_depth_plus_5_depth_plus_6_reg_out :
  _guard10 ? cond3_out :
  1'd0;
assign top_1_0_write_en = _guard13;
assign top_1_0_clk = clk;
assign top_1_0_reset = reset;
assign top_1_0_in = top_0_0_out;
assign idx_between_depth_plus_6_depth_plus_7_reg_write_en = _guard19;
assign idx_between_depth_plus_6_depth_plus_7_reg_clk = clk;
assign idx_between_depth_plus_6_depth_plus_7_reg_reset = reset;
assign idx_between_depth_plus_6_depth_plus_7_reg_in =
  _guard20 ? idx_between_depth_plus_6_depth_plus_7_comb_out :
  _guard21 ? 1'd0 :
  'x;
assign index_lt_min_depth_4_plus_3_left = idx_add_out;
assign index_lt_min_depth_4_plus_3_right = min_depth_4_plus_3_out;
assign index_lt_depth_plus_6_left = idx_add_out;
assign index_lt_depth_plus_6_right = depth_plus_6_out;
assign index_lt_min_depth_4_plus_2_left = idx_add_out;
assign index_lt_min_depth_4_plus_2_right = min_depth_4_plus_2_out;
assign done = _guard28;
assign l0_addr0 =
  _guard31 ? l0_idx_out :
  2'd0;
assign out_mem_1_addr0 =
  _guard34 ? 32'd0 :
  _guard37 ? 32'd1 :
  32'd0;
assign out_mem_0_write_data =
  _guard40 ? pe_0_1_out :
  _guard43 ? pe_0_0_out :
  32'd0;
assign l1_addr0 =
  _guard46 ? l1_idx_out :
  2'd0;
assign out_mem_1_write_data =
  _guard49 ? pe_1_0_out :
  _guard52 ? pe_1_1_out :
  32'd0;
assign out_mem_1_write_en = _guard65;
assign t0_addr0 =
  _guard68 ? t0_idx_out :
  2'd0;
assign t1_addr0 =
  _guard71 ? t1_idx_out :
  2'd0;
assign out_mem_0_write_en = _guard84;
assign out_mem_0_addr0 =
  _guard87 ? 32'd0 :
  _guard90 ? 32'd1 :
  32'd0;
assign cond_wire0_in =
  _guard91 ? idx_between_1_min_depth_4_plus_1_reg_out :
  _guard94 ? cond0_out :
  1'd0;
assign cond_wire4_in =
  _guard97 ? cond4_out :
  _guard98 ? idx_between_1_depth_plus_1_reg_out :
  1'd0;
assign cond6_write_en = _guard99;
assign cond6_clk = clk;
assign cond6_reset = reset;
assign cond6_in =
  _guard100 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond_wire13_in =
  _guard101 ? idx_between_depth_plus_6_depth_plus_7_reg_out :
  _guard104 ? cond13_out :
  1'd0;
assign cond_wire16_in =
  _guard105 ? idx_between_depth_plus_7_depth_plus_8_reg_out :
  _guard108 ? cond16_out :
  1'd0;
assign fsm_write_en = _guard111;
assign fsm_clk = clk;
assign fsm_reset = reset;
assign fsm_in =
  _guard114 ? adder_out :
  _guard121 ? 1'd0 :
  _guard124 ? adder0_out :
  1'd0;
assign adder_left =
  _guard125 ? fsm_out :
  1'd0;
assign adder_right = _guard126;
assign early_reset_static_par0_go_in = _guard127;
assign l0_idx_write_en = _guard132;
assign l0_idx_clk = clk;
assign l0_idx_reset = reset;
assign l0_idx_in =
  _guard133 ? 2'd0 :
  _guard136 ? l0_add_out :
  'x;
assign idx_between_1_min_depth_4_plus_1_reg_write_en = _guard139;
assign idx_between_1_min_depth_4_plus_1_reg_clk = clk;
assign idx_between_1_min_depth_4_plus_1_reg_reset = reset;
assign idx_between_1_min_depth_4_plus_1_reg_in =
  _guard140 ? 1'd0 :
  _guard141 ? idx_between_1_min_depth_4_plus_1_comb_out :
  'x;
assign idx_between_3_min_depth_4_plus_3_comb_left = index_ge_3_out;
assign idx_between_3_min_depth_4_plus_3_comb_right = index_lt_min_depth_4_plus_3_out;
assign cond11_write_en = _guard144;
assign cond11_clk = clk;
assign cond11_reset = reset;
assign cond11_in =
  _guard145 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond15_write_en = _guard146;
assign cond15_clk = clk;
assign cond15_reset = reset;
assign cond15_in =
  _guard147 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign pe_0_1_mul_ready =
  _guard150 ? 1'd1 :
  _guard153 ? 1'd0 :
  1'd0;
assign pe_0_1_clk = clk;
assign pe_0_1_top =
  _guard166 ? top_0_1_out :
  32'd0;
assign pe_0_1_left =
  _guard179 ? left_0_1_out :
  32'd0;
assign pe_0_1_reset = reset;
assign pe_0_1_go = _guard192;
assign idx_between_5_depth_plus_5_comb_left = index_ge_5_out;
assign idx_between_5_depth_plus_5_comb_right = index_lt_depth_plus_5_out;
assign index_ge_3_left = idx_add_out;
assign index_ge_3_right = 32'd3;
assign cond_write_en = _guard197;
assign cond_clk = clk;
assign cond_reset = reset;
assign cond_in =
  _guard198 ? idx_between_0_depth_plus_0_reg_out :
  1'd0;
assign depth_plus_5_left =
  _guard199 ? depth :
  _guard200 ? 32'd8 :
  'x;
assign depth_plus_5_right =
  _guard201 ? 32'd5 :
  _guard202 ? depth :
  'x;
assign pe_1_0_mul_ready =
  _guard205 ? 1'd1 :
  _guard208 ? 1'd0 :
  1'd0;
assign pe_1_0_clk = clk;
assign pe_1_0_top =
  _guard221 ? top_1_0_out :
  32'd0;
assign pe_1_0_left =
  _guard234 ? left_1_0_out :
  32'd0;
assign pe_1_0_reset = reset;
assign pe_1_0_go = _guard247;
assign left_1_0_write_en = _guard250;
assign left_1_0_clk = clk;
assign left_1_0_reset = reset;
assign left_1_0_in = l1_read_data;
assign left_1_1_write_en = _guard256;
assign left_1_1_clk = clk;
assign left_1_1_reset = reset;
assign left_1_1_in = left_1_0_out;
assign t1_idx_write_en = _guard264;
assign t1_idx_clk = clk;
assign t1_idx_reset = reset;
assign t1_idx_in =
  _guard265 ? 2'd0 :
  _guard268 ? t1_add_out :
  'x;
assign idx_between_depth_plus_6_depth_plus_7_comb_left = index_ge_depth_plus_6_out;
assign idx_between_depth_plus_6_depth_plus_7_comb_right = index_lt_depth_plus_7_out;
assign depth_plus_1_left = depth;
assign depth_plus_1_right = 32'd1;
assign min_depth_4_plus_2_left = min_depth_4_out;
assign min_depth_4_plus_2_right = 32'd2;
assign left_0_0_write_en = _guard277;
assign left_0_0_clk = clk;
assign left_0_0_reset = reset;
assign left_0_0_in = l0_read_data;
assign idx_between_depth_plus_5_depth_plus_6_reg_write_en = _guard283;
assign idx_between_depth_plus_5_depth_plus_6_reg_clk = clk;
assign idx_between_depth_plus_5_depth_plus_6_reg_reset = reset;
assign idx_between_depth_plus_5_depth_plus_6_reg_in =
  _guard284 ? 1'd0 :
  _guard285 ? idx_between_depth_plus_5_depth_plus_6_comb_out :
  'x;
assign index_lt_depth_plus_8_left = idx_add_out;
assign index_lt_depth_plus_8_right = depth_plus_8_out;
assign wrapper_early_reset_static_par_go_in = _guard293;
assign depth_plus_7_left = depth;
assign depth_plus_7_right = 32'd7;
assign t0_idx_write_en = _guard300;
assign t0_idx_clk = clk;
assign t0_idx_reset = reset;
assign t0_idx_in =
  _guard301 ? 2'd0 :
  _guard304 ? t0_add_out :
  'x;
assign l1_idx_write_en = _guard309;
assign l1_idx_clk = clk;
assign l1_idx_reset = reset;
assign l1_idx_in =
  _guard312 ? l1_add_out :
  _guard313 ? 2'd0 :
  'x;
assign idx_add_left = idx_out;
assign idx_add_right = 32'd1;
assign index_ge_7_left = idx_add_out;
assign index_ge_7_right = 32'd7;
assign idx_between_2_min_depth_4_plus_2_comb_left = index_ge_2_out;
assign idx_between_2_min_depth_4_plus_2_comb_right = index_lt_min_depth_4_plus_2_out;
assign cond3_write_en = _guard320;
assign cond3_clk = clk;
assign cond3_reset = reset;
assign cond3_in =
  _guard321 ? idx_between_depth_plus_5_depth_plus_6_reg_out :
  1'd0;
assign cond13_write_en = _guard322;
assign cond13_clk = clk;
assign cond13_reset = reset;
assign cond13_in =
  _guard323 ? idx_between_depth_plus_6_depth_plus_7_reg_out :
  1'd0;
assign wrapper_early_reset_static_par_done_in = _guard326;
assign early_reset_static_par0_done_in = ud0_out;
assign tdcc_go_in = go;
assign lt_iter_limit_left =
  _guard327 ? depth :
  _guard328 ? idx_add_out :
  'x;
assign lt_iter_limit_right =
  _guard329 ? 32'd4 :
  _guard330 ? iter_limit_out :
  'x;
assign idx_between_7_depth_plus_7_comb_left = index_ge_7_out;
assign idx_between_7_depth_plus_7_comb_right = index_lt_depth_plus_7_out;
assign idx_between_6_depth_plus_6_comb_left = index_ge_6_out;
assign idx_between_6_depth_plus_6_comb_right = index_lt_depth_plus_6_out;
assign index_ge_depth_plus_7_left = idx_add_out;
assign index_ge_depth_plus_7_right = depth_plus_7_out;
assign fsm0_write_en = _guard349;
assign fsm0_clk = clk;
assign fsm0_reset = reset;
assign fsm0_in =
  _guard354 ? 2'd1 :
  _guard355 ? 2'd0 :
  _guard360 ? 2'd2 :
  2'd0;
assign depth_plus_0_left = depth;
assign depth_plus_0_right = 32'd0;
assign depth_plus_8_left = depth;
assign depth_plus_8_right = 32'd8;
assign idx_write_en = _guard367;
assign idx_clk = clk;
assign idx_reset = reset;
assign idx_in =
  _guard368 ? 32'd0 :
  _guard369 ? idx_add_out :
  'x;
assign idx_between_7_depth_plus_7_reg_write_en = _guard372;
assign idx_between_7_depth_plus_7_reg_clk = clk;
assign idx_between_7_depth_plus_7_reg_reset = reset;
assign idx_between_7_depth_plus_7_reg_in =
  _guard373 ? idx_between_7_depth_plus_7_comb_out :
  _guard374 ? 1'd0 :
  'x;
assign index_lt_depth_plus_0_left = idx_add_out;
assign index_lt_depth_plus_0_right = depth_plus_0_out;
assign idx_between_1_depth_plus_1_comb_left = index_ge_1_out;
assign idx_between_1_depth_plus_1_comb_right = index_lt_depth_plus_1_out;
assign cond7_write_en = _guard379;
assign cond7_clk = clk;
assign cond7_reset = reset;
assign cond7_in =
  _guard380 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire8_in =
  _guard381 ? idx_between_depth_plus_6_depth_plus_7_reg_out :
  _guard384 ? cond8_out :
  1'd0;
assign cond9_write_en = _guard385;
assign cond9_clk = clk;
assign cond9_reset = reset;
assign cond9_in =
  _guard386 ? idx_between_1_depth_plus_1_reg_out :
  1'd0;
assign cond14_write_en = _guard387;
assign cond14_clk = clk;
assign cond14_reset = reset;
assign cond14_in =
  _guard388 ? idx_between_3_min_depth_4_plus_3_reg_out :
  1'd0;
assign min_depth_4_write_en = _guard389;
assign min_depth_4_clk = clk;
assign min_depth_4_reset = reset;
assign min_depth_4_in =
  _guard392 ? depth :
  _guard396 ? 32'd4 :
  'x;
assign top_0_1_write_en = _guard399;
assign top_0_1_clk = clk;
assign top_0_1_reset = reset;
assign top_0_1_in = t1_read_data;
assign index_ge_1_left = idx_add_out;
assign index_ge_1_right = 32'd1;
assign idx_between_3_min_depth_4_plus_3_reg_write_en = _guard407;
assign idx_between_3_min_depth_4_plus_3_reg_clk = clk;
assign idx_between_3_min_depth_4_plus_3_reg_reset = reset;
assign idx_between_3_min_depth_4_plus_3_reg_in =
  _guard408 ? idx_between_3_min_depth_4_plus_3_comb_out :
  _guard409 ? 1'd0 :
  'x;
assign cond4_write_en = _guard410;
assign cond4_clk = clk;
assign cond4_reset = reset;
assign cond4_in =
  _guard411 ? idx_between_1_depth_plus_1_reg_out :
  1'd0;
assign cond5_write_en = _guard412;
assign cond5_clk = clk;
assign cond5_reset = reset;
assign cond5_in =
  _guard413 ? idx_between_2_min_depth_4_plus_2_reg_out :
  1'd0;
assign cond_wire6_in =
  _guard416 ? cond6_out :
  _guard417 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign adder0_left =
  _guard418 ? fsm_out :
  1'd0;
assign adder0_right = _guard419;
assign early_reset_static_par_done_in = ud_out;
assign top_1_1_write_en = _guard422;
assign top_1_1_clk = clk;
assign top_1_1_reset = reset;
assign top_1_1_in = top_0_1_out;
assign t0_add_left = 2'd1;
assign t0_add_right = t0_idx_out;
assign l0_add_left = 2'd1;
assign l0_add_right = l0_idx_out;
assign idx_between_1_min_depth_4_plus_1_comb_left = index_ge_1_out;
assign idx_between_1_min_depth_4_plus_1_comb_right = index_lt_min_depth_4_plus_1_out;
assign idx_between_depth_plus_7_depth_plus_8_comb_left = index_ge_depth_plus_7_out;
assign idx_between_depth_plus_7_depth_plus_8_comb_right = index_lt_depth_plus_8_out;
assign cond_wire2_in =
  _guard444 ? cond2_out :
  _guard445 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond_wire9_in =
  _guard448 ? cond9_out :
  _guard449 ? idx_between_1_depth_plus_1_reg_out :
  1'd0;
assign cond10_write_en = _guard450;
assign cond10_clk = clk;
assign cond10_reset = reset;
assign cond10_in =
  _guard451 ? idx_between_2_min_depth_4_plus_2_reg_out :
  1'd0;
assign cond_wire11_in =
  _guard454 ? cond11_out :
  _guard455 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign signal_reg_write_en = _guard465;
assign signal_reg_clk = clk;
assign signal_reg_reset = reset;
assign signal_reg_in =
  _guard471 ? 1'd1 :
  _guard474 ? 1'd0 :
  1'd0;
assign depth_plus_6_left = depth;
assign depth_plus_6_right = 32'd6;
assign t1_add_left = 2'd1;
assign t1_add_right = t1_idx_out;
assign index_ge_2_left = idx_add_out;
assign index_ge_2_right = 32'd2;
assign index_lt_depth_plus_7_left = idx_add_out;
assign index_lt_depth_plus_7_right = depth_plus_7_out;
assign idx_between_0_depth_plus_0_reg_write_en = _guard489;
assign idx_between_0_depth_plus_0_reg_clk = clk;
assign idx_between_0_depth_plus_0_reg_reset = reset;
assign idx_between_0_depth_plus_0_reg_in =
  _guard490 ? 1'd1 :
  _guard491 ? index_lt_depth_plus_0_out :
  'x;
assign idx_between_6_depth_plus_6_reg_write_en = _guard494;
assign idx_between_6_depth_plus_6_reg_clk = clk;
assign idx_between_6_depth_plus_6_reg_reset = reset;
assign idx_between_6_depth_plus_6_reg_in =
  _guard495 ? idx_between_6_depth_plus_6_comb_out :
  _guard496 ? 1'd0 :
  'x;
assign idx_between_depth_plus_7_depth_plus_8_reg_write_en = _guard499;
assign idx_between_depth_plus_7_depth_plus_8_reg_clk = clk;
assign idx_between_depth_plus_7_depth_plus_8_reg_reset = reset;
assign idx_between_depth_plus_7_depth_plus_8_reg_in =
  _guard500 ? 1'd0 :
  _guard501 ? idx_between_depth_plus_7_depth_plus_8_comb_out :
  'x;
assign cond_wire_in =
  _guard504 ? cond_out :
  _guard505 ? idx_between_0_depth_plus_0_reg_out :
  1'd0;
assign cond_wire15_in =
  _guard508 ? cond15_out :
  _guard509 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond16_write_en = _guard510;
assign cond16_clk = clk;
assign cond16_reset = reset;
assign cond16_in =
  _guard511 ? idx_between_depth_plus_7_depth_plus_8_reg_out :
  1'd0;
assign depth_plus_2_left = depth;
assign depth_plus_2_right = 32'd2;
assign pe_0_0_mul_ready =
  _guard516 ? 1'd1 :
  _guard519 ? 1'd0 :
  1'd0;
assign pe_0_0_clk = clk;
assign pe_0_0_top =
  _guard532 ? top_0_0_out :
  32'd0;
assign pe_0_0_left =
  _guard545 ? left_0_0_out :
  32'd0;
assign pe_0_0_reset = reset;
assign pe_0_0_go = _guard558;
assign index_ge_5_left = idx_add_out;
assign index_ge_5_right = 32'd5;
assign idx_between_2_depth_plus_2_reg_write_en = _guard563;
assign idx_between_2_depth_plus_2_reg_clk = clk;
assign idx_between_2_depth_plus_2_reg_reset = reset;
assign idx_between_2_depth_plus_2_reg_in =
  _guard564 ? 1'd0 :
  _guard565 ? idx_between_2_depth_plus_2_comb_out :
  'x;
assign idx_between_2_depth_plus_2_comb_left = index_ge_2_out;
assign idx_between_2_depth_plus_2_comb_right = index_lt_depth_plus_2_out;
assign index_ge_depth_plus_6_left = idx_add_out;
assign index_ge_depth_plus_6_right = depth_plus_6_out;
assign idx_between_2_min_depth_4_plus_2_reg_write_en = _guard572;
assign idx_between_2_min_depth_4_plus_2_reg_clk = clk;
assign idx_between_2_min_depth_4_plus_2_reg_reset = reset;
assign idx_between_2_min_depth_4_plus_2_reg_in =
  _guard573 ? idx_between_2_min_depth_4_plus_2_comb_out :
  _guard574 ? 1'd0 :
  'x;
assign cond0_write_en = _guard575;
assign cond0_clk = clk;
assign cond0_reset = reset;
assign cond0_in =
  _guard576 ? idx_between_1_min_depth_4_plus_1_reg_out :
  1'd0;
assign cond_wire7_in =
  _guard579 ? cond7_out :
  _guard580 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire10_in =
  _guard583 ? cond10_out :
  _guard584 ? idx_between_2_min_depth_4_plus_2_reg_out :
  1'd0;
assign cond_wire12_in =
  _guard585 ? idx_between_6_depth_plus_6_reg_out :
  _guard588 ? cond12_out :
  1'd0;
assign tdcc_done_in = _guard589;
assign index_lt_depth_plus_5_left = idx_add_out;
assign index_lt_depth_plus_5_right = depth_plus_5_out;
assign idx_between_1_depth_plus_1_reg_write_en = _guard594;
assign idx_between_1_depth_plus_1_reg_clk = clk;
assign idx_between_1_depth_plus_1_reg_reset = reset;
assign idx_between_1_depth_plus_1_reg_in =
  _guard595 ? idx_between_1_depth_plus_1_comb_out :
  _guard596 ? 1'd0 :
  'x;
assign index_ge_depth_plus_5_left = idx_add_out;
assign index_ge_depth_plus_5_right = depth_plus_5_out;
assign index_ge_6_left = idx_add_out;
assign index_ge_6_right = 32'd6;
assign cond1_write_en = _guard601;
assign cond1_clk = clk;
assign cond1_reset = reset;
assign cond1_in =
  _guard602 ? idx_between_1_depth_plus_1_reg_out :
  1'd0;
assign cond2_write_en = _guard603;
assign cond2_clk = clk;
assign cond2_reset = reset;
assign cond2_in =
  _guard604 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond_wire5_in =
  _guard607 ? cond5_out :
  _guard608 ? idx_between_2_min_depth_4_plus_2_reg_out :
  1'd0;
assign early_reset_static_par_go_in = _guard609;
assign iter_limit_write_en = _guard610;
assign iter_limit_clk = clk;
assign iter_limit_reset = reset;
assign iter_limit_in = depth_plus_5_out;
assign min_depth_4_plus_1_left = min_depth_4_out;
assign min_depth_4_plus_1_right = 32'd1;
assign min_depth_4_plus_3_left = min_depth_4_out;
assign min_depth_4_plus_3_right = 32'd3;
assign top_0_0_write_en = _guard618;
assign top_0_0_clk = clk;
assign top_0_0_reset = reset;
assign top_0_0_in = t0_read_data;
assign pe_1_1_mul_ready =
  _guard624 ? 1'd1 :
  _guard627 ? 1'd0 :
  1'd0;
assign pe_1_1_clk = clk;
assign pe_1_1_top =
  _guard640 ? top_1_1_out :
  32'd0;
assign pe_1_1_left =
  _guard653 ? left_1_1_out :
  32'd0;
assign pe_1_1_reset = reset;
assign pe_1_1_go = _guard666;
assign index_lt_depth_plus_2_left = idx_add_out;
assign index_lt_depth_plus_2_right = depth_plus_2_out;
assign index_lt_min_depth_4_plus_1_left = idx_add_out;
assign index_lt_min_depth_4_plus_1_right = min_depth_4_plus_1_out;
assign idx_between_depth_plus_5_depth_plus_6_comb_left = index_ge_depth_plus_5_out;
assign idx_between_depth_plus_5_depth_plus_6_comb_right = index_lt_depth_plus_6_out;
assign cond_wire1_in =
  _guard673 ? idx_between_1_depth_plus_1_reg_out :
  _guard676 ? cond1_out :
  1'd0;
assign cond8_write_en = _guard677;
assign cond8_clk = clk;
assign cond8_reset = reset;
assign cond8_in =
  _guard678 ? idx_between_depth_plus_6_depth_plus_7_reg_out :
  1'd0;
assign cond12_write_en = _guard679;
assign cond12_clk = clk;
assign cond12_reset = reset;
assign cond12_in =
  _guard680 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign left_0_1_write_en = _guard683;
assign left_0_1_clk = clk;
assign left_0_1_reset = reset;
assign left_0_1_in = left_0_0_out;
assign cond_reg_write_en = _guard689;
assign cond_reg_clk = clk;
assign cond_reg_reset = reset;
assign cond_reg_in =
  _guard690 ? 1'd1 :
  _guard691 ? lt_iter_limit_out :
  'x;
assign idx_between_5_depth_plus_5_reg_write_en = _guard694;
assign idx_between_5_depth_plus_5_reg_clk = clk;
assign idx_between_5_depth_plus_5_reg_reset = reset;
assign idx_between_5_depth_plus_5_reg_in =
  _guard695 ? idx_between_5_depth_plus_5_comb_out :
  _guard696 ? 1'd0 :
  'x;
assign index_lt_depth_plus_1_left = idx_add_out;
assign index_lt_depth_plus_1_right = depth_plus_1_out;
assign cond_wire14_in =
  _guard701 ? cond14_out :
  _guard702 ? idx_between_3_min_depth_4_plus_3_reg_out :
  1'd0;
assign while_wrapper_early_reset_static_par0_go_in = _guard708;
assign while_wrapper_early_reset_static_par0_done_in = _guard712;
// COMPONENT END: systolic_array_comp
endmodule
module main(
  input logic go,
  input logic clk,
  input logic reset,
  output logic done,
  output logic [1:0] t0_addr0,
  output logic [31:0] t0_write_data,
  output logic t0_write_en,
  output logic t0_clk,
  output logic t0_reset,
  input logic [31:0] t0_read_data,
  input logic t0_done,
  output logic [1:0] t1_addr0,
  output logic [31:0] t1_write_data,
  output logic t1_write_en,
  output logic t1_clk,
  output logic t1_reset,
  input logic [31:0] t1_read_data,
  input logic t1_done,
  output logic [1:0] l0_addr0,
  output logic [31:0] l0_write_data,
  output logic l0_write_en,
  output logic l0_clk,
  output logic l0_reset,
  input logic [31:0] l0_read_data,
  input logic l0_done,
  output logic [1:0] l1_addr0,
  output logic [31:0] l1_write_data,
  output logic l1_write_en,
  output logic l1_clk,
  output logic l1_reset,
  input logic [31:0] l1_read_data,
  input logic l1_done,
  output logic [31:0] out_mem_0_addr0,
  output logic [31:0] out_mem_0_write_data,
  output logic out_mem_0_write_en,
  output logic out_mem_0_clk,
  output logic out_mem_0_reset,
  input logic [31:0] out_mem_0_read_data,
  input logic out_mem_0_done,
  output logic [31:0] out_mem_1_addr0,
  output logic [31:0] out_mem_1_write_data,
  output logic out_mem_1_write_en,
  output logic out_mem_1_clk,
  output logic out_mem_1_reset,
  input logic [31:0] out_mem_1_read_data,
  input logic out_mem_1_done
);
// COMPONENT START: main
logic [31:0] systolic_array_depth;
logic [31:0] systolic_array_t0_read_data;
logic [31:0] systolic_array_t1_read_data;
logic [31:0] systolic_array_l0_read_data;
logic [31:0] systolic_array_l1_read_data;
logic [1:0] systolic_array_t0_addr0;
logic [1:0] systolic_array_t1_addr0;
logic [1:0] systolic_array_l0_addr0;
logic [1:0] systolic_array_l1_addr0;
logic [31:0] systolic_array_out_mem_0_addr0;
logic [31:0] systolic_array_out_mem_0_write_data;
logic systolic_array_out_mem_0_write_en;
logic [31:0] systolic_array_out_mem_1_addr0;
logic [31:0] systolic_array_out_mem_1_write_data;
logic systolic_array_out_mem_1_write_en;
logic systolic_array_go;
logic systolic_array_clk;
logic systolic_array_reset;
logic systolic_array_done;
logic invoke0_go_in;
logic invoke0_go_out;
logic invoke0_done_in;
logic invoke0_done_out;
systolic_array_comp systolic_array (
    .clk(systolic_array_clk),
    .depth(systolic_array_depth),
    .done(systolic_array_done),
    .go(systolic_array_go),
    .l0_addr0(systolic_array_l0_addr0),
    .l0_read_data(systolic_array_l0_read_data),
    .l1_addr0(systolic_array_l1_addr0),
    .l1_read_data(systolic_array_l1_read_data),
    .out_mem_0_addr0(systolic_array_out_mem_0_addr0),
    .out_mem_0_write_data(systolic_array_out_mem_0_write_data),
    .out_mem_0_write_en(systolic_array_out_mem_0_write_en),
    .out_mem_1_addr0(systolic_array_out_mem_1_addr0),
    .out_mem_1_write_data(systolic_array_out_mem_1_write_data),
    .out_mem_1_write_en(systolic_array_out_mem_1_write_en),
    .reset(systolic_array_reset),
    .t0_addr0(systolic_array_t0_addr0),
    .t0_read_data(systolic_array_t0_read_data),
    .t1_addr0(systolic_array_t1_addr0),
    .t1_read_data(systolic_array_t1_read_data)
);
std_wire # (
    .WIDTH(1)
) invoke0_go (
    .in(invoke0_go_in),
    .out(invoke0_go_out)
);
std_wire # (
    .WIDTH(1)
) invoke0_done (
    .in(invoke0_done_in),
    .out(invoke0_done_out)
);
wire _guard0 = 1;
wire _guard1 = invoke0_done_out;
wire _guard2 = invoke0_go_out;
wire _guard3 = invoke0_go_out;
wire _guard4 = invoke0_go_out;
wire _guard5 = invoke0_go_out;
wire _guard6 = invoke0_go_out;
wire _guard7 = invoke0_go_out;
wire _guard8 = invoke0_go_out;
wire _guard9 = invoke0_go_out;
wire _guard10 = invoke0_go_out;
wire _guard11 = invoke0_go_out;
wire _guard12 = invoke0_go_out;
wire _guard13 = invoke0_go_out;
wire _guard14 = invoke0_go_out;
wire _guard15 = invoke0_go_out;
wire _guard16 = invoke0_go_out;
wire _guard17 = invoke0_go_out;
assign done = _guard1;
assign t0_reset = reset;
assign l0_addr0 =
  _guard2 ? systolic_array_l0_addr0 :
  2'd0;
assign out_mem_1_addr0 =
  _guard3 ? systolic_array_out_mem_1_addr0 :
  32'd0;
assign out_mem_1_clk = clk;
assign out_mem_0_write_data =
  _guard4 ? systolic_array_out_mem_0_write_data :
  32'd0;
assign t0_clk = clk;
assign out_mem_1_reset = reset;
assign l1_addr0 =
  _guard5 ? systolic_array_l1_addr0 :
  2'd0;
assign l0_reset = reset;
assign out_mem_0_clk = clk;
assign t1_reset = reset;
assign out_mem_1_write_data =
  _guard6 ? systolic_array_out_mem_1_write_data :
  32'd0;
assign out_mem_1_write_en =
  _guard7 ? systolic_array_out_mem_1_write_en :
  1'd0;
assign out_mem_0_reset = reset;
assign t0_addr0 =
  _guard8 ? systolic_array_t0_addr0 :
  2'd0;
assign t1_addr0 =
  _guard9 ? systolic_array_t1_addr0 :
  2'd0;
assign out_mem_0_write_en =
  _guard10 ? systolic_array_out_mem_0_write_en :
  1'd0;
assign t1_clk = clk;
assign l1_reset = reset;
assign out_mem_0_addr0 =
  _guard11 ? systolic_array_out_mem_0_addr0 :
  32'd0;
assign l0_clk = clk;
assign l1_clk = clk;
assign invoke0_go_in = go;
assign invoke0_done_in = systolic_array_done;
assign systolic_array_l1_read_data =
  _guard12 ? l1_read_data :
  32'd0;
assign systolic_array_depth =
  _guard13 ? 32'd2 :
  32'd0;
assign systolic_array_clk = clk;
assign systolic_array_l0_read_data =
  _guard14 ? l0_read_data :
  32'd0;
assign systolic_array_reset = reset;
assign systolic_array_go = _guard15;
assign systolic_array_t1_read_data =
  _guard16 ? t1_read_data :
  32'd0;
assign systolic_array_t0_read_data =
  _guard17 ? t0_read_data :
  32'd0;
// COMPONENT END: main
endmodule

