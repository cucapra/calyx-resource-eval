
/// This is mostly used for testing the static guarantees currently.
/// A realistic implementation would probably take four cycles.
module pipelined_mult (
    input wire clk,
    input wire reset,
    // inputs
    input wire [31:0] left,
    input wire [31:0] right,
    // The input has been committed
    output wire [31:0] out
);

logic [31:0] lt, rt, buff0, buff1, buff2, tmp_prod;

assign out = buff2;
assign tmp_prod = lt * rt;

always_ff @(posedge clk) begin
    if (reset) begin
        lt <= 0;
        rt <= 0;
        buff0 <= 0;
        buff1 <= 0;
        buff2 <= 0;
    end else begin
        lt <= left;
        rt <= right;
        buff0 <= tmp_prod;
        buff1 <= buff0;
        buff2 <= buff1;
    end
end

endmodule

module bb_pipelined_mult(
	               input wire [31:0] left,
	               input wire [31:0] right,
	               output wire [31:0] out,
	               input wire clk
	               );
`ifdef __ICARUS__
   reg [31:0] reg0;
   reg [31:0] reg1;
   reg [31:0] reg2;
   reg [31:0] reg3;
   always @( posedge clk ) begin
      reg0 <= left * right;
      reg1 <= reg0;
      reg2 <= reg1;
      reg3 <= reg2;
   end
   assign out = reg3;
`elsif VERILATOR
   reg [31:0] reg0;
   reg [31:0] reg1;
   reg [31:0] reg2;
   reg [31:0] reg3;
   always @( posedge clk ) begin
      reg0 <= left * right;
      reg1 <= reg0;
      reg2 <= reg1;
      reg3 <= reg2;
   end
   assign out = reg3;
`else
   // mul_uint32 is a black box module generated by Xilinx's IP Core generator.
   // Generation commands are in the synth.tcl file.
   mul_uint32 mul_uint32 (
                   .A(left),
                   .B(right),
                   .P(out),
                   .CLK(clk)
                   );
`endif
endmodule
/* verilator lint_off MULTITOP */
/// =================== Unsigned, Fixed Point =========================
module std_fp_add #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  assign out = left + right;
endmodule

module std_fp_sub #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module std_fp_mult_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16,
    parameter SIGNED = 0
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    input  logic             go,
    input  logic             clk,
    input  logic             reset,
    output logic [WIDTH-1:0] out,
    output logic             done
);
  logic [WIDTH-1:0]          rtmp;
  logic [WIDTH-1:0]          ltmp;
  logic [(WIDTH << 1) - 1:0] out_tmp;
  // Buffer used to walk through the 3 cycles of the pipeline.
  logic done_buf[1:0];

  assign done = done_buf[1];

  assign out = out_tmp[(WIDTH << 1) - INT_WIDTH - 1 : WIDTH - INT_WIDTH];

  // If the done buffer is completely empty and go is high then execution
  // just started.
  logic start;
  assign start = go;

  // Start sending the done signal.
  always_ff @(posedge clk) begin
    if (start)
      done_buf[0] <= 1;
    else
      done_buf[0] <= 0;
  end

  // Push the done signal through the pipeline.
  always_ff @(posedge clk) begin
    if (go) begin
      done_buf[1] <= done_buf[0];
    end else begin
      done_buf[1] <= 0;
    end
  end

  // Register the inputs
  always_ff @(posedge clk) begin
    if (reset) begin
      rtmp <= 0;
      ltmp <= 0;
    end else if (go) begin
      if (SIGNED) begin
        rtmp <= $signed(right);
        ltmp <= $signed(left);
      end else begin
        rtmp <= right;
        ltmp <= left;
      end
    end else begin
      rtmp <= 0;
      ltmp <= 0;
    end

  end

  // Compute the output and save it into out_tmp
  always_ff @(posedge clk) begin
    if (reset) begin
      out_tmp <= 0;
    end else if (go) begin
      if (SIGNED) begin
        // In the first cycle, this performs an invalid computation because
        // ltmp and rtmp only get their actual values in cycle 1
        out_tmp <= $signed(
          { {WIDTH{ltmp[WIDTH-1]}}, ltmp} *
          { {WIDTH{rtmp[WIDTH-1]}}, rtmp}
        );
      end else begin
        out_tmp <= ltmp * rtmp;
      end
    end else begin
      out_tmp <= out_tmp;
    end
  end
endmodule

/* verilator lint_off WIDTH */
module std_fp_div_pipe #(
  parameter WIDTH = 32,
  parameter INT_WIDTH = 16,
  parameter FRAC_WIDTH = 16
) (
    input  logic             go,
    input  logic             clk,
    input  logic             reset,
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out_remainder,
    output logic [WIDTH-1:0] out_quotient,
    output logic             done
);
    localparam ITERATIONS = WIDTH + FRAC_WIDTH;

    logic [WIDTH-1:0] quotient, quotient_next;
    logic [WIDTH:0] acc, acc_next;
    logic [$clog2(ITERATIONS)-1:0] idx;
    logic start, running, finished, dividend_is_zero;

    assign start = go && !running;
    assign dividend_is_zero = start && left == 0;
    assign finished = idx == ITERATIONS - 1 && running;

    always_ff @(posedge clk) begin
      if (reset || finished || dividend_is_zero)
        running <= 0;
      else if (start)
        running <= 1;
      else
        running <= running;
    end

    always_comb begin
      if (acc >= {1'b0, right}) begin
        acc_next = acc - right;
        {acc_next, quotient_next} = {acc_next[WIDTH-1:0], quotient, 1'b1};
      end else begin
        {acc_next, quotient_next} = {acc, quotient} << 1;
      end
    end

    // `done` signaling
    always_ff @(posedge clk) begin
      if (dividend_is_zero || finished)
        done <= 1;
      else
        done <= 0;
    end

    always_ff @(posedge clk) begin
      if (running)
        idx <= idx + 1;
      else
        idx <= 0;
    end

    always_ff @(posedge clk) begin
      if (reset) begin
        out_quotient <= 0;
        out_remainder <= 0;
      end else if (start) begin
        out_quotient <= 0;
        out_remainder <= left;
      end else if (go == 0) begin
        out_quotient <= out_quotient;
        out_remainder <= out_remainder;
      end else if (dividend_is_zero) begin
        out_quotient <= 0;
        out_remainder <= 0;
      end else if (finished) begin
        out_quotient <= quotient_next;
        out_remainder <= out_remainder;
      end else begin
        out_quotient <= out_quotient;
        if (right <= out_remainder)
          out_remainder <= out_remainder - right;
        else
          out_remainder <= out_remainder;
      end
    end

    always_ff @(posedge clk) begin
      if (reset) begin
        acc <= 0;
        quotient <= 0;
      end else if (start) begin
        {acc, quotient} <= {{WIDTH{1'b0}}, left, 1'b0};
      end else begin
        acc <= acc_next;
        quotient <= quotient_next;
      end
    end
endmodule

module std_fp_gt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic             out
);
  assign out = left > right;
endmodule

/// =================== Signed, Fixed Point =========================
module std_fp_sadd #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left + right);
endmodule

module std_fp_ssub #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);

  assign out = $signed(left - right);
endmodule

module std_fp_smult_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  [WIDTH-1:0]              left,
    input  [WIDTH-1:0]              right,
    input  logic                    reset,
    input  logic                    go,
    input  logic                    clk,
    output logic [WIDTH-1:0]        out,
    output logic                    done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(INT_WIDTH),
    .FRAC_WIDTH(FRAC_WIDTH),
    .SIGNED(1)
  ) comp (
    .clk(clk),
    .done(done),
    .reset(reset),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

module std_fp_sdiv_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input                     clk,
    input                     go,
    input                     reset,
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out_quotient,
    output signed [WIDTH-1:0] out_remainder,
    output logic              done
);

  logic signed [WIDTH-1:0] left_abs, right_abs, comp_out_q, comp_out_r, right_save, out_rem_intermediate;

  // Registers to figure out how to transform outputs.
  logic different_signs, left_sign, right_sign;

  // Latch the value of control registers so that their available after
  // go signal becomes low.
  always_ff @(posedge clk) begin
    if (go) begin
      right_save <= right_abs;
      left_sign <= left[WIDTH-1];
      right_sign <= right[WIDTH-1];
    end else begin
      left_sign <= left_sign;
      right_save <= right_save;
      right_sign <= right_sign;
    end
  end

  assign right_abs = right[WIDTH-1] ? -right : right;
  assign left_abs = left[WIDTH-1] ? -left : left;

  assign different_signs = left_sign ^ right_sign;
  assign out_quotient = different_signs ? -comp_out_q : comp_out_q;

  // Remainder is computed as:
  //  t0 = |left| % |right|
  //  t1 = if left * right < 0 and t0 != 0 then |right| - t0 else t0
  //  rem = if right < 0 then -t1 else t1
  assign out_rem_intermediate = different_signs & |comp_out_r ? $signed(right_save - comp_out_r) : comp_out_r;
  assign out_remainder = right_sign ? -out_rem_intermediate : out_rem_intermediate;

  std_fp_div_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(INT_WIDTH),
    .FRAC_WIDTH(FRAC_WIDTH)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left_abs),
    .right(right_abs),
    .out_quotient(comp_out_q),
    .out_remainder(comp_out_r)
  );
endmodule

module std_fp_sgt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic signed [WIDTH-1:0] left,
    input  logic signed [WIDTH-1:0] right,
    output logic signed             out
);
  assign out = $signed(left > right);
endmodule

module std_fp_slt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
   input logic signed [WIDTH-1:0] left,
   input logic signed [WIDTH-1:0] right,
   output logic signed            out
);
  assign out = $signed(left < right);
endmodule

/// =================== Unsigned, Bitnum =========================
module std_mult_pipe #(
    parameter WIDTH = 32
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    input  logic             reset,
    input  logic             go,
    input  logic             clk,
    output logic [WIDTH-1:0] out,
    output logic             done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(WIDTH),
    .FRAC_WIDTH(0),
    .SIGNED(0)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

module std_div_pipe #(
    parameter WIDTH = 32
) (
    input                    reset,
    input                    clk,
    input                    go,
    input        [WIDTH-1:0] left,
    input        [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out_remainder,
    output logic [WIDTH-1:0] out_quotient,
    output logic             done
);

  logic [WIDTH-1:0] dividend;
  logic [(WIDTH-1)*2:0] divisor;
  logic [WIDTH-1:0] quotient;
  logic [WIDTH-1:0] quotient_msk;
  logic start, running, finished, dividend_is_zero;

  assign start = go && !running;
  assign finished = quotient_msk == 0 && running;
  assign dividend_is_zero = start && left == 0;

  always_ff @(posedge clk) begin
    // Early return if the divisor is zero.
    if (finished || dividend_is_zero)
      done <= 1;
    else
      done <= 0;
  end

  always_ff @(posedge clk) begin
    if (reset || finished || dividend_is_zero)
      running <= 0;
    else if (start)
      running <= 1;
    else
      running <= running;
  end

  // Outputs
  always_ff @(posedge clk) begin
    if (dividend_is_zero || start) begin
      out_quotient <= 0;
      out_remainder <= 0;
    end else if (finished) begin
      out_quotient <= quotient;
      out_remainder <= dividend;
    end else begin
      // Otherwise, explicitly latch the values.
      out_quotient <= out_quotient;
      out_remainder <= out_remainder;
    end
  end

  // Calculate the quotient mask.
  always_ff @(posedge clk) begin
    if (start)
      quotient_msk <= 1 << WIDTH - 1;
    else if (running)
      quotient_msk <= quotient_msk >> 1;
    else
      quotient_msk <= quotient_msk;
  end

  // Calculate the quotient.
  always_ff @(posedge clk) begin
    if (start)
      quotient <= 0;
    else if (divisor <= dividend)
      quotient <= quotient | quotient_msk;
    else
      quotient <= quotient;
  end

  // Calculate the dividend.
  always_ff @(posedge clk) begin
    if (start)
      dividend <= left;
    else if (divisor <= dividend)
      dividend <= dividend - divisor;
    else
      dividend <= dividend;
  end

  always_ff @(posedge clk) begin
    if (start) begin
      divisor <= right << WIDTH - 1;
    end else if (finished) begin
      divisor <= 0;
    end else begin
      divisor <= divisor >> 1;
    end
  end

  // Simulation self test against unsynthesizable implementation.
  `ifdef VERILATOR
    logic [WIDTH-1:0] l, r;
    always_ff @(posedge clk) begin
      if (go) begin
        l <= left;
        r <= right;
      end else begin
        l <= l;
        r <= r;
      end
    end

    always @(posedge clk) begin
      if (done && $unsigned(out_remainder) != $unsigned(l % r))
        $error(
          "\nstd_div_pipe (Remainder): Computed and golden outputs do not match!\n",
          "left: %0d", $unsigned(l),
          "  right: %0d\n", $unsigned(r),
          "expected: %0d", $unsigned(l % r),
          "  computed: %0d", $unsigned(out_remainder)
        );

      if (done && $unsigned(out_quotient) != $unsigned(l / r))
        $error(
          "\nstd_div_pipe (Quotient): Computed and golden outputs do not match!\n",
          "left: %0d", $unsigned(l),
          "  right: %0d\n", $unsigned(r),
          "expected: %0d", $unsigned(l / r),
          "  computed: %0d", $unsigned(out_quotient)
        );
    end
  `endif
endmodule

/// =================== Signed, Bitnum =========================
module std_sadd #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left + right);
endmodule

module std_ssub #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left - right);
endmodule

module std_smult_pipe #(
    parameter WIDTH = 32
) (
    input  logic                    reset,
    input  logic                    go,
    input  logic                    clk,
    input  signed       [WIDTH-1:0] left,
    input  signed       [WIDTH-1:0] right,
    output logic signed [WIDTH-1:0] out,
    output logic                    done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(WIDTH),
    .FRAC_WIDTH(0),
    .SIGNED(1)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

/* verilator lint_off WIDTH */
module std_sdiv_pipe #(
    parameter WIDTH = 32
) (
    input                           reset,
    input                           clk,
    input                           go,
    input  logic signed [WIDTH-1:0] left,
    input  logic signed [WIDTH-1:0] right,
    output logic signed [WIDTH-1:0] out_quotient,
    output logic signed [WIDTH-1:0] out_remainder,
    output logic                    done
);

  logic signed [WIDTH-1:0] left_abs, right_abs, comp_out_q, comp_out_r, right_save, out_rem_intermediate;

  // Registers to figure out how to transform outputs.
  logic different_signs, left_sign, right_sign;

  // Latch the value of control registers so that their available after
  // go signal becomes low.
  always_ff @(posedge clk) begin
    if (go) begin
      right_save <= right_abs;
      left_sign <= left[WIDTH-1];
      right_sign <= right[WIDTH-1];
    end else begin
      left_sign <= left_sign;
      right_save <= right_save;
      right_sign <= right_sign;
    end
  end

  assign right_abs = right[WIDTH-1] ? -right : right;
  assign left_abs = left[WIDTH-1] ? -left : left;

  assign different_signs = left_sign ^ right_sign;
  assign out_quotient = different_signs ? -comp_out_q : comp_out_q;

  // Remainder is computed as:
  //  t0 = |left| % |right|
  //  t1 = if left * right < 0 and t0 != 0 then |right| - t0 else t0
  //  rem = if right < 0 then -t1 else t1
  assign out_rem_intermediate = different_signs & |comp_out_r ? $signed(right_save - comp_out_r) : comp_out_r;
  assign out_remainder = right_sign ? -out_rem_intermediate : out_rem_intermediate;

  std_div_pipe #(
    .WIDTH(WIDTH)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left_abs),
    .right(right_abs),
    .out_quotient(comp_out_q),
    .out_remainder(comp_out_r)
  );

  // Simulation self test against unsynthesizable implementation.
  `ifdef VERILATOR
    logic signed [WIDTH-1:0] l, r;
    always_ff @(posedge clk) begin
      if (go) begin
        l <= left;
        r <= right;
      end else begin
        l <= l;
        r <= r;
      end
    end

    always @(posedge clk) begin
      if (done && out_quotient != $signed(l / r))
        $error(
          "\nstd_sdiv_pipe (Quotient): Computed and golden outputs do not match!\n",
          "left: %0d", l,
          "  right: %0d\n", r,
          "expected: %0d", $signed(l / r),
          "  computed: %0d", $signed(out_quotient),
        );
      if (done && out_remainder != $signed(((l % r) + r) % r))
        $error(
          "\nstd_sdiv_pipe (Remainder): Computed and golden outputs do not match!\n",
          "left: %0d", l,
          "  right: %0d\n", r,
          "expected: %0d", $signed(((l % r) + r) % r),
          "  computed: %0d", $signed(out_remainder),
        );
    end
  `endif
endmodule

module std_sgt #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left > right);
endmodule

module std_slt #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left < right);
endmodule

module std_seq #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left == right);
endmodule

module std_sneq #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left != right);
endmodule

module std_sge #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left >= right);
endmodule

module std_sle #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left <= right);
endmodule

module std_slsh #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = left <<< right;
endmodule

module std_srsh #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = left >>> right;
endmodule

/**
 * Core primitives for Calyx.
 * Implements core primitives used by the compiler.
 *
 * Conventions:
 * - All parameter names must be SNAKE_CASE and all caps.
 * - Port names must be snake_case, no caps.
 */
`default_nettype none

module std_slice #(
    parameter IN_WIDTH  = 32,
    parameter OUT_WIDTH = 32
) (
   input wire                   logic [ IN_WIDTH-1:0] in,
   output logic [OUT_WIDTH-1:0] out
);
  assign out = in[OUT_WIDTH-1:0];

  `ifdef VERILATOR
    always_comb begin
      if (IN_WIDTH < OUT_WIDTH)
        $error(
          "std_slice: Input width less than output width\n",
          "IN_WIDTH: %0d", IN_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_pad #(
    parameter IN_WIDTH  = 32,
    parameter OUT_WIDTH = 32
) (
   input wire logic [IN_WIDTH-1:0]  in,
   output logic     [OUT_WIDTH-1:0] out
);
  localparam EXTEND = OUT_WIDTH - IN_WIDTH;
  assign out = { {EXTEND {1'b0}}, in};

  `ifdef VERILATOR
    always_comb begin
      if (IN_WIDTH > OUT_WIDTH)
        $error(
          "std_pad: Output width less than input width\n",
          "IN_WIDTH: %0d", IN_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_cat #(
  parameter LEFT_WIDTH  = 32,
  parameter RIGHT_WIDTH = 32,
  parameter OUT_WIDTH = 64
) (
  input wire logic [LEFT_WIDTH-1:0] left,
  input wire logic [RIGHT_WIDTH-1:0] right,
  output logic [OUT_WIDTH-1:0] out
);
  assign out = {left, right};

  `ifdef VERILATOR
    always_comb begin
      if (LEFT_WIDTH + RIGHT_WIDTH != OUT_WIDTH)
        $error(
          "std_cat: Output width must equal sum of input widths\n",
          "LEFT_WIDTH: %0d", LEFT_WIDTH,
          "RIGHT_WIDTH: %0d", RIGHT_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_not #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] in,
   output logic [WIDTH-1:0] out
);
  assign out = ~in;
endmodule

module std_and #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left & right;
endmodule

module std_or #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left | right;
endmodule

module std_xor #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left ^ right;
endmodule

module std_sub #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module std_gt #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left > right;
endmodule

module std_lt #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left < right;
endmodule

module std_eq #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left == right;
endmodule

module std_neq #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left != right;
endmodule

module std_ge #(
    parameter WIDTH = 32
) (
    input wire   logic [WIDTH-1:0] left,
    input wire   logic [WIDTH-1:0] right,
    output logic out
);
  assign out = left >= right;
endmodule

module std_le #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left <= right;
endmodule

module std_lsh #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left << right;
endmodule

module std_rsh #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left >> right;
endmodule

/// this primitive is intended to be used
/// for lowering purposes (not in source programs)
module std_mux #(
    parameter WIDTH = 32
) (
   input wire               logic cond,
   input wire               logic [WIDTH-1:0] tru,
   input wire               logic [WIDTH-1:0] fal,
   output logic [WIDTH-1:0] out
);
  assign out = cond ? tru : fal;
endmodule

module std_mem_d1 #(
    parameter WIDTH = 32,
    parameter SIZE = 16,
    parameter IDX_SIZE = 4
) (
   input wire                logic [IDX_SIZE-1:0] addr0,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  logic [WIDTH-1:0] mem[SIZE-1:0];

  /* verilator lint_off WIDTH */
  assign read_data = mem[addr0];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= SIZE)
        $error(
          "std_mem_d1: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "SIZE: %0d", SIZE
        );
    end
  `endif
endmodule

module std_mem_d2 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0];

  assign read_data = mem[addr0][addr1];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d2: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d2: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
    end
  `endif
endmodule

module std_mem_d3 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D2_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4,
    parameter D2_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [D2_IDX_SIZE-1:0] addr2,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0][D2_SIZE-1:0];

  assign read_data = mem[addr0][addr1][addr2];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1][addr2] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
      if (addr2 >= D2_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr2: %0d\n", addr2,
          "D2_SIZE: %0d", D2_SIZE
        );
    end
  `endif
endmodule

module std_mem_d4 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D2_SIZE = 16,
    parameter D3_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4,
    parameter D2_IDX_SIZE = 4,
    parameter D3_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [D2_IDX_SIZE-1:0] addr2,
   input wire                logic [D3_IDX_SIZE-1:0] addr3,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0][D2_SIZE-1:0][D3_SIZE-1:0];

  assign read_data = mem[addr0][addr1][addr2][addr3];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1][addr2][addr3] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
      if (addr2 >= D2_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr2: %0d\n", addr2,
          "D2_SIZE: %0d", D2_SIZE
        );
      if (addr3 >= D3_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr3: %0d\n", addr3,
          "D3_SIZE: %0d", D3_SIZE
        );
    end
  `endif
endmodule

`default_nettype wire

module undef #(
    parameter WIDTH = 32
) (
   output logic [WIDTH-1:0] out
);
assign out = 'x;
endmodule

module std_const #(
    parameter WIDTH = 32,
    parameter VALUE = 32
) (
   output logic [WIDTH-1:0] out
);
assign out = VALUE;
endmodule

module std_wire #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] in,
   output logic [WIDTH-1:0] out
);
assign out = in;
endmodule

module std_add #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] left,
   input logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
assign out = left + right;
endmodule

module std_reg #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] in,
   input logic write_en,
   input logic clk,
   input logic reset,
   output logic [WIDTH-1:0] out,
   output logic done
);
always_ff @(posedge clk) begin
    if (reset) begin
       out <= 0;
       done <= 0;
    end else if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module mac_pe(
  input logic [31:0] top,
  input logic [31:0] left,
  input logic mul_ready,
  output logic [31:0] out,
  input logic go,
  input logic clk,
  input logic reset,
  output logic done
);
// COMPONENT START: mac_pe
logic [31:0] acc_in;
logic acc_write_en;
logic acc_clk;
logic acc_reset;
logic [31:0] acc_out;
logic acc_done;
logic [31:0] add_left;
logic [31:0] add_right;
logic [31:0] add_out;
logic mul_clk;
logic [31:0] mul_left;
logic [31:0] mul_right;
logic [31:0] mul_out;
logic fsm_in;
logic fsm_write_en;
logic fsm_clk;
logic fsm_reset;
logic fsm_out;
logic fsm_done;
logic ud_out;
logic adder_left;
logic adder_right;
logic adder_out;
logic signal_reg_in;
logic signal_reg_write_en;
logic signal_reg_clk;
logic signal_reg_reset;
logic signal_reg_out;
logic signal_reg_done;
logic early_reset_static_par_go_in;
logic early_reset_static_par_go_out;
logic early_reset_static_par_done_in;
logic early_reset_static_par_done_out;
logic wrapper_early_reset_static_par_go_in;
logic wrapper_early_reset_static_par_go_out;
logic wrapper_early_reset_static_par_done_in;
logic wrapper_early_reset_static_par_done_out;
std_reg # (
    .WIDTH(32)
) acc (
    .clk(acc_clk),
    .done(acc_done),
    .in(acc_in),
    .out(acc_out),
    .reset(acc_reset),
    .write_en(acc_write_en)
);
std_add # (
    .WIDTH(32)
) add (
    .left(add_left),
    .out(add_out),
    .right(add_right)
);
bb_pipelined_mult mul (
    .clk(mul_clk),
    .left(mul_left),
    .out(mul_out),
    .right(mul_right)
);
std_reg # (
    .WIDTH(1)
) fsm (
    .clk(fsm_clk),
    .done(fsm_done),
    .in(fsm_in),
    .out(fsm_out),
    .reset(fsm_reset),
    .write_en(fsm_write_en)
);
undef # (
    .WIDTH(1)
) ud (
    .out(ud_out)
);
std_add # (
    .WIDTH(1)
) adder (
    .left(adder_left),
    .out(adder_out),
    .right(adder_right)
);
std_reg # (
    .WIDTH(1)
) signal_reg (
    .clk(signal_reg_clk),
    .done(signal_reg_done),
    .in(signal_reg_in),
    .out(signal_reg_out),
    .reset(signal_reg_reset),
    .write_en(signal_reg_write_en)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_go (
    .in(early_reset_static_par_go_in),
    .out(early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_done (
    .in(early_reset_static_par_done_in),
    .out(early_reset_static_par_done_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_go (
    .in(wrapper_early_reset_static_par_go_in),
    .out(wrapper_early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_done (
    .in(wrapper_early_reset_static_par_done_in),
    .out(wrapper_early_reset_static_par_done_out)
);
wire _guard0 = 1;
wire _guard1 = early_reset_static_par_go_out;
wire _guard2 = early_reset_static_par_go_out;
wire _guard3 = wrapper_early_reset_static_par_done_out;
wire _guard4 = early_reset_static_par_go_out;
wire _guard5 = fsm_out != 1'd0;
wire _guard6 = early_reset_static_par_go_out;
wire _guard7 = _guard5 & _guard6;
wire _guard8 = fsm_out == 1'd0;
wire _guard9 = early_reset_static_par_go_out;
wire _guard10 = _guard8 & _guard9;
wire _guard11 = early_reset_static_par_go_out;
wire _guard12 = early_reset_static_par_go_out;
wire _guard13 = fsm_out == 1'd0;
wire _guard14 = signal_reg_out;
wire _guard15 = _guard13 & _guard14;
wire _guard16 = fsm_out == 1'd0;
wire _guard17 = signal_reg_out;
wire _guard18 = _guard16 & _guard17;
wire _guard19 = fsm_out == 1'd0;
wire _guard20 = signal_reg_out;
wire _guard21 = ~_guard20;
wire _guard22 = _guard19 & _guard21;
wire _guard23 = wrapper_early_reset_static_par_go_out;
wire _guard24 = _guard22 & _guard23;
wire _guard25 = _guard18 | _guard24;
wire _guard26 = fsm_out == 1'd0;
wire _guard27 = signal_reg_out;
wire _guard28 = ~_guard27;
wire _guard29 = _guard26 & _guard28;
wire _guard30 = wrapper_early_reset_static_par_go_out;
wire _guard31 = _guard29 & _guard30;
wire _guard32 = fsm_out == 1'd0;
wire _guard33 = signal_reg_out;
wire _guard34 = _guard32 & _guard33;
wire _guard35 = early_reset_static_par_go_out;
wire _guard36 = early_reset_static_par_go_out;
wire _guard37 = early_reset_static_par_go_out;
wire _guard38 = early_reset_static_par_go_out;
wire _guard39 = wrapper_early_reset_static_par_go_out;
assign acc_write_en =
  _guard1 ? mul_ready :
  1'd0;
assign acc_clk = clk;
assign acc_reset = reset;
assign acc_in = add_out;
assign done = _guard3;
assign out = acc_out;
assign fsm_write_en = _guard4;
assign fsm_clk = clk;
assign fsm_reset = reset;
assign fsm_in =
  _guard7 ? adder_out :
  _guard10 ? 1'd0 :
  1'd0;
assign adder_left =
  _guard11 ? fsm_out :
  1'd0;
assign adder_right = _guard12;
assign wrapper_early_reset_static_par_go_in = go;
assign wrapper_early_reset_static_par_done_in = _guard15;
assign early_reset_static_par_done_in = ud_out;
assign signal_reg_write_en = _guard25;
assign signal_reg_clk = clk;
assign signal_reg_reset = reset;
assign signal_reg_in =
  _guard31 ? 1'd1 :
  _guard34 ? 1'd0 :
  1'd0;
assign add_left = acc_out;
assign add_right = mul_out;
assign mul_clk = clk;
assign mul_left =
  _guard37 ? top :
  32'd0;
assign mul_right =
  _guard38 ? left :
  32'd0;
assign early_reset_static_par_go_in = _guard39;
// COMPONENT END: mac_pe
endmodule
module systolic_array_comp(
  input logic [31:0] depth,
  input logic [31:0] t0_read_data,
  input logic [31:0] t1_read_data,
  input logic [31:0] t2_read_data,
  input logic [31:0] t3_read_data,
  input logic [31:0] t4_read_data,
  input logic [31:0] t5_read_data,
  input logic [31:0] t6_read_data,
  input logic [31:0] t7_read_data,
  input logic [31:0] l0_read_data,
  input logic [31:0] l1_read_data,
  input logic [31:0] l2_read_data,
  input logic [31:0] l3_read_data,
  input logic [31:0] l4_read_data,
  input logic [31:0] l5_read_data,
  input logic [31:0] l6_read_data,
  input logic [31:0] l7_read_data,
  output logic [3:0] t0_addr0,
  output logic [3:0] t1_addr0,
  output logic [3:0] t2_addr0,
  output logic [3:0] t3_addr0,
  output logic [3:0] t4_addr0,
  output logic [3:0] t5_addr0,
  output logic [3:0] t6_addr0,
  output logic [3:0] t7_addr0,
  output logic [3:0] l0_addr0,
  output logic [3:0] l1_addr0,
  output logic [3:0] l2_addr0,
  output logic [3:0] l3_addr0,
  output logic [3:0] l4_addr0,
  output logic [3:0] l5_addr0,
  output logic [3:0] l6_addr0,
  output logic [3:0] l7_addr0,
  output logic [31:0] out_mem_0_addr0,
  output logic [31:0] out_mem_0_write_data,
  output logic out_mem_0_write_en,
  output logic [31:0] out_mem_1_addr0,
  output logic [31:0] out_mem_1_write_data,
  output logic out_mem_1_write_en,
  output logic [31:0] out_mem_2_addr0,
  output logic [31:0] out_mem_2_write_data,
  output logic out_mem_2_write_en,
  output logic [31:0] out_mem_3_addr0,
  output logic [31:0] out_mem_3_write_data,
  output logic out_mem_3_write_en,
  output logic [31:0] out_mem_4_addr0,
  output logic [31:0] out_mem_4_write_data,
  output logic out_mem_4_write_en,
  output logic [31:0] out_mem_5_addr0,
  output logic [31:0] out_mem_5_write_data,
  output logic out_mem_5_write_en,
  output logic [31:0] out_mem_6_addr0,
  output logic [31:0] out_mem_6_write_data,
  output logic out_mem_6_write_en,
  output logic [31:0] out_mem_7_addr0,
  output logic [31:0] out_mem_7_write_data,
  output logic out_mem_7_write_en,
  input logic go,
  input logic clk,
  input logic reset,
  output logic done
);
// COMPONENT START: systolic_array_comp
logic [31:0] min_depth_4_in;
logic min_depth_4_write_en;
logic min_depth_4_clk;
logic min_depth_4_reset;
logic [31:0] min_depth_4_out;
logic min_depth_4_done;
logic [31:0] iter_limit_in;
logic iter_limit_write_en;
logic iter_limit_clk;
logic iter_limit_reset;
logic [31:0] iter_limit_out;
logic iter_limit_done;
logic [31:0] depth_plus_16_left;
logic [31:0] depth_plus_16_right;
logic [31:0] depth_plus_16_out;
logic [31:0] depth_plus_17_left;
logic [31:0] depth_plus_17_right;
logic [31:0] depth_plus_17_out;
logic [31:0] depth_plus_12_left;
logic [31:0] depth_plus_12_right;
logic [31:0] depth_plus_12_out;
logic [31:0] depth_plus_13_left;
logic [31:0] depth_plus_13_right;
logic [31:0] depth_plus_13_out;
logic [31:0] depth_plus_8_left;
logic [31:0] depth_plus_8_right;
logic [31:0] depth_plus_8_out;
logic [31:0] depth_plus_9_left;
logic [31:0] depth_plus_9_right;
logic [31:0] depth_plus_9_out;
logic [31:0] min_depth_4_plus_2_left;
logic [31:0] min_depth_4_plus_2_right;
logic [31:0] min_depth_4_plus_2_out;
logic [31:0] depth_plus_2_left;
logic [31:0] depth_plus_2_right;
logic [31:0] depth_plus_2_out;
logic [31:0] depth_plus_18_left;
logic [31:0] depth_plus_18_right;
logic [31:0] depth_plus_18_out;
logic [31:0] depth_plus_11_left;
logic [31:0] depth_plus_11_right;
logic [31:0] depth_plus_11_out;
logic [31:0] min_depth_4_plus_11_left;
logic [31:0] min_depth_4_plus_11_right;
logic [31:0] min_depth_4_plus_11_out;
logic [31:0] depth_plus_14_left;
logic [31:0] depth_plus_14_right;
logic [31:0] depth_plus_14_out;
logic [31:0] depth_plus_7_left;
logic [31:0] depth_plus_7_right;
logic [31:0] depth_plus_7_out;
logic [31:0] min_depth_4_plus_7_left;
logic [31:0] min_depth_4_plus_7_right;
logic [31:0] min_depth_4_plus_7_out;
logic [31:0] depth_plus_19_left;
logic [31:0] depth_plus_19_right;
logic [31:0] depth_plus_19_out;
logic [31:0] depth_plus_3_left;
logic [31:0] depth_plus_3_right;
logic [31:0] depth_plus_3_out;
logic [31:0] min_depth_4_plus_3_left;
logic [31:0] min_depth_4_plus_3_right;
logic [31:0] min_depth_4_plus_3_out;
logic [31:0] min_depth_4_plus_12_left;
logic [31:0] min_depth_4_plus_12_right;
logic [31:0] min_depth_4_plus_12_out;
logic [31:0] depth_plus_5_left;
logic [31:0] depth_plus_5_right;
logic [31:0] depth_plus_5_out;
logic [31:0] depth_plus_6_left;
logic [31:0] depth_plus_6_right;
logic [31:0] depth_plus_6_out;
logic [31:0] depth_plus_15_left;
logic [31:0] depth_plus_15_right;
logic [31:0] depth_plus_15_out;
logic [31:0] depth_plus_10_left;
logic [31:0] depth_plus_10_right;
logic [31:0] depth_plus_10_out;
logic [31:0] min_depth_4_plus_8_left;
logic [31:0] min_depth_4_plus_8_right;
logic [31:0] min_depth_4_plus_8_out;
logic [31:0] depth_plus_20_left;
logic [31:0] depth_plus_20_right;
logic [31:0] depth_plus_20_out;
logic [31:0] min_depth_4_plus_6_left;
logic [31:0] min_depth_4_plus_6_right;
logic [31:0] min_depth_4_plus_6_out;
logic [31:0] min_depth_4_plus_13_left;
logic [31:0] min_depth_4_plus_13_right;
logic [31:0] min_depth_4_plus_13_out;
logic [31:0] depth_plus_4_left;
logic [31:0] depth_plus_4_right;
logic [31:0] depth_plus_4_out;
logic [31:0] min_depth_4_plus_4_left;
logic [31:0] min_depth_4_plus_4_right;
logic [31:0] min_depth_4_plus_4_out;
logic [31:0] min_depth_4_plus_5_left;
logic [31:0] min_depth_4_plus_5_right;
logic [31:0] min_depth_4_plus_5_out;
logic [31:0] min_depth_4_plus_14_left;
logic [31:0] min_depth_4_plus_14_right;
logic [31:0] min_depth_4_plus_14_out;
logic [31:0] depth_plus_0_left;
logic [31:0] depth_plus_0_right;
logic [31:0] depth_plus_0_out;
logic [31:0] min_depth_4_plus_9_left;
logic [31:0] min_depth_4_plus_9_right;
logic [31:0] min_depth_4_plus_9_out;
logic [31:0] depth_plus_1_left;
logic [31:0] depth_plus_1_right;
logic [31:0] depth_plus_1_out;
logic [31:0] min_depth_4_plus_1_left;
logic [31:0] min_depth_4_plus_1_right;
logic [31:0] min_depth_4_plus_1_out;
logic [31:0] min_depth_4_plus_10_left;
logic [31:0] min_depth_4_plus_10_right;
logic [31:0] min_depth_4_plus_10_out;
logic [31:0] min_depth_4_plus_15_left;
logic [31:0] min_depth_4_plus_15_right;
logic [31:0] min_depth_4_plus_15_out;
logic [31:0] pe_0_0_top;
logic [31:0] pe_0_0_left;
logic pe_0_0_mul_ready;
logic [31:0] pe_0_0_out;
logic pe_0_0_go;
logic pe_0_0_clk;
logic pe_0_0_reset;
logic pe_0_0_done;
logic [31:0] top_0_0_in;
logic top_0_0_write_en;
logic top_0_0_clk;
logic top_0_0_reset;
logic [31:0] top_0_0_out;
logic top_0_0_done;
logic [31:0] left_0_0_in;
logic left_0_0_write_en;
logic left_0_0_clk;
logic left_0_0_reset;
logic [31:0] left_0_0_out;
logic left_0_0_done;
logic [31:0] pe_0_1_top;
logic [31:0] pe_0_1_left;
logic pe_0_1_mul_ready;
logic [31:0] pe_0_1_out;
logic pe_0_1_go;
logic pe_0_1_clk;
logic pe_0_1_reset;
logic pe_0_1_done;
logic [31:0] top_0_1_in;
logic top_0_1_write_en;
logic top_0_1_clk;
logic top_0_1_reset;
logic [31:0] top_0_1_out;
logic top_0_1_done;
logic [31:0] left_0_1_in;
logic left_0_1_write_en;
logic left_0_1_clk;
logic left_0_1_reset;
logic [31:0] left_0_1_out;
logic left_0_1_done;
logic [31:0] pe_0_2_top;
logic [31:0] pe_0_2_left;
logic pe_0_2_mul_ready;
logic [31:0] pe_0_2_out;
logic pe_0_2_go;
logic pe_0_2_clk;
logic pe_0_2_reset;
logic pe_0_2_done;
logic [31:0] top_0_2_in;
logic top_0_2_write_en;
logic top_0_2_clk;
logic top_0_2_reset;
logic [31:0] top_0_2_out;
logic top_0_2_done;
logic [31:0] left_0_2_in;
logic left_0_2_write_en;
logic left_0_2_clk;
logic left_0_2_reset;
logic [31:0] left_0_2_out;
logic left_0_2_done;
logic [31:0] pe_0_3_top;
logic [31:0] pe_0_3_left;
logic pe_0_3_mul_ready;
logic [31:0] pe_0_3_out;
logic pe_0_3_go;
logic pe_0_3_clk;
logic pe_0_3_reset;
logic pe_0_3_done;
logic [31:0] top_0_3_in;
logic top_0_3_write_en;
logic top_0_3_clk;
logic top_0_3_reset;
logic [31:0] top_0_3_out;
logic top_0_3_done;
logic [31:0] left_0_3_in;
logic left_0_3_write_en;
logic left_0_3_clk;
logic left_0_3_reset;
logic [31:0] left_0_3_out;
logic left_0_3_done;
logic [31:0] pe_0_4_top;
logic [31:0] pe_0_4_left;
logic pe_0_4_mul_ready;
logic [31:0] pe_0_4_out;
logic pe_0_4_go;
logic pe_0_4_clk;
logic pe_0_4_reset;
logic pe_0_4_done;
logic [31:0] top_0_4_in;
logic top_0_4_write_en;
logic top_0_4_clk;
logic top_0_4_reset;
logic [31:0] top_0_4_out;
logic top_0_4_done;
logic [31:0] left_0_4_in;
logic left_0_4_write_en;
logic left_0_4_clk;
logic left_0_4_reset;
logic [31:0] left_0_4_out;
logic left_0_4_done;
logic [31:0] pe_0_5_top;
logic [31:0] pe_0_5_left;
logic pe_0_5_mul_ready;
logic [31:0] pe_0_5_out;
logic pe_0_5_go;
logic pe_0_5_clk;
logic pe_0_5_reset;
logic pe_0_5_done;
logic [31:0] top_0_5_in;
logic top_0_5_write_en;
logic top_0_5_clk;
logic top_0_5_reset;
logic [31:0] top_0_5_out;
logic top_0_5_done;
logic [31:0] left_0_5_in;
logic left_0_5_write_en;
logic left_0_5_clk;
logic left_0_5_reset;
logic [31:0] left_0_5_out;
logic left_0_5_done;
logic [31:0] pe_0_6_top;
logic [31:0] pe_0_6_left;
logic pe_0_6_mul_ready;
logic [31:0] pe_0_6_out;
logic pe_0_6_go;
logic pe_0_6_clk;
logic pe_0_6_reset;
logic pe_0_6_done;
logic [31:0] top_0_6_in;
logic top_0_6_write_en;
logic top_0_6_clk;
logic top_0_6_reset;
logic [31:0] top_0_6_out;
logic top_0_6_done;
logic [31:0] left_0_6_in;
logic left_0_6_write_en;
logic left_0_6_clk;
logic left_0_6_reset;
logic [31:0] left_0_6_out;
logic left_0_6_done;
logic [31:0] pe_0_7_top;
logic [31:0] pe_0_7_left;
logic pe_0_7_mul_ready;
logic [31:0] pe_0_7_out;
logic pe_0_7_go;
logic pe_0_7_clk;
logic pe_0_7_reset;
logic pe_0_7_done;
logic [31:0] top_0_7_in;
logic top_0_7_write_en;
logic top_0_7_clk;
logic top_0_7_reset;
logic [31:0] top_0_7_out;
logic top_0_7_done;
logic [31:0] left_0_7_in;
logic left_0_7_write_en;
logic left_0_7_clk;
logic left_0_7_reset;
logic [31:0] left_0_7_out;
logic left_0_7_done;
logic [31:0] pe_1_0_top;
logic [31:0] pe_1_0_left;
logic pe_1_0_mul_ready;
logic [31:0] pe_1_0_out;
logic pe_1_0_go;
logic pe_1_0_clk;
logic pe_1_0_reset;
logic pe_1_0_done;
logic [31:0] top_1_0_in;
logic top_1_0_write_en;
logic top_1_0_clk;
logic top_1_0_reset;
logic [31:0] top_1_0_out;
logic top_1_0_done;
logic [31:0] left_1_0_in;
logic left_1_0_write_en;
logic left_1_0_clk;
logic left_1_0_reset;
logic [31:0] left_1_0_out;
logic left_1_0_done;
logic [31:0] pe_1_1_top;
logic [31:0] pe_1_1_left;
logic pe_1_1_mul_ready;
logic [31:0] pe_1_1_out;
logic pe_1_1_go;
logic pe_1_1_clk;
logic pe_1_1_reset;
logic pe_1_1_done;
logic [31:0] top_1_1_in;
logic top_1_1_write_en;
logic top_1_1_clk;
logic top_1_1_reset;
logic [31:0] top_1_1_out;
logic top_1_1_done;
logic [31:0] left_1_1_in;
logic left_1_1_write_en;
logic left_1_1_clk;
logic left_1_1_reset;
logic [31:0] left_1_1_out;
logic left_1_1_done;
logic [31:0] pe_1_2_top;
logic [31:0] pe_1_2_left;
logic pe_1_2_mul_ready;
logic [31:0] pe_1_2_out;
logic pe_1_2_go;
logic pe_1_2_clk;
logic pe_1_2_reset;
logic pe_1_2_done;
logic [31:0] top_1_2_in;
logic top_1_2_write_en;
logic top_1_2_clk;
logic top_1_2_reset;
logic [31:0] top_1_2_out;
logic top_1_2_done;
logic [31:0] left_1_2_in;
logic left_1_2_write_en;
logic left_1_2_clk;
logic left_1_2_reset;
logic [31:0] left_1_2_out;
logic left_1_2_done;
logic [31:0] pe_1_3_top;
logic [31:0] pe_1_3_left;
logic pe_1_3_mul_ready;
logic [31:0] pe_1_3_out;
logic pe_1_3_go;
logic pe_1_3_clk;
logic pe_1_3_reset;
logic pe_1_3_done;
logic [31:0] top_1_3_in;
logic top_1_3_write_en;
logic top_1_3_clk;
logic top_1_3_reset;
logic [31:0] top_1_3_out;
logic top_1_3_done;
logic [31:0] left_1_3_in;
logic left_1_3_write_en;
logic left_1_3_clk;
logic left_1_3_reset;
logic [31:0] left_1_3_out;
logic left_1_3_done;
logic [31:0] pe_1_4_top;
logic [31:0] pe_1_4_left;
logic pe_1_4_mul_ready;
logic [31:0] pe_1_4_out;
logic pe_1_4_go;
logic pe_1_4_clk;
logic pe_1_4_reset;
logic pe_1_4_done;
logic [31:0] top_1_4_in;
logic top_1_4_write_en;
logic top_1_4_clk;
logic top_1_4_reset;
logic [31:0] top_1_4_out;
logic top_1_4_done;
logic [31:0] left_1_4_in;
logic left_1_4_write_en;
logic left_1_4_clk;
logic left_1_4_reset;
logic [31:0] left_1_4_out;
logic left_1_4_done;
logic [31:0] pe_1_5_top;
logic [31:0] pe_1_5_left;
logic pe_1_5_mul_ready;
logic [31:0] pe_1_5_out;
logic pe_1_5_go;
logic pe_1_5_clk;
logic pe_1_5_reset;
logic pe_1_5_done;
logic [31:0] top_1_5_in;
logic top_1_5_write_en;
logic top_1_5_clk;
logic top_1_5_reset;
logic [31:0] top_1_5_out;
logic top_1_5_done;
logic [31:0] left_1_5_in;
logic left_1_5_write_en;
logic left_1_5_clk;
logic left_1_5_reset;
logic [31:0] left_1_5_out;
logic left_1_5_done;
logic [31:0] pe_1_6_top;
logic [31:0] pe_1_6_left;
logic pe_1_6_mul_ready;
logic [31:0] pe_1_6_out;
logic pe_1_6_go;
logic pe_1_6_clk;
logic pe_1_6_reset;
logic pe_1_6_done;
logic [31:0] top_1_6_in;
logic top_1_6_write_en;
logic top_1_6_clk;
logic top_1_6_reset;
logic [31:0] top_1_6_out;
logic top_1_6_done;
logic [31:0] left_1_6_in;
logic left_1_6_write_en;
logic left_1_6_clk;
logic left_1_6_reset;
logic [31:0] left_1_6_out;
logic left_1_6_done;
logic [31:0] pe_1_7_top;
logic [31:0] pe_1_7_left;
logic pe_1_7_mul_ready;
logic [31:0] pe_1_7_out;
logic pe_1_7_go;
logic pe_1_7_clk;
logic pe_1_7_reset;
logic pe_1_7_done;
logic [31:0] top_1_7_in;
logic top_1_7_write_en;
logic top_1_7_clk;
logic top_1_7_reset;
logic [31:0] top_1_7_out;
logic top_1_7_done;
logic [31:0] left_1_7_in;
logic left_1_7_write_en;
logic left_1_7_clk;
logic left_1_7_reset;
logic [31:0] left_1_7_out;
logic left_1_7_done;
logic [31:0] pe_2_0_top;
logic [31:0] pe_2_0_left;
logic pe_2_0_mul_ready;
logic [31:0] pe_2_0_out;
logic pe_2_0_go;
logic pe_2_0_clk;
logic pe_2_0_reset;
logic pe_2_0_done;
logic [31:0] top_2_0_in;
logic top_2_0_write_en;
logic top_2_0_clk;
logic top_2_0_reset;
logic [31:0] top_2_0_out;
logic top_2_0_done;
logic [31:0] left_2_0_in;
logic left_2_0_write_en;
logic left_2_0_clk;
logic left_2_0_reset;
logic [31:0] left_2_0_out;
logic left_2_0_done;
logic [31:0] pe_2_1_top;
logic [31:0] pe_2_1_left;
logic pe_2_1_mul_ready;
logic [31:0] pe_2_1_out;
logic pe_2_1_go;
logic pe_2_1_clk;
logic pe_2_1_reset;
logic pe_2_1_done;
logic [31:0] top_2_1_in;
logic top_2_1_write_en;
logic top_2_1_clk;
logic top_2_1_reset;
logic [31:0] top_2_1_out;
logic top_2_1_done;
logic [31:0] left_2_1_in;
logic left_2_1_write_en;
logic left_2_1_clk;
logic left_2_1_reset;
logic [31:0] left_2_1_out;
logic left_2_1_done;
logic [31:0] pe_2_2_top;
logic [31:0] pe_2_2_left;
logic pe_2_2_mul_ready;
logic [31:0] pe_2_2_out;
logic pe_2_2_go;
logic pe_2_2_clk;
logic pe_2_2_reset;
logic pe_2_2_done;
logic [31:0] top_2_2_in;
logic top_2_2_write_en;
logic top_2_2_clk;
logic top_2_2_reset;
logic [31:0] top_2_2_out;
logic top_2_2_done;
logic [31:0] left_2_2_in;
logic left_2_2_write_en;
logic left_2_2_clk;
logic left_2_2_reset;
logic [31:0] left_2_2_out;
logic left_2_2_done;
logic [31:0] pe_2_3_top;
logic [31:0] pe_2_3_left;
logic pe_2_3_mul_ready;
logic [31:0] pe_2_3_out;
logic pe_2_3_go;
logic pe_2_3_clk;
logic pe_2_3_reset;
logic pe_2_3_done;
logic [31:0] top_2_3_in;
logic top_2_3_write_en;
logic top_2_3_clk;
logic top_2_3_reset;
logic [31:0] top_2_3_out;
logic top_2_3_done;
logic [31:0] left_2_3_in;
logic left_2_3_write_en;
logic left_2_3_clk;
logic left_2_3_reset;
logic [31:0] left_2_3_out;
logic left_2_3_done;
logic [31:0] pe_2_4_top;
logic [31:0] pe_2_4_left;
logic pe_2_4_mul_ready;
logic [31:0] pe_2_4_out;
logic pe_2_4_go;
logic pe_2_4_clk;
logic pe_2_4_reset;
logic pe_2_4_done;
logic [31:0] top_2_4_in;
logic top_2_4_write_en;
logic top_2_4_clk;
logic top_2_4_reset;
logic [31:0] top_2_4_out;
logic top_2_4_done;
logic [31:0] left_2_4_in;
logic left_2_4_write_en;
logic left_2_4_clk;
logic left_2_4_reset;
logic [31:0] left_2_4_out;
logic left_2_4_done;
logic [31:0] pe_2_5_top;
logic [31:0] pe_2_5_left;
logic pe_2_5_mul_ready;
logic [31:0] pe_2_5_out;
logic pe_2_5_go;
logic pe_2_5_clk;
logic pe_2_5_reset;
logic pe_2_5_done;
logic [31:0] top_2_5_in;
logic top_2_5_write_en;
logic top_2_5_clk;
logic top_2_5_reset;
logic [31:0] top_2_5_out;
logic top_2_5_done;
logic [31:0] left_2_5_in;
logic left_2_5_write_en;
logic left_2_5_clk;
logic left_2_5_reset;
logic [31:0] left_2_5_out;
logic left_2_5_done;
logic [31:0] pe_2_6_top;
logic [31:0] pe_2_6_left;
logic pe_2_6_mul_ready;
logic [31:0] pe_2_6_out;
logic pe_2_6_go;
logic pe_2_6_clk;
logic pe_2_6_reset;
logic pe_2_6_done;
logic [31:0] top_2_6_in;
logic top_2_6_write_en;
logic top_2_6_clk;
logic top_2_6_reset;
logic [31:0] top_2_6_out;
logic top_2_6_done;
logic [31:0] left_2_6_in;
logic left_2_6_write_en;
logic left_2_6_clk;
logic left_2_6_reset;
logic [31:0] left_2_6_out;
logic left_2_6_done;
logic [31:0] pe_2_7_top;
logic [31:0] pe_2_7_left;
logic pe_2_7_mul_ready;
logic [31:0] pe_2_7_out;
logic pe_2_7_go;
logic pe_2_7_clk;
logic pe_2_7_reset;
logic pe_2_7_done;
logic [31:0] top_2_7_in;
logic top_2_7_write_en;
logic top_2_7_clk;
logic top_2_7_reset;
logic [31:0] top_2_7_out;
logic top_2_7_done;
logic [31:0] left_2_7_in;
logic left_2_7_write_en;
logic left_2_7_clk;
logic left_2_7_reset;
logic [31:0] left_2_7_out;
logic left_2_7_done;
logic [31:0] pe_3_0_top;
logic [31:0] pe_3_0_left;
logic pe_3_0_mul_ready;
logic [31:0] pe_3_0_out;
logic pe_3_0_go;
logic pe_3_0_clk;
logic pe_3_0_reset;
logic pe_3_0_done;
logic [31:0] top_3_0_in;
logic top_3_0_write_en;
logic top_3_0_clk;
logic top_3_0_reset;
logic [31:0] top_3_0_out;
logic top_3_0_done;
logic [31:0] left_3_0_in;
logic left_3_0_write_en;
logic left_3_0_clk;
logic left_3_0_reset;
logic [31:0] left_3_0_out;
logic left_3_0_done;
logic [31:0] pe_3_1_top;
logic [31:0] pe_3_1_left;
logic pe_3_1_mul_ready;
logic [31:0] pe_3_1_out;
logic pe_3_1_go;
logic pe_3_1_clk;
logic pe_3_1_reset;
logic pe_3_1_done;
logic [31:0] top_3_1_in;
logic top_3_1_write_en;
logic top_3_1_clk;
logic top_3_1_reset;
logic [31:0] top_3_1_out;
logic top_3_1_done;
logic [31:0] left_3_1_in;
logic left_3_1_write_en;
logic left_3_1_clk;
logic left_3_1_reset;
logic [31:0] left_3_1_out;
logic left_3_1_done;
logic [31:0] pe_3_2_top;
logic [31:0] pe_3_2_left;
logic pe_3_2_mul_ready;
logic [31:0] pe_3_2_out;
logic pe_3_2_go;
logic pe_3_2_clk;
logic pe_3_2_reset;
logic pe_3_2_done;
logic [31:0] top_3_2_in;
logic top_3_2_write_en;
logic top_3_2_clk;
logic top_3_2_reset;
logic [31:0] top_3_2_out;
logic top_3_2_done;
logic [31:0] left_3_2_in;
logic left_3_2_write_en;
logic left_3_2_clk;
logic left_3_2_reset;
logic [31:0] left_3_2_out;
logic left_3_2_done;
logic [31:0] pe_3_3_top;
logic [31:0] pe_3_3_left;
logic pe_3_3_mul_ready;
logic [31:0] pe_3_3_out;
logic pe_3_3_go;
logic pe_3_3_clk;
logic pe_3_3_reset;
logic pe_3_3_done;
logic [31:0] top_3_3_in;
logic top_3_3_write_en;
logic top_3_3_clk;
logic top_3_3_reset;
logic [31:0] top_3_3_out;
logic top_3_3_done;
logic [31:0] left_3_3_in;
logic left_3_3_write_en;
logic left_3_3_clk;
logic left_3_3_reset;
logic [31:0] left_3_3_out;
logic left_3_3_done;
logic [31:0] pe_3_4_top;
logic [31:0] pe_3_4_left;
logic pe_3_4_mul_ready;
logic [31:0] pe_3_4_out;
logic pe_3_4_go;
logic pe_3_4_clk;
logic pe_3_4_reset;
logic pe_3_4_done;
logic [31:0] top_3_4_in;
logic top_3_4_write_en;
logic top_3_4_clk;
logic top_3_4_reset;
logic [31:0] top_3_4_out;
logic top_3_4_done;
logic [31:0] left_3_4_in;
logic left_3_4_write_en;
logic left_3_4_clk;
logic left_3_4_reset;
logic [31:0] left_3_4_out;
logic left_3_4_done;
logic [31:0] pe_3_5_top;
logic [31:0] pe_3_5_left;
logic pe_3_5_mul_ready;
logic [31:0] pe_3_5_out;
logic pe_3_5_go;
logic pe_3_5_clk;
logic pe_3_5_reset;
logic pe_3_5_done;
logic [31:0] top_3_5_in;
logic top_3_5_write_en;
logic top_3_5_clk;
logic top_3_5_reset;
logic [31:0] top_3_5_out;
logic top_3_5_done;
logic [31:0] left_3_5_in;
logic left_3_5_write_en;
logic left_3_5_clk;
logic left_3_5_reset;
logic [31:0] left_3_5_out;
logic left_3_5_done;
logic [31:0] pe_3_6_top;
logic [31:0] pe_3_6_left;
logic pe_3_6_mul_ready;
logic [31:0] pe_3_6_out;
logic pe_3_6_go;
logic pe_3_6_clk;
logic pe_3_6_reset;
logic pe_3_6_done;
logic [31:0] top_3_6_in;
logic top_3_6_write_en;
logic top_3_6_clk;
logic top_3_6_reset;
logic [31:0] top_3_6_out;
logic top_3_6_done;
logic [31:0] left_3_6_in;
logic left_3_6_write_en;
logic left_3_6_clk;
logic left_3_6_reset;
logic [31:0] left_3_6_out;
logic left_3_6_done;
logic [31:0] pe_3_7_top;
logic [31:0] pe_3_7_left;
logic pe_3_7_mul_ready;
logic [31:0] pe_3_7_out;
logic pe_3_7_go;
logic pe_3_7_clk;
logic pe_3_7_reset;
logic pe_3_7_done;
logic [31:0] top_3_7_in;
logic top_3_7_write_en;
logic top_3_7_clk;
logic top_3_7_reset;
logic [31:0] top_3_7_out;
logic top_3_7_done;
logic [31:0] left_3_7_in;
logic left_3_7_write_en;
logic left_3_7_clk;
logic left_3_7_reset;
logic [31:0] left_3_7_out;
logic left_3_7_done;
logic [31:0] pe_4_0_top;
logic [31:0] pe_4_0_left;
logic pe_4_0_mul_ready;
logic [31:0] pe_4_0_out;
logic pe_4_0_go;
logic pe_4_0_clk;
logic pe_4_0_reset;
logic pe_4_0_done;
logic [31:0] top_4_0_in;
logic top_4_0_write_en;
logic top_4_0_clk;
logic top_4_0_reset;
logic [31:0] top_4_0_out;
logic top_4_0_done;
logic [31:0] left_4_0_in;
logic left_4_0_write_en;
logic left_4_0_clk;
logic left_4_0_reset;
logic [31:0] left_4_0_out;
logic left_4_0_done;
logic [31:0] pe_4_1_top;
logic [31:0] pe_4_1_left;
logic pe_4_1_mul_ready;
logic [31:0] pe_4_1_out;
logic pe_4_1_go;
logic pe_4_1_clk;
logic pe_4_1_reset;
logic pe_4_1_done;
logic [31:0] top_4_1_in;
logic top_4_1_write_en;
logic top_4_1_clk;
logic top_4_1_reset;
logic [31:0] top_4_1_out;
logic top_4_1_done;
logic [31:0] left_4_1_in;
logic left_4_1_write_en;
logic left_4_1_clk;
logic left_4_1_reset;
logic [31:0] left_4_1_out;
logic left_4_1_done;
logic [31:0] pe_4_2_top;
logic [31:0] pe_4_2_left;
logic pe_4_2_mul_ready;
logic [31:0] pe_4_2_out;
logic pe_4_2_go;
logic pe_4_2_clk;
logic pe_4_2_reset;
logic pe_4_2_done;
logic [31:0] top_4_2_in;
logic top_4_2_write_en;
logic top_4_2_clk;
logic top_4_2_reset;
logic [31:0] top_4_2_out;
logic top_4_2_done;
logic [31:0] left_4_2_in;
logic left_4_2_write_en;
logic left_4_2_clk;
logic left_4_2_reset;
logic [31:0] left_4_2_out;
logic left_4_2_done;
logic [31:0] pe_4_3_top;
logic [31:0] pe_4_3_left;
logic pe_4_3_mul_ready;
logic [31:0] pe_4_3_out;
logic pe_4_3_go;
logic pe_4_3_clk;
logic pe_4_3_reset;
logic pe_4_3_done;
logic [31:0] top_4_3_in;
logic top_4_3_write_en;
logic top_4_3_clk;
logic top_4_3_reset;
logic [31:0] top_4_3_out;
logic top_4_3_done;
logic [31:0] left_4_3_in;
logic left_4_3_write_en;
logic left_4_3_clk;
logic left_4_3_reset;
logic [31:0] left_4_3_out;
logic left_4_3_done;
logic [31:0] pe_4_4_top;
logic [31:0] pe_4_4_left;
logic pe_4_4_mul_ready;
logic [31:0] pe_4_4_out;
logic pe_4_4_go;
logic pe_4_4_clk;
logic pe_4_4_reset;
logic pe_4_4_done;
logic [31:0] top_4_4_in;
logic top_4_4_write_en;
logic top_4_4_clk;
logic top_4_4_reset;
logic [31:0] top_4_4_out;
logic top_4_4_done;
logic [31:0] left_4_4_in;
logic left_4_4_write_en;
logic left_4_4_clk;
logic left_4_4_reset;
logic [31:0] left_4_4_out;
logic left_4_4_done;
logic [31:0] pe_4_5_top;
logic [31:0] pe_4_5_left;
logic pe_4_5_mul_ready;
logic [31:0] pe_4_5_out;
logic pe_4_5_go;
logic pe_4_5_clk;
logic pe_4_5_reset;
logic pe_4_5_done;
logic [31:0] top_4_5_in;
logic top_4_5_write_en;
logic top_4_5_clk;
logic top_4_5_reset;
logic [31:0] top_4_5_out;
logic top_4_5_done;
logic [31:0] left_4_5_in;
logic left_4_5_write_en;
logic left_4_5_clk;
logic left_4_5_reset;
logic [31:0] left_4_5_out;
logic left_4_5_done;
logic [31:0] pe_4_6_top;
logic [31:0] pe_4_6_left;
logic pe_4_6_mul_ready;
logic [31:0] pe_4_6_out;
logic pe_4_6_go;
logic pe_4_6_clk;
logic pe_4_6_reset;
logic pe_4_6_done;
logic [31:0] top_4_6_in;
logic top_4_6_write_en;
logic top_4_6_clk;
logic top_4_6_reset;
logic [31:0] top_4_6_out;
logic top_4_6_done;
logic [31:0] left_4_6_in;
logic left_4_6_write_en;
logic left_4_6_clk;
logic left_4_6_reset;
logic [31:0] left_4_6_out;
logic left_4_6_done;
logic [31:0] pe_4_7_top;
logic [31:0] pe_4_7_left;
logic pe_4_7_mul_ready;
logic [31:0] pe_4_7_out;
logic pe_4_7_go;
logic pe_4_7_clk;
logic pe_4_7_reset;
logic pe_4_7_done;
logic [31:0] top_4_7_in;
logic top_4_7_write_en;
logic top_4_7_clk;
logic top_4_7_reset;
logic [31:0] top_4_7_out;
logic top_4_7_done;
logic [31:0] left_4_7_in;
logic left_4_7_write_en;
logic left_4_7_clk;
logic left_4_7_reset;
logic [31:0] left_4_7_out;
logic left_4_7_done;
logic [31:0] pe_5_0_top;
logic [31:0] pe_5_0_left;
logic pe_5_0_mul_ready;
logic [31:0] pe_5_0_out;
logic pe_5_0_go;
logic pe_5_0_clk;
logic pe_5_0_reset;
logic pe_5_0_done;
logic [31:0] top_5_0_in;
logic top_5_0_write_en;
logic top_5_0_clk;
logic top_5_0_reset;
logic [31:0] top_5_0_out;
logic top_5_0_done;
logic [31:0] left_5_0_in;
logic left_5_0_write_en;
logic left_5_0_clk;
logic left_5_0_reset;
logic [31:0] left_5_0_out;
logic left_5_0_done;
logic [31:0] pe_5_1_top;
logic [31:0] pe_5_1_left;
logic pe_5_1_mul_ready;
logic [31:0] pe_5_1_out;
logic pe_5_1_go;
logic pe_5_1_clk;
logic pe_5_1_reset;
logic pe_5_1_done;
logic [31:0] top_5_1_in;
logic top_5_1_write_en;
logic top_5_1_clk;
logic top_5_1_reset;
logic [31:0] top_5_1_out;
logic top_5_1_done;
logic [31:0] left_5_1_in;
logic left_5_1_write_en;
logic left_5_1_clk;
logic left_5_1_reset;
logic [31:0] left_5_1_out;
logic left_5_1_done;
logic [31:0] pe_5_2_top;
logic [31:0] pe_5_2_left;
logic pe_5_2_mul_ready;
logic [31:0] pe_5_2_out;
logic pe_5_2_go;
logic pe_5_2_clk;
logic pe_5_2_reset;
logic pe_5_2_done;
logic [31:0] top_5_2_in;
logic top_5_2_write_en;
logic top_5_2_clk;
logic top_5_2_reset;
logic [31:0] top_5_2_out;
logic top_5_2_done;
logic [31:0] left_5_2_in;
logic left_5_2_write_en;
logic left_5_2_clk;
logic left_5_2_reset;
logic [31:0] left_5_2_out;
logic left_5_2_done;
logic [31:0] pe_5_3_top;
logic [31:0] pe_5_3_left;
logic pe_5_3_mul_ready;
logic [31:0] pe_5_3_out;
logic pe_5_3_go;
logic pe_5_3_clk;
logic pe_5_3_reset;
logic pe_5_3_done;
logic [31:0] top_5_3_in;
logic top_5_3_write_en;
logic top_5_3_clk;
logic top_5_3_reset;
logic [31:0] top_5_3_out;
logic top_5_3_done;
logic [31:0] left_5_3_in;
logic left_5_3_write_en;
logic left_5_3_clk;
logic left_5_3_reset;
logic [31:0] left_5_3_out;
logic left_5_3_done;
logic [31:0] pe_5_4_top;
logic [31:0] pe_5_4_left;
logic pe_5_4_mul_ready;
logic [31:0] pe_5_4_out;
logic pe_5_4_go;
logic pe_5_4_clk;
logic pe_5_4_reset;
logic pe_5_4_done;
logic [31:0] top_5_4_in;
logic top_5_4_write_en;
logic top_5_4_clk;
logic top_5_4_reset;
logic [31:0] top_5_4_out;
logic top_5_4_done;
logic [31:0] left_5_4_in;
logic left_5_4_write_en;
logic left_5_4_clk;
logic left_5_4_reset;
logic [31:0] left_5_4_out;
logic left_5_4_done;
logic [31:0] pe_5_5_top;
logic [31:0] pe_5_5_left;
logic pe_5_5_mul_ready;
logic [31:0] pe_5_5_out;
logic pe_5_5_go;
logic pe_5_5_clk;
logic pe_5_5_reset;
logic pe_5_5_done;
logic [31:0] top_5_5_in;
logic top_5_5_write_en;
logic top_5_5_clk;
logic top_5_5_reset;
logic [31:0] top_5_5_out;
logic top_5_5_done;
logic [31:0] left_5_5_in;
logic left_5_5_write_en;
logic left_5_5_clk;
logic left_5_5_reset;
logic [31:0] left_5_5_out;
logic left_5_5_done;
logic [31:0] pe_5_6_top;
logic [31:0] pe_5_6_left;
logic pe_5_6_mul_ready;
logic [31:0] pe_5_6_out;
logic pe_5_6_go;
logic pe_5_6_clk;
logic pe_5_6_reset;
logic pe_5_6_done;
logic [31:0] top_5_6_in;
logic top_5_6_write_en;
logic top_5_6_clk;
logic top_5_6_reset;
logic [31:0] top_5_6_out;
logic top_5_6_done;
logic [31:0] left_5_6_in;
logic left_5_6_write_en;
logic left_5_6_clk;
logic left_5_6_reset;
logic [31:0] left_5_6_out;
logic left_5_6_done;
logic [31:0] pe_5_7_top;
logic [31:0] pe_5_7_left;
logic pe_5_7_mul_ready;
logic [31:0] pe_5_7_out;
logic pe_5_7_go;
logic pe_5_7_clk;
logic pe_5_7_reset;
logic pe_5_7_done;
logic [31:0] top_5_7_in;
logic top_5_7_write_en;
logic top_5_7_clk;
logic top_5_7_reset;
logic [31:0] top_5_7_out;
logic top_5_7_done;
logic [31:0] left_5_7_in;
logic left_5_7_write_en;
logic left_5_7_clk;
logic left_5_7_reset;
logic [31:0] left_5_7_out;
logic left_5_7_done;
logic [31:0] pe_6_0_top;
logic [31:0] pe_6_0_left;
logic pe_6_0_mul_ready;
logic [31:0] pe_6_0_out;
logic pe_6_0_go;
logic pe_6_0_clk;
logic pe_6_0_reset;
logic pe_6_0_done;
logic [31:0] top_6_0_in;
logic top_6_0_write_en;
logic top_6_0_clk;
logic top_6_0_reset;
logic [31:0] top_6_0_out;
logic top_6_0_done;
logic [31:0] left_6_0_in;
logic left_6_0_write_en;
logic left_6_0_clk;
logic left_6_0_reset;
logic [31:0] left_6_0_out;
logic left_6_0_done;
logic [31:0] pe_6_1_top;
logic [31:0] pe_6_1_left;
logic pe_6_1_mul_ready;
logic [31:0] pe_6_1_out;
logic pe_6_1_go;
logic pe_6_1_clk;
logic pe_6_1_reset;
logic pe_6_1_done;
logic [31:0] top_6_1_in;
logic top_6_1_write_en;
logic top_6_1_clk;
logic top_6_1_reset;
logic [31:0] top_6_1_out;
logic top_6_1_done;
logic [31:0] left_6_1_in;
logic left_6_1_write_en;
logic left_6_1_clk;
logic left_6_1_reset;
logic [31:0] left_6_1_out;
logic left_6_1_done;
logic [31:0] pe_6_2_top;
logic [31:0] pe_6_2_left;
logic pe_6_2_mul_ready;
logic [31:0] pe_6_2_out;
logic pe_6_2_go;
logic pe_6_2_clk;
logic pe_6_2_reset;
logic pe_6_2_done;
logic [31:0] top_6_2_in;
logic top_6_2_write_en;
logic top_6_2_clk;
logic top_6_2_reset;
logic [31:0] top_6_2_out;
logic top_6_2_done;
logic [31:0] left_6_2_in;
logic left_6_2_write_en;
logic left_6_2_clk;
logic left_6_2_reset;
logic [31:0] left_6_2_out;
logic left_6_2_done;
logic [31:0] pe_6_3_top;
logic [31:0] pe_6_3_left;
logic pe_6_3_mul_ready;
logic [31:0] pe_6_3_out;
logic pe_6_3_go;
logic pe_6_3_clk;
logic pe_6_3_reset;
logic pe_6_3_done;
logic [31:0] top_6_3_in;
logic top_6_3_write_en;
logic top_6_3_clk;
logic top_6_3_reset;
logic [31:0] top_6_3_out;
logic top_6_3_done;
logic [31:0] left_6_3_in;
logic left_6_3_write_en;
logic left_6_3_clk;
logic left_6_3_reset;
logic [31:0] left_6_3_out;
logic left_6_3_done;
logic [31:0] pe_6_4_top;
logic [31:0] pe_6_4_left;
logic pe_6_4_mul_ready;
logic [31:0] pe_6_4_out;
logic pe_6_4_go;
logic pe_6_4_clk;
logic pe_6_4_reset;
logic pe_6_4_done;
logic [31:0] top_6_4_in;
logic top_6_4_write_en;
logic top_6_4_clk;
logic top_6_4_reset;
logic [31:0] top_6_4_out;
logic top_6_4_done;
logic [31:0] left_6_4_in;
logic left_6_4_write_en;
logic left_6_4_clk;
logic left_6_4_reset;
logic [31:0] left_6_4_out;
logic left_6_4_done;
logic [31:0] pe_6_5_top;
logic [31:0] pe_6_5_left;
logic pe_6_5_mul_ready;
logic [31:0] pe_6_5_out;
logic pe_6_5_go;
logic pe_6_5_clk;
logic pe_6_5_reset;
logic pe_6_5_done;
logic [31:0] top_6_5_in;
logic top_6_5_write_en;
logic top_6_5_clk;
logic top_6_5_reset;
logic [31:0] top_6_5_out;
logic top_6_5_done;
logic [31:0] left_6_5_in;
logic left_6_5_write_en;
logic left_6_5_clk;
logic left_6_5_reset;
logic [31:0] left_6_5_out;
logic left_6_5_done;
logic [31:0] pe_6_6_top;
logic [31:0] pe_6_6_left;
logic pe_6_6_mul_ready;
logic [31:0] pe_6_6_out;
logic pe_6_6_go;
logic pe_6_6_clk;
logic pe_6_6_reset;
logic pe_6_6_done;
logic [31:0] top_6_6_in;
logic top_6_6_write_en;
logic top_6_6_clk;
logic top_6_6_reset;
logic [31:0] top_6_6_out;
logic top_6_6_done;
logic [31:0] left_6_6_in;
logic left_6_6_write_en;
logic left_6_6_clk;
logic left_6_6_reset;
logic [31:0] left_6_6_out;
logic left_6_6_done;
logic [31:0] pe_6_7_top;
logic [31:0] pe_6_7_left;
logic pe_6_7_mul_ready;
logic [31:0] pe_6_7_out;
logic pe_6_7_go;
logic pe_6_7_clk;
logic pe_6_7_reset;
logic pe_6_7_done;
logic [31:0] top_6_7_in;
logic top_6_7_write_en;
logic top_6_7_clk;
logic top_6_7_reset;
logic [31:0] top_6_7_out;
logic top_6_7_done;
logic [31:0] left_6_7_in;
logic left_6_7_write_en;
logic left_6_7_clk;
logic left_6_7_reset;
logic [31:0] left_6_7_out;
logic left_6_7_done;
logic [31:0] pe_7_0_top;
logic [31:0] pe_7_0_left;
logic pe_7_0_mul_ready;
logic [31:0] pe_7_0_out;
logic pe_7_0_go;
logic pe_7_0_clk;
logic pe_7_0_reset;
logic pe_7_0_done;
logic [31:0] top_7_0_in;
logic top_7_0_write_en;
logic top_7_0_clk;
logic top_7_0_reset;
logic [31:0] top_7_0_out;
logic top_7_0_done;
logic [31:0] left_7_0_in;
logic left_7_0_write_en;
logic left_7_0_clk;
logic left_7_0_reset;
logic [31:0] left_7_0_out;
logic left_7_0_done;
logic [31:0] pe_7_1_top;
logic [31:0] pe_7_1_left;
logic pe_7_1_mul_ready;
logic [31:0] pe_7_1_out;
logic pe_7_1_go;
logic pe_7_1_clk;
logic pe_7_1_reset;
logic pe_7_1_done;
logic [31:0] top_7_1_in;
logic top_7_1_write_en;
logic top_7_1_clk;
logic top_7_1_reset;
logic [31:0] top_7_1_out;
logic top_7_1_done;
logic [31:0] left_7_1_in;
logic left_7_1_write_en;
logic left_7_1_clk;
logic left_7_1_reset;
logic [31:0] left_7_1_out;
logic left_7_1_done;
logic [31:0] pe_7_2_top;
logic [31:0] pe_7_2_left;
logic pe_7_2_mul_ready;
logic [31:0] pe_7_2_out;
logic pe_7_2_go;
logic pe_7_2_clk;
logic pe_7_2_reset;
logic pe_7_2_done;
logic [31:0] top_7_2_in;
logic top_7_2_write_en;
logic top_7_2_clk;
logic top_7_2_reset;
logic [31:0] top_7_2_out;
logic top_7_2_done;
logic [31:0] left_7_2_in;
logic left_7_2_write_en;
logic left_7_2_clk;
logic left_7_2_reset;
logic [31:0] left_7_2_out;
logic left_7_2_done;
logic [31:0] pe_7_3_top;
logic [31:0] pe_7_3_left;
logic pe_7_3_mul_ready;
logic [31:0] pe_7_3_out;
logic pe_7_3_go;
logic pe_7_3_clk;
logic pe_7_3_reset;
logic pe_7_3_done;
logic [31:0] top_7_3_in;
logic top_7_3_write_en;
logic top_7_3_clk;
logic top_7_3_reset;
logic [31:0] top_7_3_out;
logic top_7_3_done;
logic [31:0] left_7_3_in;
logic left_7_3_write_en;
logic left_7_3_clk;
logic left_7_3_reset;
logic [31:0] left_7_3_out;
logic left_7_3_done;
logic [31:0] pe_7_4_top;
logic [31:0] pe_7_4_left;
logic pe_7_4_mul_ready;
logic [31:0] pe_7_4_out;
logic pe_7_4_go;
logic pe_7_4_clk;
logic pe_7_4_reset;
logic pe_7_4_done;
logic [31:0] top_7_4_in;
logic top_7_4_write_en;
logic top_7_4_clk;
logic top_7_4_reset;
logic [31:0] top_7_4_out;
logic top_7_4_done;
logic [31:0] left_7_4_in;
logic left_7_4_write_en;
logic left_7_4_clk;
logic left_7_4_reset;
logic [31:0] left_7_4_out;
logic left_7_4_done;
logic [31:0] pe_7_5_top;
logic [31:0] pe_7_5_left;
logic pe_7_5_mul_ready;
logic [31:0] pe_7_5_out;
logic pe_7_5_go;
logic pe_7_5_clk;
logic pe_7_5_reset;
logic pe_7_5_done;
logic [31:0] top_7_5_in;
logic top_7_5_write_en;
logic top_7_5_clk;
logic top_7_5_reset;
logic [31:0] top_7_5_out;
logic top_7_5_done;
logic [31:0] left_7_5_in;
logic left_7_5_write_en;
logic left_7_5_clk;
logic left_7_5_reset;
logic [31:0] left_7_5_out;
logic left_7_5_done;
logic [31:0] pe_7_6_top;
logic [31:0] pe_7_6_left;
logic pe_7_6_mul_ready;
logic [31:0] pe_7_6_out;
logic pe_7_6_go;
logic pe_7_6_clk;
logic pe_7_6_reset;
logic pe_7_6_done;
logic [31:0] top_7_6_in;
logic top_7_6_write_en;
logic top_7_6_clk;
logic top_7_6_reset;
logic [31:0] top_7_6_out;
logic top_7_6_done;
logic [31:0] left_7_6_in;
logic left_7_6_write_en;
logic left_7_6_clk;
logic left_7_6_reset;
logic [31:0] left_7_6_out;
logic left_7_6_done;
logic [31:0] pe_7_7_top;
logic [31:0] pe_7_7_left;
logic pe_7_7_mul_ready;
logic [31:0] pe_7_7_out;
logic pe_7_7_go;
logic pe_7_7_clk;
logic pe_7_7_reset;
logic pe_7_7_done;
logic [31:0] top_7_7_in;
logic top_7_7_write_en;
logic top_7_7_clk;
logic top_7_7_reset;
logic [31:0] top_7_7_out;
logic top_7_7_done;
logic [31:0] left_7_7_in;
logic left_7_7_write_en;
logic left_7_7_clk;
logic left_7_7_reset;
logic [31:0] left_7_7_out;
logic left_7_7_done;
logic [3:0] t0_idx_in;
logic t0_idx_write_en;
logic t0_idx_clk;
logic t0_idx_reset;
logic [3:0] t0_idx_out;
logic t0_idx_done;
logic [3:0] t0_add_left;
logic [3:0] t0_add_right;
logic [3:0] t0_add_out;
logic [3:0] t1_idx_in;
logic t1_idx_write_en;
logic t1_idx_clk;
logic t1_idx_reset;
logic [3:0] t1_idx_out;
logic t1_idx_done;
logic [3:0] t1_add_left;
logic [3:0] t1_add_right;
logic [3:0] t1_add_out;
logic [3:0] t2_idx_in;
logic t2_idx_write_en;
logic t2_idx_clk;
logic t2_idx_reset;
logic [3:0] t2_idx_out;
logic t2_idx_done;
logic [3:0] t2_add_left;
logic [3:0] t2_add_right;
logic [3:0] t2_add_out;
logic [3:0] t3_idx_in;
logic t3_idx_write_en;
logic t3_idx_clk;
logic t3_idx_reset;
logic [3:0] t3_idx_out;
logic t3_idx_done;
logic [3:0] t3_add_left;
logic [3:0] t3_add_right;
logic [3:0] t3_add_out;
logic [3:0] t4_idx_in;
logic t4_idx_write_en;
logic t4_idx_clk;
logic t4_idx_reset;
logic [3:0] t4_idx_out;
logic t4_idx_done;
logic [3:0] t4_add_left;
logic [3:0] t4_add_right;
logic [3:0] t4_add_out;
logic [3:0] t5_idx_in;
logic t5_idx_write_en;
logic t5_idx_clk;
logic t5_idx_reset;
logic [3:0] t5_idx_out;
logic t5_idx_done;
logic [3:0] t5_add_left;
logic [3:0] t5_add_right;
logic [3:0] t5_add_out;
logic [3:0] t6_idx_in;
logic t6_idx_write_en;
logic t6_idx_clk;
logic t6_idx_reset;
logic [3:0] t6_idx_out;
logic t6_idx_done;
logic [3:0] t6_add_left;
logic [3:0] t6_add_right;
logic [3:0] t6_add_out;
logic [3:0] t7_idx_in;
logic t7_idx_write_en;
logic t7_idx_clk;
logic t7_idx_reset;
logic [3:0] t7_idx_out;
logic t7_idx_done;
logic [3:0] t7_add_left;
logic [3:0] t7_add_right;
logic [3:0] t7_add_out;
logic [3:0] l0_idx_in;
logic l0_idx_write_en;
logic l0_idx_clk;
logic l0_idx_reset;
logic [3:0] l0_idx_out;
logic l0_idx_done;
logic [3:0] l0_add_left;
logic [3:0] l0_add_right;
logic [3:0] l0_add_out;
logic [3:0] l1_idx_in;
logic l1_idx_write_en;
logic l1_idx_clk;
logic l1_idx_reset;
logic [3:0] l1_idx_out;
logic l1_idx_done;
logic [3:0] l1_add_left;
logic [3:0] l1_add_right;
logic [3:0] l1_add_out;
logic [3:0] l2_idx_in;
logic l2_idx_write_en;
logic l2_idx_clk;
logic l2_idx_reset;
logic [3:0] l2_idx_out;
logic l2_idx_done;
logic [3:0] l2_add_left;
logic [3:0] l2_add_right;
logic [3:0] l2_add_out;
logic [3:0] l3_idx_in;
logic l3_idx_write_en;
logic l3_idx_clk;
logic l3_idx_reset;
logic [3:0] l3_idx_out;
logic l3_idx_done;
logic [3:0] l3_add_left;
logic [3:0] l3_add_right;
logic [3:0] l3_add_out;
logic [3:0] l4_idx_in;
logic l4_idx_write_en;
logic l4_idx_clk;
logic l4_idx_reset;
logic [3:0] l4_idx_out;
logic l4_idx_done;
logic [3:0] l4_add_left;
logic [3:0] l4_add_right;
logic [3:0] l4_add_out;
logic [3:0] l5_idx_in;
logic l5_idx_write_en;
logic l5_idx_clk;
logic l5_idx_reset;
logic [3:0] l5_idx_out;
logic l5_idx_done;
logic [3:0] l5_add_left;
logic [3:0] l5_add_right;
logic [3:0] l5_add_out;
logic [3:0] l6_idx_in;
logic l6_idx_write_en;
logic l6_idx_clk;
logic l6_idx_reset;
logic [3:0] l6_idx_out;
logic l6_idx_done;
logic [3:0] l6_add_left;
logic [3:0] l6_add_right;
logic [3:0] l6_add_out;
logic [3:0] l7_idx_in;
logic l7_idx_write_en;
logic l7_idx_clk;
logic l7_idx_reset;
logic [3:0] l7_idx_out;
logic l7_idx_done;
logic [3:0] l7_add_left;
logic [3:0] l7_add_right;
logic [3:0] l7_add_out;
logic [31:0] idx_in;
logic idx_write_en;
logic idx_clk;
logic idx_reset;
logic [31:0] idx_out;
logic idx_done;
logic [31:0] idx_add_left;
logic [31:0] idx_add_right;
logic [31:0] idx_add_out;
logic [31:0] lt_iter_limit_left;
logic [31:0] lt_iter_limit_right;
logic lt_iter_limit_out;
logic cond_reg_in;
logic cond_reg_write_en;
logic cond_reg_clk;
logic cond_reg_reset;
logic cond_reg_out;
logic cond_reg_done;
logic idx_between_depth_plus_16_depth_plus_17_reg_in;
logic idx_between_depth_plus_16_depth_plus_17_reg_write_en;
logic idx_between_depth_plus_16_depth_plus_17_reg_clk;
logic idx_between_depth_plus_16_depth_plus_17_reg_reset;
logic idx_between_depth_plus_16_depth_plus_17_reg_out;
logic idx_between_depth_plus_16_depth_plus_17_reg_done;
logic [31:0] index_lt_depth_plus_17_left;
logic [31:0] index_lt_depth_plus_17_right;
logic index_lt_depth_plus_17_out;
logic [31:0] index_ge_depth_plus_16_left;
logic [31:0] index_ge_depth_plus_16_right;
logic index_ge_depth_plus_16_out;
logic idx_between_depth_plus_16_depth_plus_17_comb_left;
logic idx_between_depth_plus_16_depth_plus_17_comb_right;
logic idx_between_depth_plus_16_depth_plus_17_comb_out;
logic idx_between_depth_plus_12_depth_plus_13_reg_in;
logic idx_between_depth_plus_12_depth_plus_13_reg_write_en;
logic idx_between_depth_plus_12_depth_plus_13_reg_clk;
logic idx_between_depth_plus_12_depth_plus_13_reg_reset;
logic idx_between_depth_plus_12_depth_plus_13_reg_out;
logic idx_between_depth_plus_12_depth_plus_13_reg_done;
logic [31:0] index_lt_depth_plus_13_left;
logic [31:0] index_lt_depth_plus_13_right;
logic index_lt_depth_plus_13_out;
logic [31:0] index_ge_depth_plus_12_left;
logic [31:0] index_ge_depth_plus_12_right;
logic index_ge_depth_plus_12_out;
logic idx_between_depth_plus_12_depth_plus_13_comb_left;
logic idx_between_depth_plus_12_depth_plus_13_comb_right;
logic idx_between_depth_plus_12_depth_plus_13_comb_out;
logic idx_between_depth_plus_8_depth_plus_9_reg_in;
logic idx_between_depth_plus_8_depth_plus_9_reg_write_en;
logic idx_between_depth_plus_8_depth_plus_9_reg_clk;
logic idx_between_depth_plus_8_depth_plus_9_reg_reset;
logic idx_between_depth_plus_8_depth_plus_9_reg_out;
logic idx_between_depth_plus_8_depth_plus_9_reg_done;
logic [31:0] index_lt_depth_plus_9_left;
logic [31:0] index_lt_depth_plus_9_right;
logic index_lt_depth_plus_9_out;
logic [31:0] index_ge_depth_plus_8_left;
logic [31:0] index_ge_depth_plus_8_right;
logic index_ge_depth_plus_8_out;
logic idx_between_depth_plus_8_depth_plus_9_comb_left;
logic idx_between_depth_plus_8_depth_plus_9_comb_right;
logic idx_between_depth_plus_8_depth_plus_9_comb_out;
logic idx_between_2_min_depth_4_plus_2_reg_in;
logic idx_between_2_min_depth_4_plus_2_reg_write_en;
logic idx_between_2_min_depth_4_plus_2_reg_clk;
logic idx_between_2_min_depth_4_plus_2_reg_reset;
logic idx_between_2_min_depth_4_plus_2_reg_out;
logic idx_between_2_min_depth_4_plus_2_reg_done;
logic [31:0] index_lt_min_depth_4_plus_2_left;
logic [31:0] index_lt_min_depth_4_plus_2_right;
logic index_lt_min_depth_4_plus_2_out;
logic [31:0] index_ge_2_left;
logic [31:0] index_ge_2_right;
logic index_ge_2_out;
logic idx_between_2_min_depth_4_plus_2_comb_left;
logic idx_between_2_min_depth_4_plus_2_comb_right;
logic idx_between_2_min_depth_4_plus_2_comb_out;
logic idx_between_2_depth_plus_2_reg_in;
logic idx_between_2_depth_plus_2_reg_write_en;
logic idx_between_2_depth_plus_2_reg_clk;
logic idx_between_2_depth_plus_2_reg_reset;
logic idx_between_2_depth_plus_2_reg_out;
logic idx_between_2_depth_plus_2_reg_done;
logic [31:0] index_lt_depth_plus_2_left;
logic [31:0] index_lt_depth_plus_2_right;
logic index_lt_depth_plus_2_out;
logic idx_between_2_depth_plus_2_comb_left;
logic idx_between_2_depth_plus_2_comb_right;
logic idx_between_2_depth_plus_2_comb_out;
logic idx_between_depth_plus_17_depth_plus_18_reg_in;
logic idx_between_depth_plus_17_depth_plus_18_reg_write_en;
logic idx_between_depth_plus_17_depth_plus_18_reg_clk;
logic idx_between_depth_plus_17_depth_plus_18_reg_reset;
logic idx_between_depth_plus_17_depth_plus_18_reg_out;
logic idx_between_depth_plus_17_depth_plus_18_reg_done;
logic [31:0] index_lt_depth_plus_18_left;
logic [31:0] index_lt_depth_plus_18_right;
logic index_lt_depth_plus_18_out;
logic [31:0] index_ge_depth_plus_17_left;
logic [31:0] index_ge_depth_plus_17_right;
logic index_ge_depth_plus_17_out;
logic idx_between_depth_plus_17_depth_plus_18_comb_left;
logic idx_between_depth_plus_17_depth_plus_18_comb_right;
logic idx_between_depth_plus_17_depth_plus_18_comb_out;
logic idx_between_11_depth_plus_11_reg_in;
logic idx_between_11_depth_plus_11_reg_write_en;
logic idx_between_11_depth_plus_11_reg_clk;
logic idx_between_11_depth_plus_11_reg_reset;
logic idx_between_11_depth_plus_11_reg_out;
logic idx_between_11_depth_plus_11_reg_done;
logic [31:0] index_lt_depth_plus_11_left;
logic [31:0] index_lt_depth_plus_11_right;
logic index_lt_depth_plus_11_out;
logic [31:0] index_ge_11_left;
logic [31:0] index_ge_11_right;
logic index_ge_11_out;
logic idx_between_11_depth_plus_11_comb_left;
logic idx_between_11_depth_plus_11_comb_right;
logic idx_between_11_depth_plus_11_comb_out;
logic idx_between_11_min_depth_4_plus_11_reg_in;
logic idx_between_11_min_depth_4_plus_11_reg_write_en;
logic idx_between_11_min_depth_4_plus_11_reg_clk;
logic idx_between_11_min_depth_4_plus_11_reg_reset;
logic idx_between_11_min_depth_4_plus_11_reg_out;
logic idx_between_11_min_depth_4_plus_11_reg_done;
logic [31:0] index_lt_min_depth_4_plus_11_left;
logic [31:0] index_lt_min_depth_4_plus_11_right;
logic index_lt_min_depth_4_plus_11_out;
logic idx_between_11_min_depth_4_plus_11_comb_left;
logic idx_between_11_min_depth_4_plus_11_comb_right;
logic idx_between_11_min_depth_4_plus_11_comb_out;
logic idx_between_depth_plus_13_depth_plus_14_reg_in;
logic idx_between_depth_plus_13_depth_plus_14_reg_write_en;
logic idx_between_depth_plus_13_depth_plus_14_reg_clk;
logic idx_between_depth_plus_13_depth_plus_14_reg_reset;
logic idx_between_depth_plus_13_depth_plus_14_reg_out;
logic idx_between_depth_plus_13_depth_plus_14_reg_done;
logic [31:0] index_lt_depth_plus_14_left;
logic [31:0] index_lt_depth_plus_14_right;
logic index_lt_depth_plus_14_out;
logic [31:0] index_ge_depth_plus_13_left;
logic [31:0] index_ge_depth_plus_13_right;
logic index_ge_depth_plus_13_out;
logic idx_between_depth_plus_13_depth_plus_14_comb_left;
logic idx_between_depth_plus_13_depth_plus_14_comb_right;
logic idx_between_depth_plus_13_depth_plus_14_comb_out;
logic idx_between_7_depth_plus_7_reg_in;
logic idx_between_7_depth_plus_7_reg_write_en;
logic idx_between_7_depth_plus_7_reg_clk;
logic idx_between_7_depth_plus_7_reg_reset;
logic idx_between_7_depth_plus_7_reg_out;
logic idx_between_7_depth_plus_7_reg_done;
logic [31:0] index_lt_depth_plus_7_left;
logic [31:0] index_lt_depth_plus_7_right;
logic index_lt_depth_plus_7_out;
logic [31:0] index_ge_7_left;
logic [31:0] index_ge_7_right;
logic index_ge_7_out;
logic idx_between_7_depth_plus_7_comb_left;
logic idx_between_7_depth_plus_7_comb_right;
logic idx_between_7_depth_plus_7_comb_out;
logic idx_between_7_min_depth_4_plus_7_reg_in;
logic idx_between_7_min_depth_4_plus_7_reg_write_en;
logic idx_between_7_min_depth_4_plus_7_reg_clk;
logic idx_between_7_min_depth_4_plus_7_reg_reset;
logic idx_between_7_min_depth_4_plus_7_reg_out;
logic idx_between_7_min_depth_4_plus_7_reg_done;
logic [31:0] index_lt_min_depth_4_plus_7_left;
logic [31:0] index_lt_min_depth_4_plus_7_right;
logic index_lt_min_depth_4_plus_7_out;
logic idx_between_7_min_depth_4_plus_7_comb_left;
logic idx_between_7_min_depth_4_plus_7_comb_right;
logic idx_between_7_min_depth_4_plus_7_comb_out;
logic idx_between_16_depth_plus_16_reg_in;
logic idx_between_16_depth_plus_16_reg_write_en;
logic idx_between_16_depth_plus_16_reg_clk;
logic idx_between_16_depth_plus_16_reg_reset;
logic idx_between_16_depth_plus_16_reg_out;
logic idx_between_16_depth_plus_16_reg_done;
logic [31:0] index_lt_depth_plus_16_left;
logic [31:0] index_lt_depth_plus_16_right;
logic index_lt_depth_plus_16_out;
logic [31:0] index_ge_16_left;
logic [31:0] index_ge_16_right;
logic index_ge_16_out;
logic idx_between_16_depth_plus_16_comb_left;
logic idx_between_16_depth_plus_16_comb_right;
logic idx_between_16_depth_plus_16_comb_out;
logic idx_between_depth_plus_18_depth_plus_19_reg_in;
logic idx_between_depth_plus_18_depth_plus_19_reg_write_en;
logic idx_between_depth_plus_18_depth_plus_19_reg_clk;
logic idx_between_depth_plus_18_depth_plus_19_reg_reset;
logic idx_between_depth_plus_18_depth_plus_19_reg_out;
logic idx_between_depth_plus_18_depth_plus_19_reg_done;
logic [31:0] index_lt_depth_plus_19_left;
logic [31:0] index_lt_depth_plus_19_right;
logic index_lt_depth_plus_19_out;
logic [31:0] index_ge_depth_plus_18_left;
logic [31:0] index_ge_depth_plus_18_right;
logic index_ge_depth_plus_18_out;
logic idx_between_depth_plus_18_depth_plus_19_comb_left;
logic idx_between_depth_plus_18_depth_plus_19_comb_right;
logic idx_between_depth_plus_18_depth_plus_19_comb_out;
logic idx_between_3_depth_plus_3_reg_in;
logic idx_between_3_depth_plus_3_reg_write_en;
logic idx_between_3_depth_plus_3_reg_clk;
logic idx_between_3_depth_plus_3_reg_reset;
logic idx_between_3_depth_plus_3_reg_out;
logic idx_between_3_depth_plus_3_reg_done;
logic [31:0] index_lt_depth_plus_3_left;
logic [31:0] index_lt_depth_plus_3_right;
logic index_lt_depth_plus_3_out;
logic [31:0] index_ge_3_left;
logic [31:0] index_ge_3_right;
logic index_ge_3_out;
logic idx_between_3_depth_plus_3_comb_left;
logic idx_between_3_depth_plus_3_comb_right;
logic idx_between_3_depth_plus_3_comb_out;
logic idx_between_12_depth_plus_12_reg_in;
logic idx_between_12_depth_plus_12_reg_write_en;
logic idx_between_12_depth_plus_12_reg_clk;
logic idx_between_12_depth_plus_12_reg_reset;
logic idx_between_12_depth_plus_12_reg_out;
logic idx_between_12_depth_plus_12_reg_done;
logic [31:0] index_lt_depth_plus_12_left;
logic [31:0] index_lt_depth_plus_12_right;
logic index_lt_depth_plus_12_out;
logic [31:0] index_ge_12_left;
logic [31:0] index_ge_12_right;
logic index_ge_12_out;
logic idx_between_12_depth_plus_12_comb_left;
logic idx_between_12_depth_plus_12_comb_right;
logic idx_between_12_depth_plus_12_comb_out;
logic idx_between_3_min_depth_4_plus_3_reg_in;
logic idx_between_3_min_depth_4_plus_3_reg_write_en;
logic idx_between_3_min_depth_4_plus_3_reg_clk;
logic idx_between_3_min_depth_4_plus_3_reg_reset;
logic idx_between_3_min_depth_4_plus_3_reg_out;
logic idx_between_3_min_depth_4_plus_3_reg_done;
logic [31:0] index_lt_min_depth_4_plus_3_left;
logic [31:0] index_lt_min_depth_4_plus_3_right;
logic index_lt_min_depth_4_plus_3_out;
logic idx_between_3_min_depth_4_plus_3_comb_left;
logic idx_between_3_min_depth_4_plus_3_comb_right;
logic idx_between_3_min_depth_4_plus_3_comb_out;
logic idx_between_12_min_depth_4_plus_12_reg_in;
logic idx_between_12_min_depth_4_plus_12_reg_write_en;
logic idx_between_12_min_depth_4_plus_12_reg_clk;
logic idx_between_12_min_depth_4_plus_12_reg_reset;
logic idx_between_12_min_depth_4_plus_12_reg_out;
logic idx_between_12_min_depth_4_plus_12_reg_done;
logic [31:0] index_lt_min_depth_4_plus_12_left;
logic [31:0] index_lt_min_depth_4_plus_12_right;
logic index_lt_min_depth_4_plus_12_out;
logic idx_between_12_min_depth_4_plus_12_comb_left;
logic idx_between_12_min_depth_4_plus_12_comb_right;
logic idx_between_12_min_depth_4_plus_12_comb_out;
logic idx_between_depth_plus_5_depth_plus_6_reg_in;
logic idx_between_depth_plus_5_depth_plus_6_reg_write_en;
logic idx_between_depth_plus_5_depth_plus_6_reg_clk;
logic idx_between_depth_plus_5_depth_plus_6_reg_reset;
logic idx_between_depth_plus_5_depth_plus_6_reg_out;
logic idx_between_depth_plus_5_depth_plus_6_reg_done;
logic [31:0] index_lt_depth_plus_6_left;
logic [31:0] index_lt_depth_plus_6_right;
logic index_lt_depth_plus_6_out;
logic [31:0] index_ge_depth_plus_5_left;
logic [31:0] index_ge_depth_plus_5_right;
logic index_ge_depth_plus_5_out;
logic idx_between_depth_plus_5_depth_plus_6_comb_left;
logic idx_between_depth_plus_5_depth_plus_6_comb_right;
logic idx_between_depth_plus_5_depth_plus_6_comb_out;
logic idx_between_depth_plus_14_depth_plus_15_reg_in;
logic idx_between_depth_plus_14_depth_plus_15_reg_write_en;
logic idx_between_depth_plus_14_depth_plus_15_reg_clk;
logic idx_between_depth_plus_14_depth_plus_15_reg_reset;
logic idx_between_depth_plus_14_depth_plus_15_reg_out;
logic idx_between_depth_plus_14_depth_plus_15_reg_done;
logic [31:0] index_lt_depth_plus_15_left;
logic [31:0] index_lt_depth_plus_15_right;
logic index_lt_depth_plus_15_out;
logic [31:0] index_ge_depth_plus_14_left;
logic [31:0] index_ge_depth_plus_14_right;
logic index_ge_depth_plus_14_out;
logic idx_between_depth_plus_14_depth_plus_15_comb_left;
logic idx_between_depth_plus_14_depth_plus_15_comb_right;
logic idx_between_depth_plus_14_depth_plus_15_comb_out;
logic idx_between_depth_plus_9_depth_plus_10_reg_in;
logic idx_between_depth_plus_9_depth_plus_10_reg_write_en;
logic idx_between_depth_plus_9_depth_plus_10_reg_clk;
logic idx_between_depth_plus_9_depth_plus_10_reg_reset;
logic idx_between_depth_plus_9_depth_plus_10_reg_out;
logic idx_between_depth_plus_9_depth_plus_10_reg_done;
logic [31:0] index_lt_depth_plus_10_left;
logic [31:0] index_lt_depth_plus_10_right;
logic index_lt_depth_plus_10_out;
logic [31:0] index_ge_depth_plus_9_left;
logic [31:0] index_ge_depth_plus_9_right;
logic index_ge_depth_plus_9_out;
logic idx_between_depth_plus_9_depth_plus_10_comb_left;
logic idx_between_depth_plus_9_depth_plus_10_comb_right;
logic idx_between_depth_plus_9_depth_plus_10_comb_out;
logic idx_between_8_depth_plus_8_reg_in;
logic idx_between_8_depth_plus_8_reg_write_en;
logic idx_between_8_depth_plus_8_reg_clk;
logic idx_between_8_depth_plus_8_reg_reset;
logic idx_between_8_depth_plus_8_reg_out;
logic idx_between_8_depth_plus_8_reg_done;
logic [31:0] index_lt_depth_plus_8_left;
logic [31:0] index_lt_depth_plus_8_right;
logic index_lt_depth_plus_8_out;
logic [31:0] index_ge_8_left;
logic [31:0] index_ge_8_right;
logic index_ge_8_out;
logic idx_between_8_depth_plus_8_comb_left;
logic idx_between_8_depth_plus_8_comb_right;
logic idx_between_8_depth_plus_8_comb_out;
logic idx_between_8_min_depth_4_plus_8_reg_in;
logic idx_between_8_min_depth_4_plus_8_reg_write_en;
logic idx_between_8_min_depth_4_plus_8_reg_clk;
logic idx_between_8_min_depth_4_plus_8_reg_reset;
logic idx_between_8_min_depth_4_plus_8_reg_out;
logic idx_between_8_min_depth_4_plus_8_reg_done;
logic [31:0] index_lt_min_depth_4_plus_8_left;
logic [31:0] index_lt_min_depth_4_plus_8_right;
logic index_lt_min_depth_4_plus_8_out;
logic idx_between_8_min_depth_4_plus_8_comb_left;
logic idx_between_8_min_depth_4_plus_8_comb_right;
logic idx_between_8_min_depth_4_plus_8_comb_out;
logic idx_between_17_depth_plus_17_reg_in;
logic idx_between_17_depth_plus_17_reg_write_en;
logic idx_between_17_depth_plus_17_reg_clk;
logic idx_between_17_depth_plus_17_reg_reset;
logic idx_between_17_depth_plus_17_reg_out;
logic idx_between_17_depth_plus_17_reg_done;
logic [31:0] index_ge_17_left;
logic [31:0] index_ge_17_right;
logic index_ge_17_out;
logic idx_between_17_depth_plus_17_comb_left;
logic idx_between_17_depth_plus_17_comb_right;
logic idx_between_17_depth_plus_17_comb_out;
logic idx_between_depth_plus_10_depth_plus_11_reg_in;
logic idx_between_depth_plus_10_depth_plus_11_reg_write_en;
logic idx_between_depth_plus_10_depth_plus_11_reg_clk;
logic idx_between_depth_plus_10_depth_plus_11_reg_reset;
logic idx_between_depth_plus_10_depth_plus_11_reg_out;
logic idx_between_depth_plus_10_depth_plus_11_reg_done;
logic [31:0] index_ge_depth_plus_10_left;
logic [31:0] index_ge_depth_plus_10_right;
logic index_ge_depth_plus_10_out;
logic idx_between_depth_plus_10_depth_plus_11_comb_left;
logic idx_between_depth_plus_10_depth_plus_11_comb_right;
logic idx_between_depth_plus_10_depth_plus_11_comb_out;
logic idx_between_depth_plus_19_depth_plus_20_reg_in;
logic idx_between_depth_plus_19_depth_plus_20_reg_write_en;
logic idx_between_depth_plus_19_depth_plus_20_reg_clk;
logic idx_between_depth_plus_19_depth_plus_20_reg_reset;
logic idx_between_depth_plus_19_depth_plus_20_reg_out;
logic idx_between_depth_plus_19_depth_plus_20_reg_done;
logic [31:0] index_lt_depth_plus_20_left;
logic [31:0] index_lt_depth_plus_20_right;
logic index_lt_depth_plus_20_out;
logic [31:0] index_ge_depth_plus_19_left;
logic [31:0] index_ge_depth_plus_19_right;
logic index_ge_depth_plus_19_out;
logic idx_between_depth_plus_19_depth_plus_20_comb_left;
logic idx_between_depth_plus_19_depth_plus_20_comb_right;
logic idx_between_depth_plus_19_depth_plus_20_comb_out;
logic idx_between_6_min_depth_4_plus_6_reg_in;
logic idx_between_6_min_depth_4_plus_6_reg_write_en;
logic idx_between_6_min_depth_4_plus_6_reg_clk;
logic idx_between_6_min_depth_4_plus_6_reg_reset;
logic idx_between_6_min_depth_4_plus_6_reg_out;
logic idx_between_6_min_depth_4_plus_6_reg_done;
logic [31:0] index_lt_min_depth_4_plus_6_left;
logic [31:0] index_lt_min_depth_4_plus_6_right;
logic index_lt_min_depth_4_plus_6_out;
logic [31:0] index_ge_6_left;
logic [31:0] index_ge_6_right;
logic index_ge_6_out;
logic idx_between_6_min_depth_4_plus_6_comb_left;
logic idx_between_6_min_depth_4_plus_6_comb_right;
logic idx_between_6_min_depth_4_plus_6_comb_out;
logic idx_between_13_depth_plus_13_reg_in;
logic idx_between_13_depth_plus_13_reg_write_en;
logic idx_between_13_depth_plus_13_reg_clk;
logic idx_between_13_depth_plus_13_reg_reset;
logic idx_between_13_depth_plus_13_reg_out;
logic idx_between_13_depth_plus_13_reg_done;
logic [31:0] index_ge_13_left;
logic [31:0] index_ge_13_right;
logic index_ge_13_out;
logic idx_between_13_depth_plus_13_comb_left;
logic idx_between_13_depth_plus_13_comb_right;
logic idx_between_13_depth_plus_13_comb_out;
logic idx_between_13_min_depth_4_plus_13_reg_in;
logic idx_between_13_min_depth_4_plus_13_reg_write_en;
logic idx_between_13_min_depth_4_plus_13_reg_clk;
logic idx_between_13_min_depth_4_plus_13_reg_reset;
logic idx_between_13_min_depth_4_plus_13_reg_out;
logic idx_between_13_min_depth_4_plus_13_reg_done;
logic [31:0] index_lt_min_depth_4_plus_13_left;
logic [31:0] index_lt_min_depth_4_plus_13_right;
logic index_lt_min_depth_4_plus_13_out;
logic idx_between_13_min_depth_4_plus_13_comb_left;
logic idx_between_13_min_depth_4_plus_13_comb_right;
logic idx_between_13_min_depth_4_plus_13_comb_out;
logic idx_between_depth_plus_6_depth_plus_7_reg_in;
logic idx_between_depth_plus_6_depth_plus_7_reg_write_en;
logic idx_between_depth_plus_6_depth_plus_7_reg_clk;
logic idx_between_depth_plus_6_depth_plus_7_reg_reset;
logic idx_between_depth_plus_6_depth_plus_7_reg_out;
logic idx_between_depth_plus_6_depth_plus_7_reg_done;
logic [31:0] index_ge_depth_plus_6_left;
logic [31:0] index_ge_depth_plus_6_right;
logic index_ge_depth_plus_6_out;
logic idx_between_depth_plus_6_depth_plus_7_comb_left;
logic idx_between_depth_plus_6_depth_plus_7_comb_right;
logic idx_between_depth_plus_6_depth_plus_7_comb_out;
logic idx_between_depth_plus_15_depth_plus_16_reg_in;
logic idx_between_depth_plus_15_depth_plus_16_reg_write_en;
logic idx_between_depth_plus_15_depth_plus_16_reg_clk;
logic idx_between_depth_plus_15_depth_plus_16_reg_reset;
logic idx_between_depth_plus_15_depth_plus_16_reg_out;
logic idx_between_depth_plus_15_depth_plus_16_reg_done;
logic [31:0] index_ge_depth_plus_15_left;
logic [31:0] index_ge_depth_plus_15_right;
logic index_ge_depth_plus_15_out;
logic idx_between_depth_plus_15_depth_plus_16_comb_left;
logic idx_between_depth_plus_15_depth_plus_16_comb_right;
logic idx_between_depth_plus_15_depth_plus_16_comb_out;
logic idx_between_18_depth_plus_18_reg_in;
logic idx_between_18_depth_plus_18_reg_write_en;
logic idx_between_18_depth_plus_18_reg_clk;
logic idx_between_18_depth_plus_18_reg_reset;
logic idx_between_18_depth_plus_18_reg_out;
logic idx_between_18_depth_plus_18_reg_done;
logic [31:0] index_ge_18_left;
logic [31:0] index_ge_18_right;
logic index_ge_18_out;
logic idx_between_18_depth_plus_18_comb_left;
logic idx_between_18_depth_plus_18_comb_right;
logic idx_between_18_depth_plus_18_comb_out;
logic idx_between_15_depth_plus_15_reg_in;
logic idx_between_15_depth_plus_15_reg_write_en;
logic idx_between_15_depth_plus_15_reg_clk;
logic idx_between_15_depth_plus_15_reg_reset;
logic idx_between_15_depth_plus_15_reg_out;
logic idx_between_15_depth_plus_15_reg_done;
logic [31:0] index_ge_15_left;
logic [31:0] index_ge_15_right;
logic index_ge_15_out;
logic idx_between_15_depth_plus_15_comb_left;
logic idx_between_15_depth_plus_15_comb_right;
logic idx_between_15_depth_plus_15_comb_out;
logic idx_between_4_depth_plus_4_reg_in;
logic idx_between_4_depth_plus_4_reg_write_en;
logic idx_between_4_depth_plus_4_reg_clk;
logic idx_between_4_depth_plus_4_reg_reset;
logic idx_between_4_depth_plus_4_reg_out;
logic idx_between_4_depth_plus_4_reg_done;
logic [31:0] index_lt_depth_plus_4_left;
logic [31:0] index_lt_depth_plus_4_right;
logic index_lt_depth_plus_4_out;
logic [31:0] index_ge_4_left;
logic [31:0] index_ge_4_right;
logic index_ge_4_out;
logic idx_between_4_depth_plus_4_comb_left;
logic idx_between_4_depth_plus_4_comb_right;
logic idx_between_4_depth_plus_4_comb_out;
logic idx_between_4_min_depth_4_plus_4_reg_in;
logic idx_between_4_min_depth_4_plus_4_reg_write_en;
logic idx_between_4_min_depth_4_plus_4_reg_clk;
logic idx_between_4_min_depth_4_plus_4_reg_reset;
logic idx_between_4_min_depth_4_plus_4_reg_out;
logic idx_between_4_min_depth_4_plus_4_reg_done;
logic [31:0] index_lt_min_depth_4_plus_4_left;
logic [31:0] index_lt_min_depth_4_plus_4_right;
logic index_lt_min_depth_4_plus_4_out;
logic idx_between_4_min_depth_4_plus_4_comb_left;
logic idx_between_4_min_depth_4_plus_4_comb_right;
logic idx_between_4_min_depth_4_plus_4_comb_out;
logic idx_between_5_depth_plus_5_reg_in;
logic idx_between_5_depth_plus_5_reg_write_en;
logic idx_between_5_depth_plus_5_reg_clk;
logic idx_between_5_depth_plus_5_reg_reset;
logic idx_between_5_depth_plus_5_reg_out;
logic idx_between_5_depth_plus_5_reg_done;
logic [31:0] index_lt_depth_plus_5_left;
logic [31:0] index_lt_depth_plus_5_right;
logic index_lt_depth_plus_5_out;
logic [31:0] index_ge_5_left;
logic [31:0] index_ge_5_right;
logic index_ge_5_out;
logic idx_between_5_depth_plus_5_comb_left;
logic idx_between_5_depth_plus_5_comb_right;
logic idx_between_5_depth_plus_5_comb_out;
logic idx_between_14_depth_plus_14_reg_in;
logic idx_between_14_depth_plus_14_reg_write_en;
logic idx_between_14_depth_plus_14_reg_clk;
logic idx_between_14_depth_plus_14_reg_reset;
logic idx_between_14_depth_plus_14_reg_out;
logic idx_between_14_depth_plus_14_reg_done;
logic [31:0] index_ge_14_left;
logic [31:0] index_ge_14_right;
logic index_ge_14_out;
logic idx_between_14_depth_plus_14_comb_left;
logic idx_between_14_depth_plus_14_comb_right;
logic idx_between_14_depth_plus_14_comb_out;
logic idx_between_5_min_depth_4_plus_5_reg_in;
logic idx_between_5_min_depth_4_plus_5_reg_write_en;
logic idx_between_5_min_depth_4_plus_5_reg_clk;
logic idx_between_5_min_depth_4_plus_5_reg_reset;
logic idx_between_5_min_depth_4_plus_5_reg_out;
logic idx_between_5_min_depth_4_plus_5_reg_done;
logic [31:0] index_lt_min_depth_4_plus_5_left;
logic [31:0] index_lt_min_depth_4_plus_5_right;
logic index_lt_min_depth_4_plus_5_out;
logic idx_between_5_min_depth_4_plus_5_comb_left;
logic idx_between_5_min_depth_4_plus_5_comb_right;
logic idx_between_5_min_depth_4_plus_5_comb_out;
logic idx_between_14_min_depth_4_plus_14_reg_in;
logic idx_between_14_min_depth_4_plus_14_reg_write_en;
logic idx_between_14_min_depth_4_plus_14_reg_clk;
logic idx_between_14_min_depth_4_plus_14_reg_reset;
logic idx_between_14_min_depth_4_plus_14_reg_out;
logic idx_between_14_min_depth_4_plus_14_reg_done;
logic [31:0] index_lt_min_depth_4_plus_14_left;
logic [31:0] index_lt_min_depth_4_plus_14_right;
logic index_lt_min_depth_4_plus_14_out;
logic idx_between_14_min_depth_4_plus_14_comb_left;
logic idx_between_14_min_depth_4_plus_14_comb_right;
logic idx_between_14_min_depth_4_plus_14_comb_out;
logic idx_between_0_depth_plus_0_reg_in;
logic idx_between_0_depth_plus_0_reg_write_en;
logic idx_between_0_depth_plus_0_reg_clk;
logic idx_between_0_depth_plus_0_reg_reset;
logic idx_between_0_depth_plus_0_reg_out;
logic idx_between_0_depth_plus_0_reg_done;
logic [31:0] index_lt_depth_plus_0_left;
logic [31:0] index_lt_depth_plus_0_right;
logic index_lt_depth_plus_0_out;
logic idx_between_9_depth_plus_9_reg_in;
logic idx_between_9_depth_plus_9_reg_write_en;
logic idx_between_9_depth_plus_9_reg_clk;
logic idx_between_9_depth_plus_9_reg_reset;
logic idx_between_9_depth_plus_9_reg_out;
logic idx_between_9_depth_plus_9_reg_done;
logic [31:0] index_ge_9_left;
logic [31:0] index_ge_9_right;
logic index_ge_9_out;
logic idx_between_9_depth_plus_9_comb_left;
logic idx_between_9_depth_plus_9_comb_right;
logic idx_between_9_depth_plus_9_comb_out;
logic idx_between_9_min_depth_4_plus_9_reg_in;
logic idx_between_9_min_depth_4_plus_9_reg_write_en;
logic idx_between_9_min_depth_4_plus_9_reg_clk;
logic idx_between_9_min_depth_4_plus_9_reg_reset;
logic idx_between_9_min_depth_4_plus_9_reg_out;
logic idx_between_9_min_depth_4_plus_9_reg_done;
logic [31:0] index_lt_min_depth_4_plus_9_left;
logic [31:0] index_lt_min_depth_4_plus_9_right;
logic index_lt_min_depth_4_plus_9_out;
logic idx_between_9_min_depth_4_plus_9_comb_left;
logic idx_between_9_min_depth_4_plus_9_comb_right;
logic idx_between_9_min_depth_4_plus_9_comb_out;
logic idx_between_1_depth_plus_1_reg_in;
logic idx_between_1_depth_plus_1_reg_write_en;
logic idx_between_1_depth_plus_1_reg_clk;
logic idx_between_1_depth_plus_1_reg_reset;
logic idx_between_1_depth_plus_1_reg_out;
logic idx_between_1_depth_plus_1_reg_done;
logic [31:0] index_lt_depth_plus_1_left;
logic [31:0] index_lt_depth_plus_1_right;
logic index_lt_depth_plus_1_out;
logic [31:0] index_ge_1_left;
logic [31:0] index_ge_1_right;
logic index_ge_1_out;
logic idx_between_1_depth_plus_1_comb_left;
logic idx_between_1_depth_plus_1_comb_right;
logic idx_between_1_depth_plus_1_comb_out;
logic idx_between_1_min_depth_4_plus_1_reg_in;
logic idx_between_1_min_depth_4_plus_1_reg_write_en;
logic idx_between_1_min_depth_4_plus_1_reg_clk;
logic idx_between_1_min_depth_4_plus_1_reg_reset;
logic idx_between_1_min_depth_4_plus_1_reg_out;
logic idx_between_1_min_depth_4_plus_1_reg_done;
logic [31:0] index_lt_min_depth_4_plus_1_left;
logic [31:0] index_lt_min_depth_4_plus_1_right;
logic index_lt_min_depth_4_plus_1_out;
logic idx_between_1_min_depth_4_plus_1_comb_left;
logic idx_between_1_min_depth_4_plus_1_comb_right;
logic idx_between_1_min_depth_4_plus_1_comb_out;
logic idx_between_depth_plus_11_depth_plus_12_reg_in;
logic idx_between_depth_plus_11_depth_plus_12_reg_write_en;
logic idx_between_depth_plus_11_depth_plus_12_reg_clk;
logic idx_between_depth_plus_11_depth_plus_12_reg_reset;
logic idx_between_depth_plus_11_depth_plus_12_reg_out;
logic idx_between_depth_plus_11_depth_plus_12_reg_done;
logic [31:0] index_ge_depth_plus_11_left;
logic [31:0] index_ge_depth_plus_11_right;
logic index_ge_depth_plus_11_out;
logic idx_between_depth_plus_11_depth_plus_12_comb_left;
logic idx_between_depth_plus_11_depth_plus_12_comb_right;
logic idx_between_depth_plus_11_depth_plus_12_comb_out;
logic idx_between_10_depth_plus_10_reg_in;
logic idx_between_10_depth_plus_10_reg_write_en;
logic idx_between_10_depth_plus_10_reg_clk;
logic idx_between_10_depth_plus_10_reg_reset;
logic idx_between_10_depth_plus_10_reg_out;
logic idx_between_10_depth_plus_10_reg_done;
logic [31:0] index_ge_10_left;
logic [31:0] index_ge_10_right;
logic index_ge_10_out;
logic idx_between_10_depth_plus_10_comb_left;
logic idx_between_10_depth_plus_10_comb_right;
logic idx_between_10_depth_plus_10_comb_out;
logic idx_between_10_min_depth_4_plus_10_reg_in;
logic idx_between_10_min_depth_4_plus_10_reg_write_en;
logic idx_between_10_min_depth_4_plus_10_reg_clk;
logic idx_between_10_min_depth_4_plus_10_reg_reset;
logic idx_between_10_min_depth_4_plus_10_reg_out;
logic idx_between_10_min_depth_4_plus_10_reg_done;
logic [31:0] index_lt_min_depth_4_plus_10_left;
logic [31:0] index_lt_min_depth_4_plus_10_right;
logic index_lt_min_depth_4_plus_10_out;
logic idx_between_10_min_depth_4_plus_10_comb_left;
logic idx_between_10_min_depth_4_plus_10_comb_right;
logic idx_between_10_min_depth_4_plus_10_comb_out;
logic idx_between_19_depth_plus_19_reg_in;
logic idx_between_19_depth_plus_19_reg_write_en;
logic idx_between_19_depth_plus_19_reg_clk;
logic idx_between_19_depth_plus_19_reg_reset;
logic idx_between_19_depth_plus_19_reg_out;
logic idx_between_19_depth_plus_19_reg_done;
logic [31:0] index_ge_19_left;
logic [31:0] index_ge_19_right;
logic index_ge_19_out;
logic idx_between_19_depth_plus_19_comb_left;
logic idx_between_19_depth_plus_19_comb_right;
logic idx_between_19_depth_plus_19_comb_out;
logic idx_between_6_depth_plus_6_reg_in;
logic idx_between_6_depth_plus_6_reg_write_en;
logic idx_between_6_depth_plus_6_reg_clk;
logic idx_between_6_depth_plus_6_reg_reset;
logic idx_between_6_depth_plus_6_reg_out;
logic idx_between_6_depth_plus_6_reg_done;
logic idx_between_6_depth_plus_6_comb_left;
logic idx_between_6_depth_plus_6_comb_right;
logic idx_between_6_depth_plus_6_comb_out;
logic idx_between_depth_plus_7_depth_plus_8_reg_in;
logic idx_between_depth_plus_7_depth_plus_8_reg_write_en;
logic idx_between_depth_plus_7_depth_plus_8_reg_clk;
logic idx_between_depth_plus_7_depth_plus_8_reg_reset;
logic idx_between_depth_plus_7_depth_plus_8_reg_out;
logic idx_between_depth_plus_7_depth_plus_8_reg_done;
logic [31:0] index_ge_depth_plus_7_left;
logic [31:0] index_ge_depth_plus_7_right;
logic index_ge_depth_plus_7_out;
logic idx_between_depth_plus_7_depth_plus_8_comb_left;
logic idx_between_depth_plus_7_depth_plus_8_comb_right;
logic idx_between_depth_plus_7_depth_plus_8_comb_out;
logic idx_between_15_min_depth_4_plus_15_reg_in;
logic idx_between_15_min_depth_4_plus_15_reg_write_en;
logic idx_between_15_min_depth_4_plus_15_reg_clk;
logic idx_between_15_min_depth_4_plus_15_reg_reset;
logic idx_between_15_min_depth_4_plus_15_reg_out;
logic idx_between_15_min_depth_4_plus_15_reg_done;
logic [31:0] index_lt_min_depth_4_plus_15_left;
logic [31:0] index_lt_min_depth_4_plus_15_right;
logic index_lt_min_depth_4_plus_15_out;
logic idx_between_15_min_depth_4_plus_15_comb_left;
logic idx_between_15_min_depth_4_plus_15_comb_right;
logic idx_between_15_min_depth_4_plus_15_comb_out;
logic cond_in;
logic cond_write_en;
logic cond_clk;
logic cond_reset;
logic cond_out;
logic cond_done;
logic cond_wire_in;
logic cond_wire_out;
logic cond0_in;
logic cond0_write_en;
logic cond0_clk;
logic cond0_reset;
logic cond0_out;
logic cond0_done;
logic cond_wire0_in;
logic cond_wire0_out;
logic cond1_in;
logic cond1_write_en;
logic cond1_clk;
logic cond1_reset;
logic cond1_out;
logic cond1_done;
logic cond_wire1_in;
logic cond_wire1_out;
logic cond2_in;
logic cond2_write_en;
logic cond2_clk;
logic cond2_reset;
logic cond2_out;
logic cond2_done;
logic cond_wire2_in;
logic cond_wire2_out;
logic cond3_in;
logic cond3_write_en;
logic cond3_clk;
logic cond3_reset;
logic cond3_out;
logic cond3_done;
logic cond_wire3_in;
logic cond_wire3_out;
logic cond4_in;
logic cond4_write_en;
logic cond4_clk;
logic cond4_reset;
logic cond4_out;
logic cond4_done;
logic cond_wire4_in;
logic cond_wire4_out;
logic cond5_in;
logic cond5_write_en;
logic cond5_clk;
logic cond5_reset;
logic cond5_out;
logic cond5_done;
logic cond_wire5_in;
logic cond_wire5_out;
logic cond6_in;
logic cond6_write_en;
logic cond6_clk;
logic cond6_reset;
logic cond6_out;
logic cond6_done;
logic cond_wire6_in;
logic cond_wire6_out;
logic cond7_in;
logic cond7_write_en;
logic cond7_clk;
logic cond7_reset;
logic cond7_out;
logic cond7_done;
logic cond_wire7_in;
logic cond_wire7_out;
logic cond8_in;
logic cond8_write_en;
logic cond8_clk;
logic cond8_reset;
logic cond8_out;
logic cond8_done;
logic cond_wire8_in;
logic cond_wire8_out;
logic cond9_in;
logic cond9_write_en;
logic cond9_clk;
logic cond9_reset;
logic cond9_out;
logic cond9_done;
logic cond_wire9_in;
logic cond_wire9_out;
logic cond10_in;
logic cond10_write_en;
logic cond10_clk;
logic cond10_reset;
logic cond10_out;
logic cond10_done;
logic cond_wire10_in;
logic cond_wire10_out;
logic cond11_in;
logic cond11_write_en;
logic cond11_clk;
logic cond11_reset;
logic cond11_out;
logic cond11_done;
logic cond_wire11_in;
logic cond_wire11_out;
logic cond12_in;
logic cond12_write_en;
logic cond12_clk;
logic cond12_reset;
logic cond12_out;
logic cond12_done;
logic cond_wire12_in;
logic cond_wire12_out;
logic cond13_in;
logic cond13_write_en;
logic cond13_clk;
logic cond13_reset;
logic cond13_out;
logic cond13_done;
logic cond_wire13_in;
logic cond_wire13_out;
logic cond14_in;
logic cond14_write_en;
logic cond14_clk;
logic cond14_reset;
logic cond14_out;
logic cond14_done;
logic cond_wire14_in;
logic cond_wire14_out;
logic cond15_in;
logic cond15_write_en;
logic cond15_clk;
logic cond15_reset;
logic cond15_out;
logic cond15_done;
logic cond_wire15_in;
logic cond_wire15_out;
logic cond16_in;
logic cond16_write_en;
logic cond16_clk;
logic cond16_reset;
logic cond16_out;
logic cond16_done;
logic cond_wire16_in;
logic cond_wire16_out;
logic cond17_in;
logic cond17_write_en;
logic cond17_clk;
logic cond17_reset;
logic cond17_out;
logic cond17_done;
logic cond_wire17_in;
logic cond_wire17_out;
logic cond18_in;
logic cond18_write_en;
logic cond18_clk;
logic cond18_reset;
logic cond18_out;
logic cond18_done;
logic cond_wire18_in;
logic cond_wire18_out;
logic cond19_in;
logic cond19_write_en;
logic cond19_clk;
logic cond19_reset;
logic cond19_out;
logic cond19_done;
logic cond_wire19_in;
logic cond_wire19_out;
logic cond20_in;
logic cond20_write_en;
logic cond20_clk;
logic cond20_reset;
logic cond20_out;
logic cond20_done;
logic cond_wire20_in;
logic cond_wire20_out;
logic cond21_in;
logic cond21_write_en;
logic cond21_clk;
logic cond21_reset;
logic cond21_out;
logic cond21_done;
logic cond_wire21_in;
logic cond_wire21_out;
logic cond22_in;
logic cond22_write_en;
logic cond22_clk;
logic cond22_reset;
logic cond22_out;
logic cond22_done;
logic cond_wire22_in;
logic cond_wire22_out;
logic cond23_in;
logic cond23_write_en;
logic cond23_clk;
logic cond23_reset;
logic cond23_out;
logic cond23_done;
logic cond_wire23_in;
logic cond_wire23_out;
logic cond24_in;
logic cond24_write_en;
logic cond24_clk;
logic cond24_reset;
logic cond24_out;
logic cond24_done;
logic cond_wire24_in;
logic cond_wire24_out;
logic cond25_in;
logic cond25_write_en;
logic cond25_clk;
logic cond25_reset;
logic cond25_out;
logic cond25_done;
logic cond_wire25_in;
logic cond_wire25_out;
logic cond26_in;
logic cond26_write_en;
logic cond26_clk;
logic cond26_reset;
logic cond26_out;
logic cond26_done;
logic cond_wire26_in;
logic cond_wire26_out;
logic cond27_in;
logic cond27_write_en;
logic cond27_clk;
logic cond27_reset;
logic cond27_out;
logic cond27_done;
logic cond_wire27_in;
logic cond_wire27_out;
logic cond28_in;
logic cond28_write_en;
logic cond28_clk;
logic cond28_reset;
logic cond28_out;
logic cond28_done;
logic cond_wire28_in;
logic cond_wire28_out;
logic cond29_in;
logic cond29_write_en;
logic cond29_clk;
logic cond29_reset;
logic cond29_out;
logic cond29_done;
logic cond_wire29_in;
logic cond_wire29_out;
logic cond30_in;
logic cond30_write_en;
logic cond30_clk;
logic cond30_reset;
logic cond30_out;
logic cond30_done;
logic cond_wire30_in;
logic cond_wire30_out;
logic cond31_in;
logic cond31_write_en;
logic cond31_clk;
logic cond31_reset;
logic cond31_out;
logic cond31_done;
logic cond_wire31_in;
logic cond_wire31_out;
logic cond32_in;
logic cond32_write_en;
logic cond32_clk;
logic cond32_reset;
logic cond32_out;
logic cond32_done;
logic cond_wire32_in;
logic cond_wire32_out;
logic cond33_in;
logic cond33_write_en;
logic cond33_clk;
logic cond33_reset;
logic cond33_out;
logic cond33_done;
logic cond_wire33_in;
logic cond_wire33_out;
logic cond34_in;
logic cond34_write_en;
logic cond34_clk;
logic cond34_reset;
logic cond34_out;
logic cond34_done;
logic cond_wire34_in;
logic cond_wire34_out;
logic cond35_in;
logic cond35_write_en;
logic cond35_clk;
logic cond35_reset;
logic cond35_out;
logic cond35_done;
logic cond_wire35_in;
logic cond_wire35_out;
logic cond36_in;
logic cond36_write_en;
logic cond36_clk;
logic cond36_reset;
logic cond36_out;
logic cond36_done;
logic cond_wire36_in;
logic cond_wire36_out;
logic cond37_in;
logic cond37_write_en;
logic cond37_clk;
logic cond37_reset;
logic cond37_out;
logic cond37_done;
logic cond_wire37_in;
logic cond_wire37_out;
logic cond38_in;
logic cond38_write_en;
logic cond38_clk;
logic cond38_reset;
logic cond38_out;
logic cond38_done;
logic cond_wire38_in;
logic cond_wire38_out;
logic cond39_in;
logic cond39_write_en;
logic cond39_clk;
logic cond39_reset;
logic cond39_out;
logic cond39_done;
logic cond_wire39_in;
logic cond_wire39_out;
logic cond40_in;
logic cond40_write_en;
logic cond40_clk;
logic cond40_reset;
logic cond40_out;
logic cond40_done;
logic cond_wire40_in;
logic cond_wire40_out;
logic cond41_in;
logic cond41_write_en;
logic cond41_clk;
logic cond41_reset;
logic cond41_out;
logic cond41_done;
logic cond_wire41_in;
logic cond_wire41_out;
logic cond42_in;
logic cond42_write_en;
logic cond42_clk;
logic cond42_reset;
logic cond42_out;
logic cond42_done;
logic cond_wire42_in;
logic cond_wire42_out;
logic cond43_in;
logic cond43_write_en;
logic cond43_clk;
logic cond43_reset;
logic cond43_out;
logic cond43_done;
logic cond_wire43_in;
logic cond_wire43_out;
logic cond44_in;
logic cond44_write_en;
logic cond44_clk;
logic cond44_reset;
logic cond44_out;
logic cond44_done;
logic cond_wire44_in;
logic cond_wire44_out;
logic cond45_in;
logic cond45_write_en;
logic cond45_clk;
logic cond45_reset;
logic cond45_out;
logic cond45_done;
logic cond_wire45_in;
logic cond_wire45_out;
logic cond46_in;
logic cond46_write_en;
logic cond46_clk;
logic cond46_reset;
logic cond46_out;
logic cond46_done;
logic cond_wire46_in;
logic cond_wire46_out;
logic cond47_in;
logic cond47_write_en;
logic cond47_clk;
logic cond47_reset;
logic cond47_out;
logic cond47_done;
logic cond_wire47_in;
logic cond_wire47_out;
logic cond48_in;
logic cond48_write_en;
logic cond48_clk;
logic cond48_reset;
logic cond48_out;
logic cond48_done;
logic cond_wire48_in;
logic cond_wire48_out;
logic cond49_in;
logic cond49_write_en;
logic cond49_clk;
logic cond49_reset;
logic cond49_out;
logic cond49_done;
logic cond_wire49_in;
logic cond_wire49_out;
logic cond50_in;
logic cond50_write_en;
logic cond50_clk;
logic cond50_reset;
logic cond50_out;
logic cond50_done;
logic cond_wire50_in;
logic cond_wire50_out;
logic cond51_in;
logic cond51_write_en;
logic cond51_clk;
logic cond51_reset;
logic cond51_out;
logic cond51_done;
logic cond_wire51_in;
logic cond_wire51_out;
logic cond52_in;
logic cond52_write_en;
logic cond52_clk;
logic cond52_reset;
logic cond52_out;
logic cond52_done;
logic cond_wire52_in;
logic cond_wire52_out;
logic cond53_in;
logic cond53_write_en;
logic cond53_clk;
logic cond53_reset;
logic cond53_out;
logic cond53_done;
logic cond_wire53_in;
logic cond_wire53_out;
logic cond54_in;
logic cond54_write_en;
logic cond54_clk;
logic cond54_reset;
logic cond54_out;
logic cond54_done;
logic cond_wire54_in;
logic cond_wire54_out;
logic cond55_in;
logic cond55_write_en;
logic cond55_clk;
logic cond55_reset;
logic cond55_out;
logic cond55_done;
logic cond_wire55_in;
logic cond_wire55_out;
logic cond56_in;
logic cond56_write_en;
logic cond56_clk;
logic cond56_reset;
logic cond56_out;
logic cond56_done;
logic cond_wire56_in;
logic cond_wire56_out;
logic cond57_in;
logic cond57_write_en;
logic cond57_clk;
logic cond57_reset;
logic cond57_out;
logic cond57_done;
logic cond_wire57_in;
logic cond_wire57_out;
logic cond58_in;
logic cond58_write_en;
logic cond58_clk;
logic cond58_reset;
logic cond58_out;
logic cond58_done;
logic cond_wire58_in;
logic cond_wire58_out;
logic cond59_in;
logic cond59_write_en;
logic cond59_clk;
logic cond59_reset;
logic cond59_out;
logic cond59_done;
logic cond_wire59_in;
logic cond_wire59_out;
logic cond60_in;
logic cond60_write_en;
logic cond60_clk;
logic cond60_reset;
logic cond60_out;
logic cond60_done;
logic cond_wire60_in;
logic cond_wire60_out;
logic cond61_in;
logic cond61_write_en;
logic cond61_clk;
logic cond61_reset;
logic cond61_out;
logic cond61_done;
logic cond_wire61_in;
logic cond_wire61_out;
logic cond62_in;
logic cond62_write_en;
logic cond62_clk;
logic cond62_reset;
logic cond62_out;
logic cond62_done;
logic cond_wire62_in;
logic cond_wire62_out;
logic cond63_in;
logic cond63_write_en;
logic cond63_clk;
logic cond63_reset;
logic cond63_out;
logic cond63_done;
logic cond_wire63_in;
logic cond_wire63_out;
logic cond64_in;
logic cond64_write_en;
logic cond64_clk;
logic cond64_reset;
logic cond64_out;
logic cond64_done;
logic cond_wire64_in;
logic cond_wire64_out;
logic cond65_in;
logic cond65_write_en;
logic cond65_clk;
logic cond65_reset;
logic cond65_out;
logic cond65_done;
logic cond_wire65_in;
logic cond_wire65_out;
logic cond66_in;
logic cond66_write_en;
logic cond66_clk;
logic cond66_reset;
logic cond66_out;
logic cond66_done;
logic cond_wire66_in;
logic cond_wire66_out;
logic cond67_in;
logic cond67_write_en;
logic cond67_clk;
logic cond67_reset;
logic cond67_out;
logic cond67_done;
logic cond_wire67_in;
logic cond_wire67_out;
logic cond68_in;
logic cond68_write_en;
logic cond68_clk;
logic cond68_reset;
logic cond68_out;
logic cond68_done;
logic cond_wire68_in;
logic cond_wire68_out;
logic cond69_in;
logic cond69_write_en;
logic cond69_clk;
logic cond69_reset;
logic cond69_out;
logic cond69_done;
logic cond_wire69_in;
logic cond_wire69_out;
logic cond70_in;
logic cond70_write_en;
logic cond70_clk;
logic cond70_reset;
logic cond70_out;
logic cond70_done;
logic cond_wire70_in;
logic cond_wire70_out;
logic cond71_in;
logic cond71_write_en;
logic cond71_clk;
logic cond71_reset;
logic cond71_out;
logic cond71_done;
logic cond_wire71_in;
logic cond_wire71_out;
logic cond72_in;
logic cond72_write_en;
logic cond72_clk;
logic cond72_reset;
logic cond72_out;
logic cond72_done;
logic cond_wire72_in;
logic cond_wire72_out;
logic cond73_in;
logic cond73_write_en;
logic cond73_clk;
logic cond73_reset;
logic cond73_out;
logic cond73_done;
logic cond_wire73_in;
logic cond_wire73_out;
logic cond74_in;
logic cond74_write_en;
logic cond74_clk;
logic cond74_reset;
logic cond74_out;
logic cond74_done;
logic cond_wire74_in;
logic cond_wire74_out;
logic cond75_in;
logic cond75_write_en;
logic cond75_clk;
logic cond75_reset;
logic cond75_out;
logic cond75_done;
logic cond_wire75_in;
logic cond_wire75_out;
logic cond76_in;
logic cond76_write_en;
logic cond76_clk;
logic cond76_reset;
logic cond76_out;
logic cond76_done;
logic cond_wire76_in;
logic cond_wire76_out;
logic cond77_in;
logic cond77_write_en;
logic cond77_clk;
logic cond77_reset;
logic cond77_out;
logic cond77_done;
logic cond_wire77_in;
logic cond_wire77_out;
logic cond78_in;
logic cond78_write_en;
logic cond78_clk;
logic cond78_reset;
logic cond78_out;
logic cond78_done;
logic cond_wire78_in;
logic cond_wire78_out;
logic cond79_in;
logic cond79_write_en;
logic cond79_clk;
logic cond79_reset;
logic cond79_out;
logic cond79_done;
logic cond_wire79_in;
logic cond_wire79_out;
logic cond80_in;
logic cond80_write_en;
logic cond80_clk;
logic cond80_reset;
logic cond80_out;
logic cond80_done;
logic cond_wire80_in;
logic cond_wire80_out;
logic cond81_in;
logic cond81_write_en;
logic cond81_clk;
logic cond81_reset;
logic cond81_out;
logic cond81_done;
logic cond_wire81_in;
logic cond_wire81_out;
logic cond82_in;
logic cond82_write_en;
logic cond82_clk;
logic cond82_reset;
logic cond82_out;
logic cond82_done;
logic cond_wire82_in;
logic cond_wire82_out;
logic cond83_in;
logic cond83_write_en;
logic cond83_clk;
logic cond83_reset;
logic cond83_out;
logic cond83_done;
logic cond_wire83_in;
logic cond_wire83_out;
logic cond84_in;
logic cond84_write_en;
logic cond84_clk;
logic cond84_reset;
logic cond84_out;
logic cond84_done;
logic cond_wire84_in;
logic cond_wire84_out;
logic cond85_in;
logic cond85_write_en;
logic cond85_clk;
logic cond85_reset;
logic cond85_out;
logic cond85_done;
logic cond_wire85_in;
logic cond_wire85_out;
logic cond86_in;
logic cond86_write_en;
logic cond86_clk;
logic cond86_reset;
logic cond86_out;
logic cond86_done;
logic cond_wire86_in;
logic cond_wire86_out;
logic cond87_in;
logic cond87_write_en;
logic cond87_clk;
logic cond87_reset;
logic cond87_out;
logic cond87_done;
logic cond_wire87_in;
logic cond_wire87_out;
logic cond88_in;
logic cond88_write_en;
logic cond88_clk;
logic cond88_reset;
logic cond88_out;
logic cond88_done;
logic cond_wire88_in;
logic cond_wire88_out;
logic cond89_in;
logic cond89_write_en;
logic cond89_clk;
logic cond89_reset;
logic cond89_out;
logic cond89_done;
logic cond_wire89_in;
logic cond_wire89_out;
logic cond90_in;
logic cond90_write_en;
logic cond90_clk;
logic cond90_reset;
logic cond90_out;
logic cond90_done;
logic cond_wire90_in;
logic cond_wire90_out;
logic cond91_in;
logic cond91_write_en;
logic cond91_clk;
logic cond91_reset;
logic cond91_out;
logic cond91_done;
logic cond_wire91_in;
logic cond_wire91_out;
logic cond92_in;
logic cond92_write_en;
logic cond92_clk;
logic cond92_reset;
logic cond92_out;
logic cond92_done;
logic cond_wire92_in;
logic cond_wire92_out;
logic cond93_in;
logic cond93_write_en;
logic cond93_clk;
logic cond93_reset;
logic cond93_out;
logic cond93_done;
logic cond_wire93_in;
logic cond_wire93_out;
logic cond94_in;
logic cond94_write_en;
logic cond94_clk;
logic cond94_reset;
logic cond94_out;
logic cond94_done;
logic cond_wire94_in;
logic cond_wire94_out;
logic cond95_in;
logic cond95_write_en;
logic cond95_clk;
logic cond95_reset;
logic cond95_out;
logic cond95_done;
logic cond_wire95_in;
logic cond_wire95_out;
logic cond96_in;
logic cond96_write_en;
logic cond96_clk;
logic cond96_reset;
logic cond96_out;
logic cond96_done;
logic cond_wire96_in;
logic cond_wire96_out;
logic cond97_in;
logic cond97_write_en;
logic cond97_clk;
logic cond97_reset;
logic cond97_out;
logic cond97_done;
logic cond_wire97_in;
logic cond_wire97_out;
logic cond98_in;
logic cond98_write_en;
logic cond98_clk;
logic cond98_reset;
logic cond98_out;
logic cond98_done;
logic cond_wire98_in;
logic cond_wire98_out;
logic cond99_in;
logic cond99_write_en;
logic cond99_clk;
logic cond99_reset;
logic cond99_out;
logic cond99_done;
logic cond_wire99_in;
logic cond_wire99_out;
logic cond100_in;
logic cond100_write_en;
logic cond100_clk;
logic cond100_reset;
logic cond100_out;
logic cond100_done;
logic cond_wire100_in;
logic cond_wire100_out;
logic cond101_in;
logic cond101_write_en;
logic cond101_clk;
logic cond101_reset;
logic cond101_out;
logic cond101_done;
logic cond_wire101_in;
logic cond_wire101_out;
logic cond102_in;
logic cond102_write_en;
logic cond102_clk;
logic cond102_reset;
logic cond102_out;
logic cond102_done;
logic cond_wire102_in;
logic cond_wire102_out;
logic cond103_in;
logic cond103_write_en;
logic cond103_clk;
logic cond103_reset;
logic cond103_out;
logic cond103_done;
logic cond_wire103_in;
logic cond_wire103_out;
logic cond104_in;
logic cond104_write_en;
logic cond104_clk;
logic cond104_reset;
logic cond104_out;
logic cond104_done;
logic cond_wire104_in;
logic cond_wire104_out;
logic cond105_in;
logic cond105_write_en;
logic cond105_clk;
logic cond105_reset;
logic cond105_out;
logic cond105_done;
logic cond_wire105_in;
logic cond_wire105_out;
logic cond106_in;
logic cond106_write_en;
logic cond106_clk;
logic cond106_reset;
logic cond106_out;
logic cond106_done;
logic cond_wire106_in;
logic cond_wire106_out;
logic cond107_in;
logic cond107_write_en;
logic cond107_clk;
logic cond107_reset;
logic cond107_out;
logic cond107_done;
logic cond_wire107_in;
logic cond_wire107_out;
logic cond108_in;
logic cond108_write_en;
logic cond108_clk;
logic cond108_reset;
logic cond108_out;
logic cond108_done;
logic cond_wire108_in;
logic cond_wire108_out;
logic cond109_in;
logic cond109_write_en;
logic cond109_clk;
logic cond109_reset;
logic cond109_out;
logic cond109_done;
logic cond_wire109_in;
logic cond_wire109_out;
logic cond110_in;
logic cond110_write_en;
logic cond110_clk;
logic cond110_reset;
logic cond110_out;
logic cond110_done;
logic cond_wire110_in;
logic cond_wire110_out;
logic cond111_in;
logic cond111_write_en;
logic cond111_clk;
logic cond111_reset;
logic cond111_out;
logic cond111_done;
logic cond_wire111_in;
logic cond_wire111_out;
logic cond112_in;
logic cond112_write_en;
logic cond112_clk;
logic cond112_reset;
logic cond112_out;
logic cond112_done;
logic cond_wire112_in;
logic cond_wire112_out;
logic cond113_in;
logic cond113_write_en;
logic cond113_clk;
logic cond113_reset;
logic cond113_out;
logic cond113_done;
logic cond_wire113_in;
logic cond_wire113_out;
logic cond114_in;
logic cond114_write_en;
logic cond114_clk;
logic cond114_reset;
logic cond114_out;
logic cond114_done;
logic cond_wire114_in;
logic cond_wire114_out;
logic cond115_in;
logic cond115_write_en;
logic cond115_clk;
logic cond115_reset;
logic cond115_out;
logic cond115_done;
logic cond_wire115_in;
logic cond_wire115_out;
logic cond116_in;
logic cond116_write_en;
logic cond116_clk;
logic cond116_reset;
logic cond116_out;
logic cond116_done;
logic cond_wire116_in;
logic cond_wire116_out;
logic cond117_in;
logic cond117_write_en;
logic cond117_clk;
logic cond117_reset;
logic cond117_out;
logic cond117_done;
logic cond_wire117_in;
logic cond_wire117_out;
logic cond118_in;
logic cond118_write_en;
logic cond118_clk;
logic cond118_reset;
logic cond118_out;
logic cond118_done;
logic cond_wire118_in;
logic cond_wire118_out;
logic cond119_in;
logic cond119_write_en;
logic cond119_clk;
logic cond119_reset;
logic cond119_out;
logic cond119_done;
logic cond_wire119_in;
logic cond_wire119_out;
logic cond120_in;
logic cond120_write_en;
logic cond120_clk;
logic cond120_reset;
logic cond120_out;
logic cond120_done;
logic cond_wire120_in;
logic cond_wire120_out;
logic cond121_in;
logic cond121_write_en;
logic cond121_clk;
logic cond121_reset;
logic cond121_out;
logic cond121_done;
logic cond_wire121_in;
logic cond_wire121_out;
logic cond122_in;
logic cond122_write_en;
logic cond122_clk;
logic cond122_reset;
logic cond122_out;
logic cond122_done;
logic cond_wire122_in;
logic cond_wire122_out;
logic cond123_in;
logic cond123_write_en;
logic cond123_clk;
logic cond123_reset;
logic cond123_out;
logic cond123_done;
logic cond_wire123_in;
logic cond_wire123_out;
logic cond124_in;
logic cond124_write_en;
logic cond124_clk;
logic cond124_reset;
logic cond124_out;
logic cond124_done;
logic cond_wire124_in;
logic cond_wire124_out;
logic cond125_in;
logic cond125_write_en;
logic cond125_clk;
logic cond125_reset;
logic cond125_out;
logic cond125_done;
logic cond_wire125_in;
logic cond_wire125_out;
logic cond126_in;
logic cond126_write_en;
logic cond126_clk;
logic cond126_reset;
logic cond126_out;
logic cond126_done;
logic cond_wire126_in;
logic cond_wire126_out;
logic cond127_in;
logic cond127_write_en;
logic cond127_clk;
logic cond127_reset;
logic cond127_out;
logic cond127_done;
logic cond_wire127_in;
logic cond_wire127_out;
logic cond128_in;
logic cond128_write_en;
logic cond128_clk;
logic cond128_reset;
logic cond128_out;
logic cond128_done;
logic cond_wire128_in;
logic cond_wire128_out;
logic cond129_in;
logic cond129_write_en;
logic cond129_clk;
logic cond129_reset;
logic cond129_out;
logic cond129_done;
logic cond_wire129_in;
logic cond_wire129_out;
logic cond130_in;
logic cond130_write_en;
logic cond130_clk;
logic cond130_reset;
logic cond130_out;
logic cond130_done;
logic cond_wire130_in;
logic cond_wire130_out;
logic cond131_in;
logic cond131_write_en;
logic cond131_clk;
logic cond131_reset;
logic cond131_out;
logic cond131_done;
logic cond_wire131_in;
logic cond_wire131_out;
logic cond132_in;
logic cond132_write_en;
logic cond132_clk;
logic cond132_reset;
logic cond132_out;
logic cond132_done;
logic cond_wire132_in;
logic cond_wire132_out;
logic cond133_in;
logic cond133_write_en;
logic cond133_clk;
logic cond133_reset;
logic cond133_out;
logic cond133_done;
logic cond_wire133_in;
logic cond_wire133_out;
logic cond134_in;
logic cond134_write_en;
logic cond134_clk;
logic cond134_reset;
logic cond134_out;
logic cond134_done;
logic cond_wire134_in;
logic cond_wire134_out;
logic cond135_in;
logic cond135_write_en;
logic cond135_clk;
logic cond135_reset;
logic cond135_out;
logic cond135_done;
logic cond_wire135_in;
logic cond_wire135_out;
logic cond136_in;
logic cond136_write_en;
logic cond136_clk;
logic cond136_reset;
logic cond136_out;
logic cond136_done;
logic cond_wire136_in;
logic cond_wire136_out;
logic cond137_in;
logic cond137_write_en;
logic cond137_clk;
logic cond137_reset;
logic cond137_out;
logic cond137_done;
logic cond_wire137_in;
logic cond_wire137_out;
logic cond138_in;
logic cond138_write_en;
logic cond138_clk;
logic cond138_reset;
logic cond138_out;
logic cond138_done;
logic cond_wire138_in;
logic cond_wire138_out;
logic cond139_in;
logic cond139_write_en;
logic cond139_clk;
logic cond139_reset;
logic cond139_out;
logic cond139_done;
logic cond_wire139_in;
logic cond_wire139_out;
logic cond140_in;
logic cond140_write_en;
logic cond140_clk;
logic cond140_reset;
logic cond140_out;
logic cond140_done;
logic cond_wire140_in;
logic cond_wire140_out;
logic cond141_in;
logic cond141_write_en;
logic cond141_clk;
logic cond141_reset;
logic cond141_out;
logic cond141_done;
logic cond_wire141_in;
logic cond_wire141_out;
logic cond142_in;
logic cond142_write_en;
logic cond142_clk;
logic cond142_reset;
logic cond142_out;
logic cond142_done;
logic cond_wire142_in;
logic cond_wire142_out;
logic cond143_in;
logic cond143_write_en;
logic cond143_clk;
logic cond143_reset;
logic cond143_out;
logic cond143_done;
logic cond_wire143_in;
logic cond_wire143_out;
logic cond144_in;
logic cond144_write_en;
logic cond144_clk;
logic cond144_reset;
logic cond144_out;
logic cond144_done;
logic cond_wire144_in;
logic cond_wire144_out;
logic cond145_in;
logic cond145_write_en;
logic cond145_clk;
logic cond145_reset;
logic cond145_out;
logic cond145_done;
logic cond_wire145_in;
logic cond_wire145_out;
logic cond146_in;
logic cond146_write_en;
logic cond146_clk;
logic cond146_reset;
logic cond146_out;
logic cond146_done;
logic cond_wire146_in;
logic cond_wire146_out;
logic cond147_in;
logic cond147_write_en;
logic cond147_clk;
logic cond147_reset;
logic cond147_out;
logic cond147_done;
logic cond_wire147_in;
logic cond_wire147_out;
logic cond148_in;
logic cond148_write_en;
logic cond148_clk;
logic cond148_reset;
logic cond148_out;
logic cond148_done;
logic cond_wire148_in;
logic cond_wire148_out;
logic cond149_in;
logic cond149_write_en;
logic cond149_clk;
logic cond149_reset;
logic cond149_out;
logic cond149_done;
logic cond_wire149_in;
logic cond_wire149_out;
logic cond150_in;
logic cond150_write_en;
logic cond150_clk;
logic cond150_reset;
logic cond150_out;
logic cond150_done;
logic cond_wire150_in;
logic cond_wire150_out;
logic cond151_in;
logic cond151_write_en;
logic cond151_clk;
logic cond151_reset;
logic cond151_out;
logic cond151_done;
logic cond_wire151_in;
logic cond_wire151_out;
logic cond152_in;
logic cond152_write_en;
logic cond152_clk;
logic cond152_reset;
logic cond152_out;
logic cond152_done;
logic cond_wire152_in;
logic cond_wire152_out;
logic cond153_in;
logic cond153_write_en;
logic cond153_clk;
logic cond153_reset;
logic cond153_out;
logic cond153_done;
logic cond_wire153_in;
logic cond_wire153_out;
logic cond154_in;
logic cond154_write_en;
logic cond154_clk;
logic cond154_reset;
logic cond154_out;
logic cond154_done;
logic cond_wire154_in;
logic cond_wire154_out;
logic cond155_in;
logic cond155_write_en;
logic cond155_clk;
logic cond155_reset;
logic cond155_out;
logic cond155_done;
logic cond_wire155_in;
logic cond_wire155_out;
logic cond156_in;
logic cond156_write_en;
logic cond156_clk;
logic cond156_reset;
logic cond156_out;
logic cond156_done;
logic cond_wire156_in;
logic cond_wire156_out;
logic cond157_in;
logic cond157_write_en;
logic cond157_clk;
logic cond157_reset;
logic cond157_out;
logic cond157_done;
logic cond_wire157_in;
logic cond_wire157_out;
logic cond158_in;
logic cond158_write_en;
logic cond158_clk;
logic cond158_reset;
logic cond158_out;
logic cond158_done;
logic cond_wire158_in;
logic cond_wire158_out;
logic cond159_in;
logic cond159_write_en;
logic cond159_clk;
logic cond159_reset;
logic cond159_out;
logic cond159_done;
logic cond_wire159_in;
logic cond_wire159_out;
logic cond160_in;
logic cond160_write_en;
logic cond160_clk;
logic cond160_reset;
logic cond160_out;
logic cond160_done;
logic cond_wire160_in;
logic cond_wire160_out;
logic cond161_in;
logic cond161_write_en;
logic cond161_clk;
logic cond161_reset;
logic cond161_out;
logic cond161_done;
logic cond_wire161_in;
logic cond_wire161_out;
logic cond162_in;
logic cond162_write_en;
logic cond162_clk;
logic cond162_reset;
logic cond162_out;
logic cond162_done;
logic cond_wire162_in;
logic cond_wire162_out;
logic cond163_in;
logic cond163_write_en;
logic cond163_clk;
logic cond163_reset;
logic cond163_out;
logic cond163_done;
logic cond_wire163_in;
logic cond_wire163_out;
logic cond164_in;
logic cond164_write_en;
logic cond164_clk;
logic cond164_reset;
logic cond164_out;
logic cond164_done;
logic cond_wire164_in;
logic cond_wire164_out;
logic cond165_in;
logic cond165_write_en;
logic cond165_clk;
logic cond165_reset;
logic cond165_out;
logic cond165_done;
logic cond_wire165_in;
logic cond_wire165_out;
logic cond166_in;
logic cond166_write_en;
logic cond166_clk;
logic cond166_reset;
logic cond166_out;
logic cond166_done;
logic cond_wire166_in;
logic cond_wire166_out;
logic cond167_in;
logic cond167_write_en;
logic cond167_clk;
logic cond167_reset;
logic cond167_out;
logic cond167_done;
logic cond_wire167_in;
logic cond_wire167_out;
logic cond168_in;
logic cond168_write_en;
logic cond168_clk;
logic cond168_reset;
logic cond168_out;
logic cond168_done;
logic cond_wire168_in;
logic cond_wire168_out;
logic cond169_in;
logic cond169_write_en;
logic cond169_clk;
logic cond169_reset;
logic cond169_out;
logic cond169_done;
logic cond_wire169_in;
logic cond_wire169_out;
logic cond170_in;
logic cond170_write_en;
logic cond170_clk;
logic cond170_reset;
logic cond170_out;
logic cond170_done;
logic cond_wire170_in;
logic cond_wire170_out;
logic cond171_in;
logic cond171_write_en;
logic cond171_clk;
logic cond171_reset;
logic cond171_out;
logic cond171_done;
logic cond_wire171_in;
logic cond_wire171_out;
logic cond172_in;
logic cond172_write_en;
logic cond172_clk;
logic cond172_reset;
logic cond172_out;
logic cond172_done;
logic cond_wire172_in;
logic cond_wire172_out;
logic cond173_in;
logic cond173_write_en;
logic cond173_clk;
logic cond173_reset;
logic cond173_out;
logic cond173_done;
logic cond_wire173_in;
logic cond_wire173_out;
logic cond174_in;
logic cond174_write_en;
logic cond174_clk;
logic cond174_reset;
logic cond174_out;
logic cond174_done;
logic cond_wire174_in;
logic cond_wire174_out;
logic cond175_in;
logic cond175_write_en;
logic cond175_clk;
logic cond175_reset;
logic cond175_out;
logic cond175_done;
logic cond_wire175_in;
logic cond_wire175_out;
logic cond176_in;
logic cond176_write_en;
logic cond176_clk;
logic cond176_reset;
logic cond176_out;
logic cond176_done;
logic cond_wire176_in;
logic cond_wire176_out;
logic cond177_in;
logic cond177_write_en;
logic cond177_clk;
logic cond177_reset;
logic cond177_out;
logic cond177_done;
logic cond_wire177_in;
logic cond_wire177_out;
logic cond178_in;
logic cond178_write_en;
logic cond178_clk;
logic cond178_reset;
logic cond178_out;
logic cond178_done;
logic cond_wire178_in;
logic cond_wire178_out;
logic cond179_in;
logic cond179_write_en;
logic cond179_clk;
logic cond179_reset;
logic cond179_out;
logic cond179_done;
logic cond_wire179_in;
logic cond_wire179_out;
logic cond180_in;
logic cond180_write_en;
logic cond180_clk;
logic cond180_reset;
logic cond180_out;
logic cond180_done;
logic cond_wire180_in;
logic cond_wire180_out;
logic cond181_in;
logic cond181_write_en;
logic cond181_clk;
logic cond181_reset;
logic cond181_out;
logic cond181_done;
logic cond_wire181_in;
logic cond_wire181_out;
logic cond182_in;
logic cond182_write_en;
logic cond182_clk;
logic cond182_reset;
logic cond182_out;
logic cond182_done;
logic cond_wire182_in;
logic cond_wire182_out;
logic cond183_in;
logic cond183_write_en;
logic cond183_clk;
logic cond183_reset;
logic cond183_out;
logic cond183_done;
logic cond_wire183_in;
logic cond_wire183_out;
logic cond184_in;
logic cond184_write_en;
logic cond184_clk;
logic cond184_reset;
logic cond184_out;
logic cond184_done;
logic cond_wire184_in;
logic cond_wire184_out;
logic cond185_in;
logic cond185_write_en;
logic cond185_clk;
logic cond185_reset;
logic cond185_out;
logic cond185_done;
logic cond_wire185_in;
logic cond_wire185_out;
logic cond186_in;
logic cond186_write_en;
logic cond186_clk;
logic cond186_reset;
logic cond186_out;
logic cond186_done;
logic cond_wire186_in;
logic cond_wire186_out;
logic cond187_in;
logic cond187_write_en;
logic cond187_clk;
logic cond187_reset;
logic cond187_out;
logic cond187_done;
logic cond_wire187_in;
logic cond_wire187_out;
logic cond188_in;
logic cond188_write_en;
logic cond188_clk;
logic cond188_reset;
logic cond188_out;
logic cond188_done;
logic cond_wire188_in;
logic cond_wire188_out;
logic cond189_in;
logic cond189_write_en;
logic cond189_clk;
logic cond189_reset;
logic cond189_out;
logic cond189_done;
logic cond_wire189_in;
logic cond_wire189_out;
logic cond190_in;
logic cond190_write_en;
logic cond190_clk;
logic cond190_reset;
logic cond190_out;
logic cond190_done;
logic cond_wire190_in;
logic cond_wire190_out;
logic cond191_in;
logic cond191_write_en;
logic cond191_clk;
logic cond191_reset;
logic cond191_out;
logic cond191_done;
logic cond_wire191_in;
logic cond_wire191_out;
logic cond192_in;
logic cond192_write_en;
logic cond192_clk;
logic cond192_reset;
logic cond192_out;
logic cond192_done;
logic cond_wire192_in;
logic cond_wire192_out;
logic cond193_in;
logic cond193_write_en;
logic cond193_clk;
logic cond193_reset;
logic cond193_out;
logic cond193_done;
logic cond_wire193_in;
logic cond_wire193_out;
logic cond194_in;
logic cond194_write_en;
logic cond194_clk;
logic cond194_reset;
logic cond194_out;
logic cond194_done;
logic cond_wire194_in;
logic cond_wire194_out;
logic cond195_in;
logic cond195_write_en;
logic cond195_clk;
logic cond195_reset;
logic cond195_out;
logic cond195_done;
logic cond_wire195_in;
logic cond_wire195_out;
logic cond196_in;
logic cond196_write_en;
logic cond196_clk;
logic cond196_reset;
logic cond196_out;
logic cond196_done;
logic cond_wire196_in;
logic cond_wire196_out;
logic cond197_in;
logic cond197_write_en;
logic cond197_clk;
logic cond197_reset;
logic cond197_out;
logic cond197_done;
logic cond_wire197_in;
logic cond_wire197_out;
logic cond198_in;
logic cond198_write_en;
logic cond198_clk;
logic cond198_reset;
logic cond198_out;
logic cond198_done;
logic cond_wire198_in;
logic cond_wire198_out;
logic cond199_in;
logic cond199_write_en;
logic cond199_clk;
logic cond199_reset;
logic cond199_out;
logic cond199_done;
logic cond_wire199_in;
logic cond_wire199_out;
logic cond200_in;
logic cond200_write_en;
logic cond200_clk;
logic cond200_reset;
logic cond200_out;
logic cond200_done;
logic cond_wire200_in;
logic cond_wire200_out;
logic cond201_in;
logic cond201_write_en;
logic cond201_clk;
logic cond201_reset;
logic cond201_out;
logic cond201_done;
logic cond_wire201_in;
logic cond_wire201_out;
logic cond202_in;
logic cond202_write_en;
logic cond202_clk;
logic cond202_reset;
logic cond202_out;
logic cond202_done;
logic cond_wire202_in;
logic cond_wire202_out;
logic cond203_in;
logic cond203_write_en;
logic cond203_clk;
logic cond203_reset;
logic cond203_out;
logic cond203_done;
logic cond_wire203_in;
logic cond_wire203_out;
logic cond204_in;
logic cond204_write_en;
logic cond204_clk;
logic cond204_reset;
logic cond204_out;
logic cond204_done;
logic cond_wire204_in;
logic cond_wire204_out;
logic cond205_in;
logic cond205_write_en;
logic cond205_clk;
logic cond205_reset;
logic cond205_out;
logic cond205_done;
logic cond_wire205_in;
logic cond_wire205_out;
logic cond206_in;
logic cond206_write_en;
logic cond206_clk;
logic cond206_reset;
logic cond206_out;
logic cond206_done;
logic cond_wire206_in;
logic cond_wire206_out;
logic cond207_in;
logic cond207_write_en;
logic cond207_clk;
logic cond207_reset;
logic cond207_out;
logic cond207_done;
logic cond_wire207_in;
logic cond_wire207_out;
logic cond208_in;
logic cond208_write_en;
logic cond208_clk;
logic cond208_reset;
logic cond208_out;
logic cond208_done;
logic cond_wire208_in;
logic cond_wire208_out;
logic cond209_in;
logic cond209_write_en;
logic cond209_clk;
logic cond209_reset;
logic cond209_out;
logic cond209_done;
logic cond_wire209_in;
logic cond_wire209_out;
logic cond210_in;
logic cond210_write_en;
logic cond210_clk;
logic cond210_reset;
logic cond210_out;
logic cond210_done;
logic cond_wire210_in;
logic cond_wire210_out;
logic cond211_in;
logic cond211_write_en;
logic cond211_clk;
logic cond211_reset;
logic cond211_out;
logic cond211_done;
logic cond_wire211_in;
logic cond_wire211_out;
logic cond212_in;
logic cond212_write_en;
logic cond212_clk;
logic cond212_reset;
logic cond212_out;
logic cond212_done;
logic cond_wire212_in;
logic cond_wire212_out;
logic cond213_in;
logic cond213_write_en;
logic cond213_clk;
logic cond213_reset;
logic cond213_out;
logic cond213_done;
logic cond_wire213_in;
logic cond_wire213_out;
logic cond214_in;
logic cond214_write_en;
logic cond214_clk;
logic cond214_reset;
logic cond214_out;
logic cond214_done;
logic cond_wire214_in;
logic cond_wire214_out;
logic cond215_in;
logic cond215_write_en;
logic cond215_clk;
logic cond215_reset;
logic cond215_out;
logic cond215_done;
logic cond_wire215_in;
logic cond_wire215_out;
logic cond216_in;
logic cond216_write_en;
logic cond216_clk;
logic cond216_reset;
logic cond216_out;
logic cond216_done;
logic cond_wire216_in;
logic cond_wire216_out;
logic cond217_in;
logic cond217_write_en;
logic cond217_clk;
logic cond217_reset;
logic cond217_out;
logic cond217_done;
logic cond_wire217_in;
logic cond_wire217_out;
logic cond218_in;
logic cond218_write_en;
logic cond218_clk;
logic cond218_reset;
logic cond218_out;
logic cond218_done;
logic cond_wire218_in;
logic cond_wire218_out;
logic cond219_in;
logic cond219_write_en;
logic cond219_clk;
logic cond219_reset;
logic cond219_out;
logic cond219_done;
logic cond_wire219_in;
logic cond_wire219_out;
logic cond220_in;
logic cond220_write_en;
logic cond220_clk;
logic cond220_reset;
logic cond220_out;
logic cond220_done;
logic cond_wire220_in;
logic cond_wire220_out;
logic cond221_in;
logic cond221_write_en;
logic cond221_clk;
logic cond221_reset;
logic cond221_out;
logic cond221_done;
logic cond_wire221_in;
logic cond_wire221_out;
logic cond222_in;
logic cond222_write_en;
logic cond222_clk;
logic cond222_reset;
logic cond222_out;
logic cond222_done;
logic cond_wire222_in;
logic cond_wire222_out;
logic cond223_in;
logic cond223_write_en;
logic cond223_clk;
logic cond223_reset;
logic cond223_out;
logic cond223_done;
logic cond_wire223_in;
logic cond_wire223_out;
logic cond224_in;
logic cond224_write_en;
logic cond224_clk;
logic cond224_reset;
logic cond224_out;
logic cond224_done;
logic cond_wire224_in;
logic cond_wire224_out;
logic cond225_in;
logic cond225_write_en;
logic cond225_clk;
logic cond225_reset;
logic cond225_out;
logic cond225_done;
logic cond_wire225_in;
logic cond_wire225_out;
logic cond226_in;
logic cond226_write_en;
logic cond226_clk;
logic cond226_reset;
logic cond226_out;
logic cond226_done;
logic cond_wire226_in;
logic cond_wire226_out;
logic cond227_in;
logic cond227_write_en;
logic cond227_clk;
logic cond227_reset;
logic cond227_out;
logic cond227_done;
logic cond_wire227_in;
logic cond_wire227_out;
logic cond228_in;
logic cond228_write_en;
logic cond228_clk;
logic cond228_reset;
logic cond228_out;
logic cond228_done;
logic cond_wire228_in;
logic cond_wire228_out;
logic cond229_in;
logic cond229_write_en;
logic cond229_clk;
logic cond229_reset;
logic cond229_out;
logic cond229_done;
logic cond_wire229_in;
logic cond_wire229_out;
logic cond230_in;
logic cond230_write_en;
logic cond230_clk;
logic cond230_reset;
logic cond230_out;
logic cond230_done;
logic cond_wire230_in;
logic cond_wire230_out;
logic cond231_in;
logic cond231_write_en;
logic cond231_clk;
logic cond231_reset;
logic cond231_out;
logic cond231_done;
logic cond_wire231_in;
logic cond_wire231_out;
logic cond232_in;
logic cond232_write_en;
logic cond232_clk;
logic cond232_reset;
logic cond232_out;
logic cond232_done;
logic cond_wire232_in;
logic cond_wire232_out;
logic cond233_in;
logic cond233_write_en;
logic cond233_clk;
logic cond233_reset;
logic cond233_out;
logic cond233_done;
logic cond_wire233_in;
logic cond_wire233_out;
logic cond234_in;
logic cond234_write_en;
logic cond234_clk;
logic cond234_reset;
logic cond234_out;
logic cond234_done;
logic cond_wire234_in;
logic cond_wire234_out;
logic cond235_in;
logic cond235_write_en;
logic cond235_clk;
logic cond235_reset;
logic cond235_out;
logic cond235_done;
logic cond_wire235_in;
logic cond_wire235_out;
logic cond236_in;
logic cond236_write_en;
logic cond236_clk;
logic cond236_reset;
logic cond236_out;
logic cond236_done;
logic cond_wire236_in;
logic cond_wire236_out;
logic cond237_in;
logic cond237_write_en;
logic cond237_clk;
logic cond237_reset;
logic cond237_out;
logic cond237_done;
logic cond_wire237_in;
logic cond_wire237_out;
logic cond238_in;
logic cond238_write_en;
logic cond238_clk;
logic cond238_reset;
logic cond238_out;
logic cond238_done;
logic cond_wire238_in;
logic cond_wire238_out;
logic cond239_in;
logic cond239_write_en;
logic cond239_clk;
logic cond239_reset;
logic cond239_out;
logic cond239_done;
logic cond_wire239_in;
logic cond_wire239_out;
logic cond240_in;
logic cond240_write_en;
logic cond240_clk;
logic cond240_reset;
logic cond240_out;
logic cond240_done;
logic cond_wire240_in;
logic cond_wire240_out;
logic cond241_in;
logic cond241_write_en;
logic cond241_clk;
logic cond241_reset;
logic cond241_out;
logic cond241_done;
logic cond_wire241_in;
logic cond_wire241_out;
logic cond242_in;
logic cond242_write_en;
logic cond242_clk;
logic cond242_reset;
logic cond242_out;
logic cond242_done;
logic cond_wire242_in;
logic cond_wire242_out;
logic cond243_in;
logic cond243_write_en;
logic cond243_clk;
logic cond243_reset;
logic cond243_out;
logic cond243_done;
logic cond_wire243_in;
logic cond_wire243_out;
logic cond244_in;
logic cond244_write_en;
logic cond244_clk;
logic cond244_reset;
logic cond244_out;
logic cond244_done;
logic cond_wire244_in;
logic cond_wire244_out;
logic cond245_in;
logic cond245_write_en;
logic cond245_clk;
logic cond245_reset;
logic cond245_out;
logic cond245_done;
logic cond_wire245_in;
logic cond_wire245_out;
logic cond246_in;
logic cond246_write_en;
logic cond246_clk;
logic cond246_reset;
logic cond246_out;
logic cond246_done;
logic cond_wire246_in;
logic cond_wire246_out;
logic cond247_in;
logic cond247_write_en;
logic cond247_clk;
logic cond247_reset;
logic cond247_out;
logic cond247_done;
logic cond_wire247_in;
logic cond_wire247_out;
logic cond248_in;
logic cond248_write_en;
logic cond248_clk;
logic cond248_reset;
logic cond248_out;
logic cond248_done;
logic cond_wire248_in;
logic cond_wire248_out;
logic cond249_in;
logic cond249_write_en;
logic cond249_clk;
logic cond249_reset;
logic cond249_out;
logic cond249_done;
logic cond_wire249_in;
logic cond_wire249_out;
logic cond250_in;
logic cond250_write_en;
logic cond250_clk;
logic cond250_reset;
logic cond250_out;
logic cond250_done;
logic cond_wire250_in;
logic cond_wire250_out;
logic cond251_in;
logic cond251_write_en;
logic cond251_clk;
logic cond251_reset;
logic cond251_out;
logic cond251_done;
logic cond_wire251_in;
logic cond_wire251_out;
logic cond252_in;
logic cond252_write_en;
logic cond252_clk;
logic cond252_reset;
logic cond252_out;
logic cond252_done;
logic cond_wire252_in;
logic cond_wire252_out;
logic cond253_in;
logic cond253_write_en;
logic cond253_clk;
logic cond253_reset;
logic cond253_out;
logic cond253_done;
logic cond_wire253_in;
logic cond_wire253_out;
logic cond254_in;
logic cond254_write_en;
logic cond254_clk;
logic cond254_reset;
logic cond254_out;
logic cond254_done;
logic cond_wire254_in;
logic cond_wire254_out;
logic cond255_in;
logic cond255_write_en;
logic cond255_clk;
logic cond255_reset;
logic cond255_out;
logic cond255_done;
logic cond_wire255_in;
logic cond_wire255_out;
logic cond256_in;
logic cond256_write_en;
logic cond256_clk;
logic cond256_reset;
logic cond256_out;
logic cond256_done;
logic cond_wire256_in;
logic cond_wire256_out;
logic cond257_in;
logic cond257_write_en;
logic cond257_clk;
logic cond257_reset;
logic cond257_out;
logic cond257_done;
logic cond_wire257_in;
logic cond_wire257_out;
logic cond258_in;
logic cond258_write_en;
logic cond258_clk;
logic cond258_reset;
logic cond258_out;
logic cond258_done;
logic cond_wire258_in;
logic cond_wire258_out;
logic cond259_in;
logic cond259_write_en;
logic cond259_clk;
logic cond259_reset;
logic cond259_out;
logic cond259_done;
logic cond_wire259_in;
logic cond_wire259_out;
logic cond260_in;
logic cond260_write_en;
logic cond260_clk;
logic cond260_reset;
logic cond260_out;
logic cond260_done;
logic cond_wire260_in;
logic cond_wire260_out;
logic cond261_in;
logic cond261_write_en;
logic cond261_clk;
logic cond261_reset;
logic cond261_out;
logic cond261_done;
logic cond_wire261_in;
logic cond_wire261_out;
logic cond262_in;
logic cond262_write_en;
logic cond262_clk;
logic cond262_reset;
logic cond262_out;
logic cond262_done;
logic cond_wire262_in;
logic cond_wire262_out;
logic cond263_in;
logic cond263_write_en;
logic cond263_clk;
logic cond263_reset;
logic cond263_out;
logic cond263_done;
logic cond_wire263_in;
logic cond_wire263_out;
logic cond264_in;
logic cond264_write_en;
logic cond264_clk;
logic cond264_reset;
logic cond264_out;
logic cond264_done;
logic cond_wire264_in;
logic cond_wire264_out;
logic cond265_in;
logic cond265_write_en;
logic cond265_clk;
logic cond265_reset;
logic cond265_out;
logic cond265_done;
logic cond_wire265_in;
logic cond_wire265_out;
logic cond266_in;
logic cond266_write_en;
logic cond266_clk;
logic cond266_reset;
logic cond266_out;
logic cond266_done;
logic cond_wire266_in;
logic cond_wire266_out;
logic cond267_in;
logic cond267_write_en;
logic cond267_clk;
logic cond267_reset;
logic cond267_out;
logic cond267_done;
logic cond_wire267_in;
logic cond_wire267_out;
logic cond268_in;
logic cond268_write_en;
logic cond268_clk;
logic cond268_reset;
logic cond268_out;
logic cond268_done;
logic cond_wire268_in;
logic cond_wire268_out;
logic fsm_in;
logic fsm_write_en;
logic fsm_clk;
logic fsm_reset;
logic fsm_out;
logic fsm_done;
logic ud_out;
logic adder_left;
logic adder_right;
logic adder_out;
logic ud0_out;
logic adder0_left;
logic adder0_right;
logic adder0_out;
logic signal_reg_in;
logic signal_reg_write_en;
logic signal_reg_clk;
logic signal_reg_reset;
logic signal_reg_out;
logic signal_reg_done;
logic [1:0] fsm0_in;
logic fsm0_write_en;
logic fsm0_clk;
logic fsm0_reset;
logic [1:0] fsm0_out;
logic fsm0_done;
logic early_reset_static_par_go_in;
logic early_reset_static_par_go_out;
logic early_reset_static_par_done_in;
logic early_reset_static_par_done_out;
logic early_reset_static_par0_go_in;
logic early_reset_static_par0_go_out;
logic early_reset_static_par0_done_in;
logic early_reset_static_par0_done_out;
logic wrapper_early_reset_static_par_go_in;
logic wrapper_early_reset_static_par_go_out;
logic wrapper_early_reset_static_par_done_in;
logic wrapper_early_reset_static_par_done_out;
logic while_wrapper_early_reset_static_par0_go_in;
logic while_wrapper_early_reset_static_par0_go_out;
logic while_wrapper_early_reset_static_par0_done_in;
logic while_wrapper_early_reset_static_par0_done_out;
logic tdcc_go_in;
logic tdcc_go_out;
logic tdcc_done_in;
logic tdcc_done_out;
std_reg # (
    .WIDTH(32)
) min_depth_4 (
    .clk(min_depth_4_clk),
    .done(min_depth_4_done),
    .in(min_depth_4_in),
    .out(min_depth_4_out),
    .reset(min_depth_4_reset),
    .write_en(min_depth_4_write_en)
);
std_reg # (
    .WIDTH(32)
) iter_limit (
    .clk(iter_limit_clk),
    .done(iter_limit_done),
    .in(iter_limit_in),
    .out(iter_limit_out),
    .reset(iter_limit_reset),
    .write_en(iter_limit_write_en)
);
std_add # (
    .WIDTH(32)
) depth_plus_16 (
    .left(depth_plus_16_left),
    .out(depth_plus_16_out),
    .right(depth_plus_16_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_17 (
    .left(depth_plus_17_left),
    .out(depth_plus_17_out),
    .right(depth_plus_17_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_12 (
    .left(depth_plus_12_left),
    .out(depth_plus_12_out),
    .right(depth_plus_12_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_13 (
    .left(depth_plus_13_left),
    .out(depth_plus_13_out),
    .right(depth_plus_13_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_8 (
    .left(depth_plus_8_left),
    .out(depth_plus_8_out),
    .right(depth_plus_8_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_9 (
    .left(depth_plus_9_left),
    .out(depth_plus_9_out),
    .right(depth_plus_9_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_2 (
    .left(min_depth_4_plus_2_left),
    .out(min_depth_4_plus_2_out),
    .right(min_depth_4_plus_2_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_2 (
    .left(depth_plus_2_left),
    .out(depth_plus_2_out),
    .right(depth_plus_2_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_18 (
    .left(depth_plus_18_left),
    .out(depth_plus_18_out),
    .right(depth_plus_18_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_11 (
    .left(depth_plus_11_left),
    .out(depth_plus_11_out),
    .right(depth_plus_11_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_11 (
    .left(min_depth_4_plus_11_left),
    .out(min_depth_4_plus_11_out),
    .right(min_depth_4_plus_11_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_14 (
    .left(depth_plus_14_left),
    .out(depth_plus_14_out),
    .right(depth_plus_14_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_7 (
    .left(depth_plus_7_left),
    .out(depth_plus_7_out),
    .right(depth_plus_7_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_7 (
    .left(min_depth_4_plus_7_left),
    .out(min_depth_4_plus_7_out),
    .right(min_depth_4_plus_7_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_19 (
    .left(depth_plus_19_left),
    .out(depth_plus_19_out),
    .right(depth_plus_19_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_3 (
    .left(depth_plus_3_left),
    .out(depth_plus_3_out),
    .right(depth_plus_3_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_3 (
    .left(min_depth_4_plus_3_left),
    .out(min_depth_4_plus_3_out),
    .right(min_depth_4_plus_3_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_12 (
    .left(min_depth_4_plus_12_left),
    .out(min_depth_4_plus_12_out),
    .right(min_depth_4_plus_12_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_5 (
    .left(depth_plus_5_left),
    .out(depth_plus_5_out),
    .right(depth_plus_5_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_6 (
    .left(depth_plus_6_left),
    .out(depth_plus_6_out),
    .right(depth_plus_6_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_15 (
    .left(depth_plus_15_left),
    .out(depth_plus_15_out),
    .right(depth_plus_15_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_10 (
    .left(depth_plus_10_left),
    .out(depth_plus_10_out),
    .right(depth_plus_10_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_8 (
    .left(min_depth_4_plus_8_left),
    .out(min_depth_4_plus_8_out),
    .right(min_depth_4_plus_8_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_20 (
    .left(depth_plus_20_left),
    .out(depth_plus_20_out),
    .right(depth_plus_20_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_6 (
    .left(min_depth_4_plus_6_left),
    .out(min_depth_4_plus_6_out),
    .right(min_depth_4_plus_6_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_13 (
    .left(min_depth_4_plus_13_left),
    .out(min_depth_4_plus_13_out),
    .right(min_depth_4_plus_13_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_4 (
    .left(depth_plus_4_left),
    .out(depth_plus_4_out),
    .right(depth_plus_4_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_4 (
    .left(min_depth_4_plus_4_left),
    .out(min_depth_4_plus_4_out),
    .right(min_depth_4_plus_4_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_5 (
    .left(min_depth_4_plus_5_left),
    .out(min_depth_4_plus_5_out),
    .right(min_depth_4_plus_5_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_14 (
    .left(min_depth_4_plus_14_left),
    .out(min_depth_4_plus_14_out),
    .right(min_depth_4_plus_14_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_0 (
    .left(depth_plus_0_left),
    .out(depth_plus_0_out),
    .right(depth_plus_0_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_9 (
    .left(min_depth_4_plus_9_left),
    .out(min_depth_4_plus_9_out),
    .right(min_depth_4_plus_9_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_1 (
    .left(depth_plus_1_left),
    .out(depth_plus_1_out),
    .right(depth_plus_1_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_1 (
    .left(min_depth_4_plus_1_left),
    .out(min_depth_4_plus_1_out),
    .right(min_depth_4_plus_1_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_10 (
    .left(min_depth_4_plus_10_left),
    .out(min_depth_4_plus_10_out),
    .right(min_depth_4_plus_10_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_15 (
    .left(min_depth_4_plus_15_left),
    .out(min_depth_4_plus_15_out),
    .right(min_depth_4_plus_15_right)
);
mac_pe pe_0_0 (
    .clk(pe_0_0_clk),
    .done(pe_0_0_done),
    .go(pe_0_0_go),
    .left(pe_0_0_left),
    .mul_ready(pe_0_0_mul_ready),
    .out(pe_0_0_out),
    .reset(pe_0_0_reset),
    .top(pe_0_0_top)
);
std_reg # (
    .WIDTH(32)
) top_0_0 (
    .clk(top_0_0_clk),
    .done(top_0_0_done),
    .in(top_0_0_in),
    .out(top_0_0_out),
    .reset(top_0_0_reset),
    .write_en(top_0_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_0 (
    .clk(left_0_0_clk),
    .done(left_0_0_done),
    .in(left_0_0_in),
    .out(left_0_0_out),
    .reset(left_0_0_reset),
    .write_en(left_0_0_write_en)
);
mac_pe pe_0_1 (
    .clk(pe_0_1_clk),
    .done(pe_0_1_done),
    .go(pe_0_1_go),
    .left(pe_0_1_left),
    .mul_ready(pe_0_1_mul_ready),
    .out(pe_0_1_out),
    .reset(pe_0_1_reset),
    .top(pe_0_1_top)
);
std_reg # (
    .WIDTH(32)
) top_0_1 (
    .clk(top_0_1_clk),
    .done(top_0_1_done),
    .in(top_0_1_in),
    .out(top_0_1_out),
    .reset(top_0_1_reset),
    .write_en(top_0_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_1 (
    .clk(left_0_1_clk),
    .done(left_0_1_done),
    .in(left_0_1_in),
    .out(left_0_1_out),
    .reset(left_0_1_reset),
    .write_en(left_0_1_write_en)
);
mac_pe pe_0_2 (
    .clk(pe_0_2_clk),
    .done(pe_0_2_done),
    .go(pe_0_2_go),
    .left(pe_0_2_left),
    .mul_ready(pe_0_2_mul_ready),
    .out(pe_0_2_out),
    .reset(pe_0_2_reset),
    .top(pe_0_2_top)
);
std_reg # (
    .WIDTH(32)
) top_0_2 (
    .clk(top_0_2_clk),
    .done(top_0_2_done),
    .in(top_0_2_in),
    .out(top_0_2_out),
    .reset(top_0_2_reset),
    .write_en(top_0_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_2 (
    .clk(left_0_2_clk),
    .done(left_0_2_done),
    .in(left_0_2_in),
    .out(left_0_2_out),
    .reset(left_0_2_reset),
    .write_en(left_0_2_write_en)
);
mac_pe pe_0_3 (
    .clk(pe_0_3_clk),
    .done(pe_0_3_done),
    .go(pe_0_3_go),
    .left(pe_0_3_left),
    .mul_ready(pe_0_3_mul_ready),
    .out(pe_0_3_out),
    .reset(pe_0_3_reset),
    .top(pe_0_3_top)
);
std_reg # (
    .WIDTH(32)
) top_0_3 (
    .clk(top_0_3_clk),
    .done(top_0_3_done),
    .in(top_0_3_in),
    .out(top_0_3_out),
    .reset(top_0_3_reset),
    .write_en(top_0_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_3 (
    .clk(left_0_3_clk),
    .done(left_0_3_done),
    .in(left_0_3_in),
    .out(left_0_3_out),
    .reset(left_0_3_reset),
    .write_en(left_0_3_write_en)
);
mac_pe pe_0_4 (
    .clk(pe_0_4_clk),
    .done(pe_0_4_done),
    .go(pe_0_4_go),
    .left(pe_0_4_left),
    .mul_ready(pe_0_4_mul_ready),
    .out(pe_0_4_out),
    .reset(pe_0_4_reset),
    .top(pe_0_4_top)
);
std_reg # (
    .WIDTH(32)
) top_0_4 (
    .clk(top_0_4_clk),
    .done(top_0_4_done),
    .in(top_0_4_in),
    .out(top_0_4_out),
    .reset(top_0_4_reset),
    .write_en(top_0_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_4 (
    .clk(left_0_4_clk),
    .done(left_0_4_done),
    .in(left_0_4_in),
    .out(left_0_4_out),
    .reset(left_0_4_reset),
    .write_en(left_0_4_write_en)
);
mac_pe pe_0_5 (
    .clk(pe_0_5_clk),
    .done(pe_0_5_done),
    .go(pe_0_5_go),
    .left(pe_0_5_left),
    .mul_ready(pe_0_5_mul_ready),
    .out(pe_0_5_out),
    .reset(pe_0_5_reset),
    .top(pe_0_5_top)
);
std_reg # (
    .WIDTH(32)
) top_0_5 (
    .clk(top_0_5_clk),
    .done(top_0_5_done),
    .in(top_0_5_in),
    .out(top_0_5_out),
    .reset(top_0_5_reset),
    .write_en(top_0_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_5 (
    .clk(left_0_5_clk),
    .done(left_0_5_done),
    .in(left_0_5_in),
    .out(left_0_5_out),
    .reset(left_0_5_reset),
    .write_en(left_0_5_write_en)
);
mac_pe pe_0_6 (
    .clk(pe_0_6_clk),
    .done(pe_0_6_done),
    .go(pe_0_6_go),
    .left(pe_0_6_left),
    .mul_ready(pe_0_6_mul_ready),
    .out(pe_0_6_out),
    .reset(pe_0_6_reset),
    .top(pe_0_6_top)
);
std_reg # (
    .WIDTH(32)
) top_0_6 (
    .clk(top_0_6_clk),
    .done(top_0_6_done),
    .in(top_0_6_in),
    .out(top_0_6_out),
    .reset(top_0_6_reset),
    .write_en(top_0_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_6 (
    .clk(left_0_6_clk),
    .done(left_0_6_done),
    .in(left_0_6_in),
    .out(left_0_6_out),
    .reset(left_0_6_reset),
    .write_en(left_0_6_write_en)
);
mac_pe pe_0_7 (
    .clk(pe_0_7_clk),
    .done(pe_0_7_done),
    .go(pe_0_7_go),
    .left(pe_0_7_left),
    .mul_ready(pe_0_7_mul_ready),
    .out(pe_0_7_out),
    .reset(pe_0_7_reset),
    .top(pe_0_7_top)
);
std_reg # (
    .WIDTH(32)
) top_0_7 (
    .clk(top_0_7_clk),
    .done(top_0_7_done),
    .in(top_0_7_in),
    .out(top_0_7_out),
    .reset(top_0_7_reset),
    .write_en(top_0_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_7 (
    .clk(left_0_7_clk),
    .done(left_0_7_done),
    .in(left_0_7_in),
    .out(left_0_7_out),
    .reset(left_0_7_reset),
    .write_en(left_0_7_write_en)
);
mac_pe pe_1_0 (
    .clk(pe_1_0_clk),
    .done(pe_1_0_done),
    .go(pe_1_0_go),
    .left(pe_1_0_left),
    .mul_ready(pe_1_0_mul_ready),
    .out(pe_1_0_out),
    .reset(pe_1_0_reset),
    .top(pe_1_0_top)
);
std_reg # (
    .WIDTH(32)
) top_1_0 (
    .clk(top_1_0_clk),
    .done(top_1_0_done),
    .in(top_1_0_in),
    .out(top_1_0_out),
    .reset(top_1_0_reset),
    .write_en(top_1_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_0 (
    .clk(left_1_0_clk),
    .done(left_1_0_done),
    .in(left_1_0_in),
    .out(left_1_0_out),
    .reset(left_1_0_reset),
    .write_en(left_1_0_write_en)
);
mac_pe pe_1_1 (
    .clk(pe_1_1_clk),
    .done(pe_1_1_done),
    .go(pe_1_1_go),
    .left(pe_1_1_left),
    .mul_ready(pe_1_1_mul_ready),
    .out(pe_1_1_out),
    .reset(pe_1_1_reset),
    .top(pe_1_1_top)
);
std_reg # (
    .WIDTH(32)
) top_1_1 (
    .clk(top_1_1_clk),
    .done(top_1_1_done),
    .in(top_1_1_in),
    .out(top_1_1_out),
    .reset(top_1_1_reset),
    .write_en(top_1_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_1 (
    .clk(left_1_1_clk),
    .done(left_1_1_done),
    .in(left_1_1_in),
    .out(left_1_1_out),
    .reset(left_1_1_reset),
    .write_en(left_1_1_write_en)
);
mac_pe pe_1_2 (
    .clk(pe_1_2_clk),
    .done(pe_1_2_done),
    .go(pe_1_2_go),
    .left(pe_1_2_left),
    .mul_ready(pe_1_2_mul_ready),
    .out(pe_1_2_out),
    .reset(pe_1_2_reset),
    .top(pe_1_2_top)
);
std_reg # (
    .WIDTH(32)
) top_1_2 (
    .clk(top_1_2_clk),
    .done(top_1_2_done),
    .in(top_1_2_in),
    .out(top_1_2_out),
    .reset(top_1_2_reset),
    .write_en(top_1_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_2 (
    .clk(left_1_2_clk),
    .done(left_1_2_done),
    .in(left_1_2_in),
    .out(left_1_2_out),
    .reset(left_1_2_reset),
    .write_en(left_1_2_write_en)
);
mac_pe pe_1_3 (
    .clk(pe_1_3_clk),
    .done(pe_1_3_done),
    .go(pe_1_3_go),
    .left(pe_1_3_left),
    .mul_ready(pe_1_3_mul_ready),
    .out(pe_1_3_out),
    .reset(pe_1_3_reset),
    .top(pe_1_3_top)
);
std_reg # (
    .WIDTH(32)
) top_1_3 (
    .clk(top_1_3_clk),
    .done(top_1_3_done),
    .in(top_1_3_in),
    .out(top_1_3_out),
    .reset(top_1_3_reset),
    .write_en(top_1_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_3 (
    .clk(left_1_3_clk),
    .done(left_1_3_done),
    .in(left_1_3_in),
    .out(left_1_3_out),
    .reset(left_1_3_reset),
    .write_en(left_1_3_write_en)
);
mac_pe pe_1_4 (
    .clk(pe_1_4_clk),
    .done(pe_1_4_done),
    .go(pe_1_4_go),
    .left(pe_1_4_left),
    .mul_ready(pe_1_4_mul_ready),
    .out(pe_1_4_out),
    .reset(pe_1_4_reset),
    .top(pe_1_4_top)
);
std_reg # (
    .WIDTH(32)
) top_1_4 (
    .clk(top_1_4_clk),
    .done(top_1_4_done),
    .in(top_1_4_in),
    .out(top_1_4_out),
    .reset(top_1_4_reset),
    .write_en(top_1_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_4 (
    .clk(left_1_4_clk),
    .done(left_1_4_done),
    .in(left_1_4_in),
    .out(left_1_4_out),
    .reset(left_1_4_reset),
    .write_en(left_1_4_write_en)
);
mac_pe pe_1_5 (
    .clk(pe_1_5_clk),
    .done(pe_1_5_done),
    .go(pe_1_5_go),
    .left(pe_1_5_left),
    .mul_ready(pe_1_5_mul_ready),
    .out(pe_1_5_out),
    .reset(pe_1_5_reset),
    .top(pe_1_5_top)
);
std_reg # (
    .WIDTH(32)
) top_1_5 (
    .clk(top_1_5_clk),
    .done(top_1_5_done),
    .in(top_1_5_in),
    .out(top_1_5_out),
    .reset(top_1_5_reset),
    .write_en(top_1_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_5 (
    .clk(left_1_5_clk),
    .done(left_1_5_done),
    .in(left_1_5_in),
    .out(left_1_5_out),
    .reset(left_1_5_reset),
    .write_en(left_1_5_write_en)
);
mac_pe pe_1_6 (
    .clk(pe_1_6_clk),
    .done(pe_1_6_done),
    .go(pe_1_6_go),
    .left(pe_1_6_left),
    .mul_ready(pe_1_6_mul_ready),
    .out(pe_1_6_out),
    .reset(pe_1_6_reset),
    .top(pe_1_6_top)
);
std_reg # (
    .WIDTH(32)
) top_1_6 (
    .clk(top_1_6_clk),
    .done(top_1_6_done),
    .in(top_1_6_in),
    .out(top_1_6_out),
    .reset(top_1_6_reset),
    .write_en(top_1_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_6 (
    .clk(left_1_6_clk),
    .done(left_1_6_done),
    .in(left_1_6_in),
    .out(left_1_6_out),
    .reset(left_1_6_reset),
    .write_en(left_1_6_write_en)
);
mac_pe pe_1_7 (
    .clk(pe_1_7_clk),
    .done(pe_1_7_done),
    .go(pe_1_7_go),
    .left(pe_1_7_left),
    .mul_ready(pe_1_7_mul_ready),
    .out(pe_1_7_out),
    .reset(pe_1_7_reset),
    .top(pe_1_7_top)
);
std_reg # (
    .WIDTH(32)
) top_1_7 (
    .clk(top_1_7_clk),
    .done(top_1_7_done),
    .in(top_1_7_in),
    .out(top_1_7_out),
    .reset(top_1_7_reset),
    .write_en(top_1_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_7 (
    .clk(left_1_7_clk),
    .done(left_1_7_done),
    .in(left_1_7_in),
    .out(left_1_7_out),
    .reset(left_1_7_reset),
    .write_en(left_1_7_write_en)
);
mac_pe pe_2_0 (
    .clk(pe_2_0_clk),
    .done(pe_2_0_done),
    .go(pe_2_0_go),
    .left(pe_2_0_left),
    .mul_ready(pe_2_0_mul_ready),
    .out(pe_2_0_out),
    .reset(pe_2_0_reset),
    .top(pe_2_0_top)
);
std_reg # (
    .WIDTH(32)
) top_2_0 (
    .clk(top_2_0_clk),
    .done(top_2_0_done),
    .in(top_2_0_in),
    .out(top_2_0_out),
    .reset(top_2_0_reset),
    .write_en(top_2_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_0 (
    .clk(left_2_0_clk),
    .done(left_2_0_done),
    .in(left_2_0_in),
    .out(left_2_0_out),
    .reset(left_2_0_reset),
    .write_en(left_2_0_write_en)
);
mac_pe pe_2_1 (
    .clk(pe_2_1_clk),
    .done(pe_2_1_done),
    .go(pe_2_1_go),
    .left(pe_2_1_left),
    .mul_ready(pe_2_1_mul_ready),
    .out(pe_2_1_out),
    .reset(pe_2_1_reset),
    .top(pe_2_1_top)
);
std_reg # (
    .WIDTH(32)
) top_2_1 (
    .clk(top_2_1_clk),
    .done(top_2_1_done),
    .in(top_2_1_in),
    .out(top_2_1_out),
    .reset(top_2_1_reset),
    .write_en(top_2_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_1 (
    .clk(left_2_1_clk),
    .done(left_2_1_done),
    .in(left_2_1_in),
    .out(left_2_1_out),
    .reset(left_2_1_reset),
    .write_en(left_2_1_write_en)
);
mac_pe pe_2_2 (
    .clk(pe_2_2_clk),
    .done(pe_2_2_done),
    .go(pe_2_2_go),
    .left(pe_2_2_left),
    .mul_ready(pe_2_2_mul_ready),
    .out(pe_2_2_out),
    .reset(pe_2_2_reset),
    .top(pe_2_2_top)
);
std_reg # (
    .WIDTH(32)
) top_2_2 (
    .clk(top_2_2_clk),
    .done(top_2_2_done),
    .in(top_2_2_in),
    .out(top_2_2_out),
    .reset(top_2_2_reset),
    .write_en(top_2_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_2 (
    .clk(left_2_2_clk),
    .done(left_2_2_done),
    .in(left_2_2_in),
    .out(left_2_2_out),
    .reset(left_2_2_reset),
    .write_en(left_2_2_write_en)
);
mac_pe pe_2_3 (
    .clk(pe_2_3_clk),
    .done(pe_2_3_done),
    .go(pe_2_3_go),
    .left(pe_2_3_left),
    .mul_ready(pe_2_3_mul_ready),
    .out(pe_2_3_out),
    .reset(pe_2_3_reset),
    .top(pe_2_3_top)
);
std_reg # (
    .WIDTH(32)
) top_2_3 (
    .clk(top_2_3_clk),
    .done(top_2_3_done),
    .in(top_2_3_in),
    .out(top_2_3_out),
    .reset(top_2_3_reset),
    .write_en(top_2_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_3 (
    .clk(left_2_3_clk),
    .done(left_2_3_done),
    .in(left_2_3_in),
    .out(left_2_3_out),
    .reset(left_2_3_reset),
    .write_en(left_2_3_write_en)
);
mac_pe pe_2_4 (
    .clk(pe_2_4_clk),
    .done(pe_2_4_done),
    .go(pe_2_4_go),
    .left(pe_2_4_left),
    .mul_ready(pe_2_4_mul_ready),
    .out(pe_2_4_out),
    .reset(pe_2_4_reset),
    .top(pe_2_4_top)
);
std_reg # (
    .WIDTH(32)
) top_2_4 (
    .clk(top_2_4_clk),
    .done(top_2_4_done),
    .in(top_2_4_in),
    .out(top_2_4_out),
    .reset(top_2_4_reset),
    .write_en(top_2_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_4 (
    .clk(left_2_4_clk),
    .done(left_2_4_done),
    .in(left_2_4_in),
    .out(left_2_4_out),
    .reset(left_2_4_reset),
    .write_en(left_2_4_write_en)
);
mac_pe pe_2_5 (
    .clk(pe_2_5_clk),
    .done(pe_2_5_done),
    .go(pe_2_5_go),
    .left(pe_2_5_left),
    .mul_ready(pe_2_5_mul_ready),
    .out(pe_2_5_out),
    .reset(pe_2_5_reset),
    .top(pe_2_5_top)
);
std_reg # (
    .WIDTH(32)
) top_2_5 (
    .clk(top_2_5_clk),
    .done(top_2_5_done),
    .in(top_2_5_in),
    .out(top_2_5_out),
    .reset(top_2_5_reset),
    .write_en(top_2_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_5 (
    .clk(left_2_5_clk),
    .done(left_2_5_done),
    .in(left_2_5_in),
    .out(left_2_5_out),
    .reset(left_2_5_reset),
    .write_en(left_2_5_write_en)
);
mac_pe pe_2_6 (
    .clk(pe_2_6_clk),
    .done(pe_2_6_done),
    .go(pe_2_6_go),
    .left(pe_2_6_left),
    .mul_ready(pe_2_6_mul_ready),
    .out(pe_2_6_out),
    .reset(pe_2_6_reset),
    .top(pe_2_6_top)
);
std_reg # (
    .WIDTH(32)
) top_2_6 (
    .clk(top_2_6_clk),
    .done(top_2_6_done),
    .in(top_2_6_in),
    .out(top_2_6_out),
    .reset(top_2_6_reset),
    .write_en(top_2_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_6 (
    .clk(left_2_6_clk),
    .done(left_2_6_done),
    .in(left_2_6_in),
    .out(left_2_6_out),
    .reset(left_2_6_reset),
    .write_en(left_2_6_write_en)
);
mac_pe pe_2_7 (
    .clk(pe_2_7_clk),
    .done(pe_2_7_done),
    .go(pe_2_7_go),
    .left(pe_2_7_left),
    .mul_ready(pe_2_7_mul_ready),
    .out(pe_2_7_out),
    .reset(pe_2_7_reset),
    .top(pe_2_7_top)
);
std_reg # (
    .WIDTH(32)
) top_2_7 (
    .clk(top_2_7_clk),
    .done(top_2_7_done),
    .in(top_2_7_in),
    .out(top_2_7_out),
    .reset(top_2_7_reset),
    .write_en(top_2_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_7 (
    .clk(left_2_7_clk),
    .done(left_2_7_done),
    .in(left_2_7_in),
    .out(left_2_7_out),
    .reset(left_2_7_reset),
    .write_en(left_2_7_write_en)
);
mac_pe pe_3_0 (
    .clk(pe_3_0_clk),
    .done(pe_3_0_done),
    .go(pe_3_0_go),
    .left(pe_3_0_left),
    .mul_ready(pe_3_0_mul_ready),
    .out(pe_3_0_out),
    .reset(pe_3_0_reset),
    .top(pe_3_0_top)
);
std_reg # (
    .WIDTH(32)
) top_3_0 (
    .clk(top_3_0_clk),
    .done(top_3_0_done),
    .in(top_3_0_in),
    .out(top_3_0_out),
    .reset(top_3_0_reset),
    .write_en(top_3_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_0 (
    .clk(left_3_0_clk),
    .done(left_3_0_done),
    .in(left_3_0_in),
    .out(left_3_0_out),
    .reset(left_3_0_reset),
    .write_en(left_3_0_write_en)
);
mac_pe pe_3_1 (
    .clk(pe_3_1_clk),
    .done(pe_3_1_done),
    .go(pe_3_1_go),
    .left(pe_3_1_left),
    .mul_ready(pe_3_1_mul_ready),
    .out(pe_3_1_out),
    .reset(pe_3_1_reset),
    .top(pe_3_1_top)
);
std_reg # (
    .WIDTH(32)
) top_3_1 (
    .clk(top_3_1_clk),
    .done(top_3_1_done),
    .in(top_3_1_in),
    .out(top_3_1_out),
    .reset(top_3_1_reset),
    .write_en(top_3_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_1 (
    .clk(left_3_1_clk),
    .done(left_3_1_done),
    .in(left_3_1_in),
    .out(left_3_1_out),
    .reset(left_3_1_reset),
    .write_en(left_3_1_write_en)
);
mac_pe pe_3_2 (
    .clk(pe_3_2_clk),
    .done(pe_3_2_done),
    .go(pe_3_2_go),
    .left(pe_3_2_left),
    .mul_ready(pe_3_2_mul_ready),
    .out(pe_3_2_out),
    .reset(pe_3_2_reset),
    .top(pe_3_2_top)
);
std_reg # (
    .WIDTH(32)
) top_3_2 (
    .clk(top_3_2_clk),
    .done(top_3_2_done),
    .in(top_3_2_in),
    .out(top_3_2_out),
    .reset(top_3_2_reset),
    .write_en(top_3_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_2 (
    .clk(left_3_2_clk),
    .done(left_3_2_done),
    .in(left_3_2_in),
    .out(left_3_2_out),
    .reset(left_3_2_reset),
    .write_en(left_3_2_write_en)
);
mac_pe pe_3_3 (
    .clk(pe_3_3_clk),
    .done(pe_3_3_done),
    .go(pe_3_3_go),
    .left(pe_3_3_left),
    .mul_ready(pe_3_3_mul_ready),
    .out(pe_3_3_out),
    .reset(pe_3_3_reset),
    .top(pe_3_3_top)
);
std_reg # (
    .WIDTH(32)
) top_3_3 (
    .clk(top_3_3_clk),
    .done(top_3_3_done),
    .in(top_3_3_in),
    .out(top_3_3_out),
    .reset(top_3_3_reset),
    .write_en(top_3_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_3 (
    .clk(left_3_3_clk),
    .done(left_3_3_done),
    .in(left_3_3_in),
    .out(left_3_3_out),
    .reset(left_3_3_reset),
    .write_en(left_3_3_write_en)
);
mac_pe pe_3_4 (
    .clk(pe_3_4_clk),
    .done(pe_3_4_done),
    .go(pe_3_4_go),
    .left(pe_3_4_left),
    .mul_ready(pe_3_4_mul_ready),
    .out(pe_3_4_out),
    .reset(pe_3_4_reset),
    .top(pe_3_4_top)
);
std_reg # (
    .WIDTH(32)
) top_3_4 (
    .clk(top_3_4_clk),
    .done(top_3_4_done),
    .in(top_3_4_in),
    .out(top_3_4_out),
    .reset(top_3_4_reset),
    .write_en(top_3_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_4 (
    .clk(left_3_4_clk),
    .done(left_3_4_done),
    .in(left_3_4_in),
    .out(left_3_4_out),
    .reset(left_3_4_reset),
    .write_en(left_3_4_write_en)
);
mac_pe pe_3_5 (
    .clk(pe_3_5_clk),
    .done(pe_3_5_done),
    .go(pe_3_5_go),
    .left(pe_3_5_left),
    .mul_ready(pe_3_5_mul_ready),
    .out(pe_3_5_out),
    .reset(pe_3_5_reset),
    .top(pe_3_5_top)
);
std_reg # (
    .WIDTH(32)
) top_3_5 (
    .clk(top_3_5_clk),
    .done(top_3_5_done),
    .in(top_3_5_in),
    .out(top_3_5_out),
    .reset(top_3_5_reset),
    .write_en(top_3_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_5 (
    .clk(left_3_5_clk),
    .done(left_3_5_done),
    .in(left_3_5_in),
    .out(left_3_5_out),
    .reset(left_3_5_reset),
    .write_en(left_3_5_write_en)
);
mac_pe pe_3_6 (
    .clk(pe_3_6_clk),
    .done(pe_3_6_done),
    .go(pe_3_6_go),
    .left(pe_3_6_left),
    .mul_ready(pe_3_6_mul_ready),
    .out(pe_3_6_out),
    .reset(pe_3_6_reset),
    .top(pe_3_6_top)
);
std_reg # (
    .WIDTH(32)
) top_3_6 (
    .clk(top_3_6_clk),
    .done(top_3_6_done),
    .in(top_3_6_in),
    .out(top_3_6_out),
    .reset(top_3_6_reset),
    .write_en(top_3_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_6 (
    .clk(left_3_6_clk),
    .done(left_3_6_done),
    .in(left_3_6_in),
    .out(left_3_6_out),
    .reset(left_3_6_reset),
    .write_en(left_3_6_write_en)
);
mac_pe pe_3_7 (
    .clk(pe_3_7_clk),
    .done(pe_3_7_done),
    .go(pe_3_7_go),
    .left(pe_3_7_left),
    .mul_ready(pe_3_7_mul_ready),
    .out(pe_3_7_out),
    .reset(pe_3_7_reset),
    .top(pe_3_7_top)
);
std_reg # (
    .WIDTH(32)
) top_3_7 (
    .clk(top_3_7_clk),
    .done(top_3_7_done),
    .in(top_3_7_in),
    .out(top_3_7_out),
    .reset(top_3_7_reset),
    .write_en(top_3_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_7 (
    .clk(left_3_7_clk),
    .done(left_3_7_done),
    .in(left_3_7_in),
    .out(left_3_7_out),
    .reset(left_3_7_reset),
    .write_en(left_3_7_write_en)
);
mac_pe pe_4_0 (
    .clk(pe_4_0_clk),
    .done(pe_4_0_done),
    .go(pe_4_0_go),
    .left(pe_4_0_left),
    .mul_ready(pe_4_0_mul_ready),
    .out(pe_4_0_out),
    .reset(pe_4_0_reset),
    .top(pe_4_0_top)
);
std_reg # (
    .WIDTH(32)
) top_4_0 (
    .clk(top_4_0_clk),
    .done(top_4_0_done),
    .in(top_4_0_in),
    .out(top_4_0_out),
    .reset(top_4_0_reset),
    .write_en(top_4_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_0 (
    .clk(left_4_0_clk),
    .done(left_4_0_done),
    .in(left_4_0_in),
    .out(left_4_0_out),
    .reset(left_4_0_reset),
    .write_en(left_4_0_write_en)
);
mac_pe pe_4_1 (
    .clk(pe_4_1_clk),
    .done(pe_4_1_done),
    .go(pe_4_1_go),
    .left(pe_4_1_left),
    .mul_ready(pe_4_1_mul_ready),
    .out(pe_4_1_out),
    .reset(pe_4_1_reset),
    .top(pe_4_1_top)
);
std_reg # (
    .WIDTH(32)
) top_4_1 (
    .clk(top_4_1_clk),
    .done(top_4_1_done),
    .in(top_4_1_in),
    .out(top_4_1_out),
    .reset(top_4_1_reset),
    .write_en(top_4_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_1 (
    .clk(left_4_1_clk),
    .done(left_4_1_done),
    .in(left_4_1_in),
    .out(left_4_1_out),
    .reset(left_4_1_reset),
    .write_en(left_4_1_write_en)
);
mac_pe pe_4_2 (
    .clk(pe_4_2_clk),
    .done(pe_4_2_done),
    .go(pe_4_2_go),
    .left(pe_4_2_left),
    .mul_ready(pe_4_2_mul_ready),
    .out(pe_4_2_out),
    .reset(pe_4_2_reset),
    .top(pe_4_2_top)
);
std_reg # (
    .WIDTH(32)
) top_4_2 (
    .clk(top_4_2_clk),
    .done(top_4_2_done),
    .in(top_4_2_in),
    .out(top_4_2_out),
    .reset(top_4_2_reset),
    .write_en(top_4_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_2 (
    .clk(left_4_2_clk),
    .done(left_4_2_done),
    .in(left_4_2_in),
    .out(left_4_2_out),
    .reset(left_4_2_reset),
    .write_en(left_4_2_write_en)
);
mac_pe pe_4_3 (
    .clk(pe_4_3_clk),
    .done(pe_4_3_done),
    .go(pe_4_3_go),
    .left(pe_4_3_left),
    .mul_ready(pe_4_3_mul_ready),
    .out(pe_4_3_out),
    .reset(pe_4_3_reset),
    .top(pe_4_3_top)
);
std_reg # (
    .WIDTH(32)
) top_4_3 (
    .clk(top_4_3_clk),
    .done(top_4_3_done),
    .in(top_4_3_in),
    .out(top_4_3_out),
    .reset(top_4_3_reset),
    .write_en(top_4_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_3 (
    .clk(left_4_3_clk),
    .done(left_4_3_done),
    .in(left_4_3_in),
    .out(left_4_3_out),
    .reset(left_4_3_reset),
    .write_en(left_4_3_write_en)
);
mac_pe pe_4_4 (
    .clk(pe_4_4_clk),
    .done(pe_4_4_done),
    .go(pe_4_4_go),
    .left(pe_4_4_left),
    .mul_ready(pe_4_4_mul_ready),
    .out(pe_4_4_out),
    .reset(pe_4_4_reset),
    .top(pe_4_4_top)
);
std_reg # (
    .WIDTH(32)
) top_4_4 (
    .clk(top_4_4_clk),
    .done(top_4_4_done),
    .in(top_4_4_in),
    .out(top_4_4_out),
    .reset(top_4_4_reset),
    .write_en(top_4_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_4 (
    .clk(left_4_4_clk),
    .done(left_4_4_done),
    .in(left_4_4_in),
    .out(left_4_4_out),
    .reset(left_4_4_reset),
    .write_en(left_4_4_write_en)
);
mac_pe pe_4_5 (
    .clk(pe_4_5_clk),
    .done(pe_4_5_done),
    .go(pe_4_5_go),
    .left(pe_4_5_left),
    .mul_ready(pe_4_5_mul_ready),
    .out(pe_4_5_out),
    .reset(pe_4_5_reset),
    .top(pe_4_5_top)
);
std_reg # (
    .WIDTH(32)
) top_4_5 (
    .clk(top_4_5_clk),
    .done(top_4_5_done),
    .in(top_4_5_in),
    .out(top_4_5_out),
    .reset(top_4_5_reset),
    .write_en(top_4_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_5 (
    .clk(left_4_5_clk),
    .done(left_4_5_done),
    .in(left_4_5_in),
    .out(left_4_5_out),
    .reset(left_4_5_reset),
    .write_en(left_4_5_write_en)
);
mac_pe pe_4_6 (
    .clk(pe_4_6_clk),
    .done(pe_4_6_done),
    .go(pe_4_6_go),
    .left(pe_4_6_left),
    .mul_ready(pe_4_6_mul_ready),
    .out(pe_4_6_out),
    .reset(pe_4_6_reset),
    .top(pe_4_6_top)
);
std_reg # (
    .WIDTH(32)
) top_4_6 (
    .clk(top_4_6_clk),
    .done(top_4_6_done),
    .in(top_4_6_in),
    .out(top_4_6_out),
    .reset(top_4_6_reset),
    .write_en(top_4_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_6 (
    .clk(left_4_6_clk),
    .done(left_4_6_done),
    .in(left_4_6_in),
    .out(left_4_6_out),
    .reset(left_4_6_reset),
    .write_en(left_4_6_write_en)
);
mac_pe pe_4_7 (
    .clk(pe_4_7_clk),
    .done(pe_4_7_done),
    .go(pe_4_7_go),
    .left(pe_4_7_left),
    .mul_ready(pe_4_7_mul_ready),
    .out(pe_4_7_out),
    .reset(pe_4_7_reset),
    .top(pe_4_7_top)
);
std_reg # (
    .WIDTH(32)
) top_4_7 (
    .clk(top_4_7_clk),
    .done(top_4_7_done),
    .in(top_4_7_in),
    .out(top_4_7_out),
    .reset(top_4_7_reset),
    .write_en(top_4_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_4_7 (
    .clk(left_4_7_clk),
    .done(left_4_7_done),
    .in(left_4_7_in),
    .out(left_4_7_out),
    .reset(left_4_7_reset),
    .write_en(left_4_7_write_en)
);
mac_pe pe_5_0 (
    .clk(pe_5_0_clk),
    .done(pe_5_0_done),
    .go(pe_5_0_go),
    .left(pe_5_0_left),
    .mul_ready(pe_5_0_mul_ready),
    .out(pe_5_0_out),
    .reset(pe_5_0_reset),
    .top(pe_5_0_top)
);
std_reg # (
    .WIDTH(32)
) top_5_0 (
    .clk(top_5_0_clk),
    .done(top_5_0_done),
    .in(top_5_0_in),
    .out(top_5_0_out),
    .reset(top_5_0_reset),
    .write_en(top_5_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_0 (
    .clk(left_5_0_clk),
    .done(left_5_0_done),
    .in(left_5_0_in),
    .out(left_5_0_out),
    .reset(left_5_0_reset),
    .write_en(left_5_0_write_en)
);
mac_pe pe_5_1 (
    .clk(pe_5_1_clk),
    .done(pe_5_1_done),
    .go(pe_5_1_go),
    .left(pe_5_1_left),
    .mul_ready(pe_5_1_mul_ready),
    .out(pe_5_1_out),
    .reset(pe_5_1_reset),
    .top(pe_5_1_top)
);
std_reg # (
    .WIDTH(32)
) top_5_1 (
    .clk(top_5_1_clk),
    .done(top_5_1_done),
    .in(top_5_1_in),
    .out(top_5_1_out),
    .reset(top_5_1_reset),
    .write_en(top_5_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_1 (
    .clk(left_5_1_clk),
    .done(left_5_1_done),
    .in(left_5_1_in),
    .out(left_5_1_out),
    .reset(left_5_1_reset),
    .write_en(left_5_1_write_en)
);
mac_pe pe_5_2 (
    .clk(pe_5_2_clk),
    .done(pe_5_2_done),
    .go(pe_5_2_go),
    .left(pe_5_2_left),
    .mul_ready(pe_5_2_mul_ready),
    .out(pe_5_2_out),
    .reset(pe_5_2_reset),
    .top(pe_5_2_top)
);
std_reg # (
    .WIDTH(32)
) top_5_2 (
    .clk(top_5_2_clk),
    .done(top_5_2_done),
    .in(top_5_2_in),
    .out(top_5_2_out),
    .reset(top_5_2_reset),
    .write_en(top_5_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_2 (
    .clk(left_5_2_clk),
    .done(left_5_2_done),
    .in(left_5_2_in),
    .out(left_5_2_out),
    .reset(left_5_2_reset),
    .write_en(left_5_2_write_en)
);
mac_pe pe_5_3 (
    .clk(pe_5_3_clk),
    .done(pe_5_3_done),
    .go(pe_5_3_go),
    .left(pe_5_3_left),
    .mul_ready(pe_5_3_mul_ready),
    .out(pe_5_3_out),
    .reset(pe_5_3_reset),
    .top(pe_5_3_top)
);
std_reg # (
    .WIDTH(32)
) top_5_3 (
    .clk(top_5_3_clk),
    .done(top_5_3_done),
    .in(top_5_3_in),
    .out(top_5_3_out),
    .reset(top_5_3_reset),
    .write_en(top_5_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_3 (
    .clk(left_5_3_clk),
    .done(left_5_3_done),
    .in(left_5_3_in),
    .out(left_5_3_out),
    .reset(left_5_3_reset),
    .write_en(left_5_3_write_en)
);
mac_pe pe_5_4 (
    .clk(pe_5_4_clk),
    .done(pe_5_4_done),
    .go(pe_5_4_go),
    .left(pe_5_4_left),
    .mul_ready(pe_5_4_mul_ready),
    .out(pe_5_4_out),
    .reset(pe_5_4_reset),
    .top(pe_5_4_top)
);
std_reg # (
    .WIDTH(32)
) top_5_4 (
    .clk(top_5_4_clk),
    .done(top_5_4_done),
    .in(top_5_4_in),
    .out(top_5_4_out),
    .reset(top_5_4_reset),
    .write_en(top_5_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_4 (
    .clk(left_5_4_clk),
    .done(left_5_4_done),
    .in(left_5_4_in),
    .out(left_5_4_out),
    .reset(left_5_4_reset),
    .write_en(left_5_4_write_en)
);
mac_pe pe_5_5 (
    .clk(pe_5_5_clk),
    .done(pe_5_5_done),
    .go(pe_5_5_go),
    .left(pe_5_5_left),
    .mul_ready(pe_5_5_mul_ready),
    .out(pe_5_5_out),
    .reset(pe_5_5_reset),
    .top(pe_5_5_top)
);
std_reg # (
    .WIDTH(32)
) top_5_5 (
    .clk(top_5_5_clk),
    .done(top_5_5_done),
    .in(top_5_5_in),
    .out(top_5_5_out),
    .reset(top_5_5_reset),
    .write_en(top_5_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_5 (
    .clk(left_5_5_clk),
    .done(left_5_5_done),
    .in(left_5_5_in),
    .out(left_5_5_out),
    .reset(left_5_5_reset),
    .write_en(left_5_5_write_en)
);
mac_pe pe_5_6 (
    .clk(pe_5_6_clk),
    .done(pe_5_6_done),
    .go(pe_5_6_go),
    .left(pe_5_6_left),
    .mul_ready(pe_5_6_mul_ready),
    .out(pe_5_6_out),
    .reset(pe_5_6_reset),
    .top(pe_5_6_top)
);
std_reg # (
    .WIDTH(32)
) top_5_6 (
    .clk(top_5_6_clk),
    .done(top_5_6_done),
    .in(top_5_6_in),
    .out(top_5_6_out),
    .reset(top_5_6_reset),
    .write_en(top_5_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_6 (
    .clk(left_5_6_clk),
    .done(left_5_6_done),
    .in(left_5_6_in),
    .out(left_5_6_out),
    .reset(left_5_6_reset),
    .write_en(left_5_6_write_en)
);
mac_pe pe_5_7 (
    .clk(pe_5_7_clk),
    .done(pe_5_7_done),
    .go(pe_5_7_go),
    .left(pe_5_7_left),
    .mul_ready(pe_5_7_mul_ready),
    .out(pe_5_7_out),
    .reset(pe_5_7_reset),
    .top(pe_5_7_top)
);
std_reg # (
    .WIDTH(32)
) top_5_7 (
    .clk(top_5_7_clk),
    .done(top_5_7_done),
    .in(top_5_7_in),
    .out(top_5_7_out),
    .reset(top_5_7_reset),
    .write_en(top_5_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_5_7 (
    .clk(left_5_7_clk),
    .done(left_5_7_done),
    .in(left_5_7_in),
    .out(left_5_7_out),
    .reset(left_5_7_reset),
    .write_en(left_5_7_write_en)
);
mac_pe pe_6_0 (
    .clk(pe_6_0_clk),
    .done(pe_6_0_done),
    .go(pe_6_0_go),
    .left(pe_6_0_left),
    .mul_ready(pe_6_0_mul_ready),
    .out(pe_6_0_out),
    .reset(pe_6_0_reset),
    .top(pe_6_0_top)
);
std_reg # (
    .WIDTH(32)
) top_6_0 (
    .clk(top_6_0_clk),
    .done(top_6_0_done),
    .in(top_6_0_in),
    .out(top_6_0_out),
    .reset(top_6_0_reset),
    .write_en(top_6_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_0 (
    .clk(left_6_0_clk),
    .done(left_6_0_done),
    .in(left_6_0_in),
    .out(left_6_0_out),
    .reset(left_6_0_reset),
    .write_en(left_6_0_write_en)
);
mac_pe pe_6_1 (
    .clk(pe_6_1_clk),
    .done(pe_6_1_done),
    .go(pe_6_1_go),
    .left(pe_6_1_left),
    .mul_ready(pe_6_1_mul_ready),
    .out(pe_6_1_out),
    .reset(pe_6_1_reset),
    .top(pe_6_1_top)
);
std_reg # (
    .WIDTH(32)
) top_6_1 (
    .clk(top_6_1_clk),
    .done(top_6_1_done),
    .in(top_6_1_in),
    .out(top_6_1_out),
    .reset(top_6_1_reset),
    .write_en(top_6_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_1 (
    .clk(left_6_1_clk),
    .done(left_6_1_done),
    .in(left_6_1_in),
    .out(left_6_1_out),
    .reset(left_6_1_reset),
    .write_en(left_6_1_write_en)
);
mac_pe pe_6_2 (
    .clk(pe_6_2_clk),
    .done(pe_6_2_done),
    .go(pe_6_2_go),
    .left(pe_6_2_left),
    .mul_ready(pe_6_2_mul_ready),
    .out(pe_6_2_out),
    .reset(pe_6_2_reset),
    .top(pe_6_2_top)
);
std_reg # (
    .WIDTH(32)
) top_6_2 (
    .clk(top_6_2_clk),
    .done(top_6_2_done),
    .in(top_6_2_in),
    .out(top_6_2_out),
    .reset(top_6_2_reset),
    .write_en(top_6_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_2 (
    .clk(left_6_2_clk),
    .done(left_6_2_done),
    .in(left_6_2_in),
    .out(left_6_2_out),
    .reset(left_6_2_reset),
    .write_en(left_6_2_write_en)
);
mac_pe pe_6_3 (
    .clk(pe_6_3_clk),
    .done(pe_6_3_done),
    .go(pe_6_3_go),
    .left(pe_6_3_left),
    .mul_ready(pe_6_3_mul_ready),
    .out(pe_6_3_out),
    .reset(pe_6_3_reset),
    .top(pe_6_3_top)
);
std_reg # (
    .WIDTH(32)
) top_6_3 (
    .clk(top_6_3_clk),
    .done(top_6_3_done),
    .in(top_6_3_in),
    .out(top_6_3_out),
    .reset(top_6_3_reset),
    .write_en(top_6_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_3 (
    .clk(left_6_3_clk),
    .done(left_6_3_done),
    .in(left_6_3_in),
    .out(left_6_3_out),
    .reset(left_6_3_reset),
    .write_en(left_6_3_write_en)
);
mac_pe pe_6_4 (
    .clk(pe_6_4_clk),
    .done(pe_6_4_done),
    .go(pe_6_4_go),
    .left(pe_6_4_left),
    .mul_ready(pe_6_4_mul_ready),
    .out(pe_6_4_out),
    .reset(pe_6_4_reset),
    .top(pe_6_4_top)
);
std_reg # (
    .WIDTH(32)
) top_6_4 (
    .clk(top_6_4_clk),
    .done(top_6_4_done),
    .in(top_6_4_in),
    .out(top_6_4_out),
    .reset(top_6_4_reset),
    .write_en(top_6_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_4 (
    .clk(left_6_4_clk),
    .done(left_6_4_done),
    .in(left_6_4_in),
    .out(left_6_4_out),
    .reset(left_6_4_reset),
    .write_en(left_6_4_write_en)
);
mac_pe pe_6_5 (
    .clk(pe_6_5_clk),
    .done(pe_6_5_done),
    .go(pe_6_5_go),
    .left(pe_6_5_left),
    .mul_ready(pe_6_5_mul_ready),
    .out(pe_6_5_out),
    .reset(pe_6_5_reset),
    .top(pe_6_5_top)
);
std_reg # (
    .WIDTH(32)
) top_6_5 (
    .clk(top_6_5_clk),
    .done(top_6_5_done),
    .in(top_6_5_in),
    .out(top_6_5_out),
    .reset(top_6_5_reset),
    .write_en(top_6_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_5 (
    .clk(left_6_5_clk),
    .done(left_6_5_done),
    .in(left_6_5_in),
    .out(left_6_5_out),
    .reset(left_6_5_reset),
    .write_en(left_6_5_write_en)
);
mac_pe pe_6_6 (
    .clk(pe_6_6_clk),
    .done(pe_6_6_done),
    .go(pe_6_6_go),
    .left(pe_6_6_left),
    .mul_ready(pe_6_6_mul_ready),
    .out(pe_6_6_out),
    .reset(pe_6_6_reset),
    .top(pe_6_6_top)
);
std_reg # (
    .WIDTH(32)
) top_6_6 (
    .clk(top_6_6_clk),
    .done(top_6_6_done),
    .in(top_6_6_in),
    .out(top_6_6_out),
    .reset(top_6_6_reset),
    .write_en(top_6_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_6 (
    .clk(left_6_6_clk),
    .done(left_6_6_done),
    .in(left_6_6_in),
    .out(left_6_6_out),
    .reset(left_6_6_reset),
    .write_en(left_6_6_write_en)
);
mac_pe pe_6_7 (
    .clk(pe_6_7_clk),
    .done(pe_6_7_done),
    .go(pe_6_7_go),
    .left(pe_6_7_left),
    .mul_ready(pe_6_7_mul_ready),
    .out(pe_6_7_out),
    .reset(pe_6_7_reset),
    .top(pe_6_7_top)
);
std_reg # (
    .WIDTH(32)
) top_6_7 (
    .clk(top_6_7_clk),
    .done(top_6_7_done),
    .in(top_6_7_in),
    .out(top_6_7_out),
    .reset(top_6_7_reset),
    .write_en(top_6_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_6_7 (
    .clk(left_6_7_clk),
    .done(left_6_7_done),
    .in(left_6_7_in),
    .out(left_6_7_out),
    .reset(left_6_7_reset),
    .write_en(left_6_7_write_en)
);
mac_pe pe_7_0 (
    .clk(pe_7_0_clk),
    .done(pe_7_0_done),
    .go(pe_7_0_go),
    .left(pe_7_0_left),
    .mul_ready(pe_7_0_mul_ready),
    .out(pe_7_0_out),
    .reset(pe_7_0_reset),
    .top(pe_7_0_top)
);
std_reg # (
    .WIDTH(32)
) top_7_0 (
    .clk(top_7_0_clk),
    .done(top_7_0_done),
    .in(top_7_0_in),
    .out(top_7_0_out),
    .reset(top_7_0_reset),
    .write_en(top_7_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_0 (
    .clk(left_7_0_clk),
    .done(left_7_0_done),
    .in(left_7_0_in),
    .out(left_7_0_out),
    .reset(left_7_0_reset),
    .write_en(left_7_0_write_en)
);
mac_pe pe_7_1 (
    .clk(pe_7_1_clk),
    .done(pe_7_1_done),
    .go(pe_7_1_go),
    .left(pe_7_1_left),
    .mul_ready(pe_7_1_mul_ready),
    .out(pe_7_1_out),
    .reset(pe_7_1_reset),
    .top(pe_7_1_top)
);
std_reg # (
    .WIDTH(32)
) top_7_1 (
    .clk(top_7_1_clk),
    .done(top_7_1_done),
    .in(top_7_1_in),
    .out(top_7_1_out),
    .reset(top_7_1_reset),
    .write_en(top_7_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_1 (
    .clk(left_7_1_clk),
    .done(left_7_1_done),
    .in(left_7_1_in),
    .out(left_7_1_out),
    .reset(left_7_1_reset),
    .write_en(left_7_1_write_en)
);
mac_pe pe_7_2 (
    .clk(pe_7_2_clk),
    .done(pe_7_2_done),
    .go(pe_7_2_go),
    .left(pe_7_2_left),
    .mul_ready(pe_7_2_mul_ready),
    .out(pe_7_2_out),
    .reset(pe_7_2_reset),
    .top(pe_7_2_top)
);
std_reg # (
    .WIDTH(32)
) top_7_2 (
    .clk(top_7_2_clk),
    .done(top_7_2_done),
    .in(top_7_2_in),
    .out(top_7_2_out),
    .reset(top_7_2_reset),
    .write_en(top_7_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_2 (
    .clk(left_7_2_clk),
    .done(left_7_2_done),
    .in(left_7_2_in),
    .out(left_7_2_out),
    .reset(left_7_2_reset),
    .write_en(left_7_2_write_en)
);
mac_pe pe_7_3 (
    .clk(pe_7_3_clk),
    .done(pe_7_3_done),
    .go(pe_7_3_go),
    .left(pe_7_3_left),
    .mul_ready(pe_7_3_mul_ready),
    .out(pe_7_3_out),
    .reset(pe_7_3_reset),
    .top(pe_7_3_top)
);
std_reg # (
    .WIDTH(32)
) top_7_3 (
    .clk(top_7_3_clk),
    .done(top_7_3_done),
    .in(top_7_3_in),
    .out(top_7_3_out),
    .reset(top_7_3_reset),
    .write_en(top_7_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_3 (
    .clk(left_7_3_clk),
    .done(left_7_3_done),
    .in(left_7_3_in),
    .out(left_7_3_out),
    .reset(left_7_3_reset),
    .write_en(left_7_3_write_en)
);
mac_pe pe_7_4 (
    .clk(pe_7_4_clk),
    .done(pe_7_4_done),
    .go(pe_7_4_go),
    .left(pe_7_4_left),
    .mul_ready(pe_7_4_mul_ready),
    .out(pe_7_4_out),
    .reset(pe_7_4_reset),
    .top(pe_7_4_top)
);
std_reg # (
    .WIDTH(32)
) top_7_4 (
    .clk(top_7_4_clk),
    .done(top_7_4_done),
    .in(top_7_4_in),
    .out(top_7_4_out),
    .reset(top_7_4_reset),
    .write_en(top_7_4_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_4 (
    .clk(left_7_4_clk),
    .done(left_7_4_done),
    .in(left_7_4_in),
    .out(left_7_4_out),
    .reset(left_7_4_reset),
    .write_en(left_7_4_write_en)
);
mac_pe pe_7_5 (
    .clk(pe_7_5_clk),
    .done(pe_7_5_done),
    .go(pe_7_5_go),
    .left(pe_7_5_left),
    .mul_ready(pe_7_5_mul_ready),
    .out(pe_7_5_out),
    .reset(pe_7_5_reset),
    .top(pe_7_5_top)
);
std_reg # (
    .WIDTH(32)
) top_7_5 (
    .clk(top_7_5_clk),
    .done(top_7_5_done),
    .in(top_7_5_in),
    .out(top_7_5_out),
    .reset(top_7_5_reset),
    .write_en(top_7_5_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_5 (
    .clk(left_7_5_clk),
    .done(left_7_5_done),
    .in(left_7_5_in),
    .out(left_7_5_out),
    .reset(left_7_5_reset),
    .write_en(left_7_5_write_en)
);
mac_pe pe_7_6 (
    .clk(pe_7_6_clk),
    .done(pe_7_6_done),
    .go(pe_7_6_go),
    .left(pe_7_6_left),
    .mul_ready(pe_7_6_mul_ready),
    .out(pe_7_6_out),
    .reset(pe_7_6_reset),
    .top(pe_7_6_top)
);
std_reg # (
    .WIDTH(32)
) top_7_6 (
    .clk(top_7_6_clk),
    .done(top_7_6_done),
    .in(top_7_6_in),
    .out(top_7_6_out),
    .reset(top_7_6_reset),
    .write_en(top_7_6_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_6 (
    .clk(left_7_6_clk),
    .done(left_7_6_done),
    .in(left_7_6_in),
    .out(left_7_6_out),
    .reset(left_7_6_reset),
    .write_en(left_7_6_write_en)
);
mac_pe pe_7_7 (
    .clk(pe_7_7_clk),
    .done(pe_7_7_done),
    .go(pe_7_7_go),
    .left(pe_7_7_left),
    .mul_ready(pe_7_7_mul_ready),
    .out(pe_7_7_out),
    .reset(pe_7_7_reset),
    .top(pe_7_7_top)
);
std_reg # (
    .WIDTH(32)
) top_7_7 (
    .clk(top_7_7_clk),
    .done(top_7_7_done),
    .in(top_7_7_in),
    .out(top_7_7_out),
    .reset(top_7_7_reset),
    .write_en(top_7_7_write_en)
);
std_reg # (
    .WIDTH(32)
) left_7_7 (
    .clk(left_7_7_clk),
    .done(left_7_7_done),
    .in(left_7_7_in),
    .out(left_7_7_out),
    .reset(left_7_7_reset),
    .write_en(left_7_7_write_en)
);
std_reg # (
    .WIDTH(4)
) t0_idx (
    .clk(t0_idx_clk),
    .done(t0_idx_done),
    .in(t0_idx_in),
    .out(t0_idx_out),
    .reset(t0_idx_reset),
    .write_en(t0_idx_write_en)
);
std_add # (
    .WIDTH(4)
) t0_add (
    .left(t0_add_left),
    .out(t0_add_out),
    .right(t0_add_right)
);
std_reg # (
    .WIDTH(4)
) t1_idx (
    .clk(t1_idx_clk),
    .done(t1_idx_done),
    .in(t1_idx_in),
    .out(t1_idx_out),
    .reset(t1_idx_reset),
    .write_en(t1_idx_write_en)
);
std_add # (
    .WIDTH(4)
) t1_add (
    .left(t1_add_left),
    .out(t1_add_out),
    .right(t1_add_right)
);
std_reg # (
    .WIDTH(4)
) t2_idx (
    .clk(t2_idx_clk),
    .done(t2_idx_done),
    .in(t2_idx_in),
    .out(t2_idx_out),
    .reset(t2_idx_reset),
    .write_en(t2_idx_write_en)
);
std_add # (
    .WIDTH(4)
) t2_add (
    .left(t2_add_left),
    .out(t2_add_out),
    .right(t2_add_right)
);
std_reg # (
    .WIDTH(4)
) t3_idx (
    .clk(t3_idx_clk),
    .done(t3_idx_done),
    .in(t3_idx_in),
    .out(t3_idx_out),
    .reset(t3_idx_reset),
    .write_en(t3_idx_write_en)
);
std_add # (
    .WIDTH(4)
) t3_add (
    .left(t3_add_left),
    .out(t3_add_out),
    .right(t3_add_right)
);
std_reg # (
    .WIDTH(4)
) t4_idx (
    .clk(t4_idx_clk),
    .done(t4_idx_done),
    .in(t4_idx_in),
    .out(t4_idx_out),
    .reset(t4_idx_reset),
    .write_en(t4_idx_write_en)
);
std_add # (
    .WIDTH(4)
) t4_add (
    .left(t4_add_left),
    .out(t4_add_out),
    .right(t4_add_right)
);
std_reg # (
    .WIDTH(4)
) t5_idx (
    .clk(t5_idx_clk),
    .done(t5_idx_done),
    .in(t5_idx_in),
    .out(t5_idx_out),
    .reset(t5_idx_reset),
    .write_en(t5_idx_write_en)
);
std_add # (
    .WIDTH(4)
) t5_add (
    .left(t5_add_left),
    .out(t5_add_out),
    .right(t5_add_right)
);
std_reg # (
    .WIDTH(4)
) t6_idx (
    .clk(t6_idx_clk),
    .done(t6_idx_done),
    .in(t6_idx_in),
    .out(t6_idx_out),
    .reset(t6_idx_reset),
    .write_en(t6_idx_write_en)
);
std_add # (
    .WIDTH(4)
) t6_add (
    .left(t6_add_left),
    .out(t6_add_out),
    .right(t6_add_right)
);
std_reg # (
    .WIDTH(4)
) t7_idx (
    .clk(t7_idx_clk),
    .done(t7_idx_done),
    .in(t7_idx_in),
    .out(t7_idx_out),
    .reset(t7_idx_reset),
    .write_en(t7_idx_write_en)
);
std_add # (
    .WIDTH(4)
) t7_add (
    .left(t7_add_left),
    .out(t7_add_out),
    .right(t7_add_right)
);
std_reg # (
    .WIDTH(4)
) l0_idx (
    .clk(l0_idx_clk),
    .done(l0_idx_done),
    .in(l0_idx_in),
    .out(l0_idx_out),
    .reset(l0_idx_reset),
    .write_en(l0_idx_write_en)
);
std_add # (
    .WIDTH(4)
) l0_add (
    .left(l0_add_left),
    .out(l0_add_out),
    .right(l0_add_right)
);
std_reg # (
    .WIDTH(4)
) l1_idx (
    .clk(l1_idx_clk),
    .done(l1_idx_done),
    .in(l1_idx_in),
    .out(l1_idx_out),
    .reset(l1_idx_reset),
    .write_en(l1_idx_write_en)
);
std_add # (
    .WIDTH(4)
) l1_add (
    .left(l1_add_left),
    .out(l1_add_out),
    .right(l1_add_right)
);
std_reg # (
    .WIDTH(4)
) l2_idx (
    .clk(l2_idx_clk),
    .done(l2_idx_done),
    .in(l2_idx_in),
    .out(l2_idx_out),
    .reset(l2_idx_reset),
    .write_en(l2_idx_write_en)
);
std_add # (
    .WIDTH(4)
) l2_add (
    .left(l2_add_left),
    .out(l2_add_out),
    .right(l2_add_right)
);
std_reg # (
    .WIDTH(4)
) l3_idx (
    .clk(l3_idx_clk),
    .done(l3_idx_done),
    .in(l3_idx_in),
    .out(l3_idx_out),
    .reset(l3_idx_reset),
    .write_en(l3_idx_write_en)
);
std_add # (
    .WIDTH(4)
) l3_add (
    .left(l3_add_left),
    .out(l3_add_out),
    .right(l3_add_right)
);
std_reg # (
    .WIDTH(4)
) l4_idx (
    .clk(l4_idx_clk),
    .done(l4_idx_done),
    .in(l4_idx_in),
    .out(l4_idx_out),
    .reset(l4_idx_reset),
    .write_en(l4_idx_write_en)
);
std_add # (
    .WIDTH(4)
) l4_add (
    .left(l4_add_left),
    .out(l4_add_out),
    .right(l4_add_right)
);
std_reg # (
    .WIDTH(4)
) l5_idx (
    .clk(l5_idx_clk),
    .done(l5_idx_done),
    .in(l5_idx_in),
    .out(l5_idx_out),
    .reset(l5_idx_reset),
    .write_en(l5_idx_write_en)
);
std_add # (
    .WIDTH(4)
) l5_add (
    .left(l5_add_left),
    .out(l5_add_out),
    .right(l5_add_right)
);
std_reg # (
    .WIDTH(4)
) l6_idx (
    .clk(l6_idx_clk),
    .done(l6_idx_done),
    .in(l6_idx_in),
    .out(l6_idx_out),
    .reset(l6_idx_reset),
    .write_en(l6_idx_write_en)
);
std_add # (
    .WIDTH(4)
) l6_add (
    .left(l6_add_left),
    .out(l6_add_out),
    .right(l6_add_right)
);
std_reg # (
    .WIDTH(4)
) l7_idx (
    .clk(l7_idx_clk),
    .done(l7_idx_done),
    .in(l7_idx_in),
    .out(l7_idx_out),
    .reset(l7_idx_reset),
    .write_en(l7_idx_write_en)
);
std_add # (
    .WIDTH(4)
) l7_add (
    .left(l7_add_left),
    .out(l7_add_out),
    .right(l7_add_right)
);
std_reg # (
    .WIDTH(32)
) idx (
    .clk(idx_clk),
    .done(idx_done),
    .in(idx_in),
    .out(idx_out),
    .reset(idx_reset),
    .write_en(idx_write_en)
);
std_add # (
    .WIDTH(32)
) idx_add (
    .left(idx_add_left),
    .out(idx_add_out),
    .right(idx_add_right)
);
std_lt # (
    .WIDTH(32)
) lt_iter_limit (
    .left(lt_iter_limit_left),
    .out(lt_iter_limit_out),
    .right(lt_iter_limit_right)
);
std_reg # (
    .WIDTH(1)
) cond_reg (
    .clk(cond_reg_clk),
    .done(cond_reg_done),
    .in(cond_reg_in),
    .out(cond_reg_out),
    .reset(cond_reg_reset),
    .write_en(cond_reg_write_en)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_16_depth_plus_17_reg (
    .clk(idx_between_depth_plus_16_depth_plus_17_reg_clk),
    .done(idx_between_depth_plus_16_depth_plus_17_reg_done),
    .in(idx_between_depth_plus_16_depth_plus_17_reg_in),
    .out(idx_between_depth_plus_16_depth_plus_17_reg_out),
    .reset(idx_between_depth_plus_16_depth_plus_17_reg_reset),
    .write_en(idx_between_depth_plus_16_depth_plus_17_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_17 (
    .left(index_lt_depth_plus_17_left),
    .out(index_lt_depth_plus_17_out),
    .right(index_lt_depth_plus_17_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_16 (
    .left(index_ge_depth_plus_16_left),
    .out(index_ge_depth_plus_16_out),
    .right(index_ge_depth_plus_16_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_16_depth_plus_17_comb (
    .left(idx_between_depth_plus_16_depth_plus_17_comb_left),
    .out(idx_between_depth_plus_16_depth_plus_17_comb_out),
    .right(idx_between_depth_plus_16_depth_plus_17_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_12_depth_plus_13_reg (
    .clk(idx_between_depth_plus_12_depth_plus_13_reg_clk),
    .done(idx_between_depth_plus_12_depth_plus_13_reg_done),
    .in(idx_between_depth_plus_12_depth_plus_13_reg_in),
    .out(idx_between_depth_plus_12_depth_plus_13_reg_out),
    .reset(idx_between_depth_plus_12_depth_plus_13_reg_reset),
    .write_en(idx_between_depth_plus_12_depth_plus_13_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_13 (
    .left(index_lt_depth_plus_13_left),
    .out(index_lt_depth_plus_13_out),
    .right(index_lt_depth_plus_13_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_12 (
    .left(index_ge_depth_plus_12_left),
    .out(index_ge_depth_plus_12_out),
    .right(index_ge_depth_plus_12_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_12_depth_plus_13_comb (
    .left(idx_between_depth_plus_12_depth_plus_13_comb_left),
    .out(idx_between_depth_plus_12_depth_plus_13_comb_out),
    .right(idx_between_depth_plus_12_depth_plus_13_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_8_depth_plus_9_reg (
    .clk(idx_between_depth_plus_8_depth_plus_9_reg_clk),
    .done(idx_between_depth_plus_8_depth_plus_9_reg_done),
    .in(idx_between_depth_plus_8_depth_plus_9_reg_in),
    .out(idx_between_depth_plus_8_depth_plus_9_reg_out),
    .reset(idx_between_depth_plus_8_depth_plus_9_reg_reset),
    .write_en(idx_between_depth_plus_8_depth_plus_9_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_9 (
    .left(index_lt_depth_plus_9_left),
    .out(index_lt_depth_plus_9_out),
    .right(index_lt_depth_plus_9_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_8 (
    .left(index_ge_depth_plus_8_left),
    .out(index_ge_depth_plus_8_out),
    .right(index_ge_depth_plus_8_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_8_depth_plus_9_comb (
    .left(idx_between_depth_plus_8_depth_plus_9_comb_left),
    .out(idx_between_depth_plus_8_depth_plus_9_comb_out),
    .right(idx_between_depth_plus_8_depth_plus_9_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_2_min_depth_4_plus_2_reg (
    .clk(idx_between_2_min_depth_4_plus_2_reg_clk),
    .done(idx_between_2_min_depth_4_plus_2_reg_done),
    .in(idx_between_2_min_depth_4_plus_2_reg_in),
    .out(idx_between_2_min_depth_4_plus_2_reg_out),
    .reset(idx_between_2_min_depth_4_plus_2_reg_reset),
    .write_en(idx_between_2_min_depth_4_plus_2_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_2 (
    .left(index_lt_min_depth_4_plus_2_left),
    .out(index_lt_min_depth_4_plus_2_out),
    .right(index_lt_min_depth_4_plus_2_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_2 (
    .left(index_ge_2_left),
    .out(index_ge_2_out),
    .right(index_ge_2_right)
);
std_and # (
    .WIDTH(1)
) idx_between_2_min_depth_4_plus_2_comb (
    .left(idx_between_2_min_depth_4_plus_2_comb_left),
    .out(idx_between_2_min_depth_4_plus_2_comb_out),
    .right(idx_between_2_min_depth_4_plus_2_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_2_depth_plus_2_reg (
    .clk(idx_between_2_depth_plus_2_reg_clk),
    .done(idx_between_2_depth_plus_2_reg_done),
    .in(idx_between_2_depth_plus_2_reg_in),
    .out(idx_between_2_depth_plus_2_reg_out),
    .reset(idx_between_2_depth_plus_2_reg_reset),
    .write_en(idx_between_2_depth_plus_2_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_2 (
    .left(index_lt_depth_plus_2_left),
    .out(index_lt_depth_plus_2_out),
    .right(index_lt_depth_plus_2_right)
);
std_and # (
    .WIDTH(1)
) idx_between_2_depth_plus_2_comb (
    .left(idx_between_2_depth_plus_2_comb_left),
    .out(idx_between_2_depth_plus_2_comb_out),
    .right(idx_between_2_depth_plus_2_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_17_depth_plus_18_reg (
    .clk(idx_between_depth_plus_17_depth_plus_18_reg_clk),
    .done(idx_between_depth_plus_17_depth_plus_18_reg_done),
    .in(idx_between_depth_plus_17_depth_plus_18_reg_in),
    .out(idx_between_depth_plus_17_depth_plus_18_reg_out),
    .reset(idx_between_depth_plus_17_depth_plus_18_reg_reset),
    .write_en(idx_between_depth_plus_17_depth_plus_18_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_18 (
    .left(index_lt_depth_plus_18_left),
    .out(index_lt_depth_plus_18_out),
    .right(index_lt_depth_plus_18_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_17 (
    .left(index_ge_depth_plus_17_left),
    .out(index_ge_depth_plus_17_out),
    .right(index_ge_depth_plus_17_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_17_depth_plus_18_comb (
    .left(idx_between_depth_plus_17_depth_plus_18_comb_left),
    .out(idx_between_depth_plus_17_depth_plus_18_comb_out),
    .right(idx_between_depth_plus_17_depth_plus_18_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_11_depth_plus_11_reg (
    .clk(idx_between_11_depth_plus_11_reg_clk),
    .done(idx_between_11_depth_plus_11_reg_done),
    .in(idx_between_11_depth_plus_11_reg_in),
    .out(idx_between_11_depth_plus_11_reg_out),
    .reset(idx_between_11_depth_plus_11_reg_reset),
    .write_en(idx_between_11_depth_plus_11_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_11 (
    .left(index_lt_depth_plus_11_left),
    .out(index_lt_depth_plus_11_out),
    .right(index_lt_depth_plus_11_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_11 (
    .left(index_ge_11_left),
    .out(index_ge_11_out),
    .right(index_ge_11_right)
);
std_and # (
    .WIDTH(1)
) idx_between_11_depth_plus_11_comb (
    .left(idx_between_11_depth_plus_11_comb_left),
    .out(idx_between_11_depth_plus_11_comb_out),
    .right(idx_between_11_depth_plus_11_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_11_min_depth_4_plus_11_reg (
    .clk(idx_between_11_min_depth_4_plus_11_reg_clk),
    .done(idx_between_11_min_depth_4_plus_11_reg_done),
    .in(idx_between_11_min_depth_4_plus_11_reg_in),
    .out(idx_between_11_min_depth_4_plus_11_reg_out),
    .reset(idx_between_11_min_depth_4_plus_11_reg_reset),
    .write_en(idx_between_11_min_depth_4_plus_11_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_11 (
    .left(index_lt_min_depth_4_plus_11_left),
    .out(index_lt_min_depth_4_plus_11_out),
    .right(index_lt_min_depth_4_plus_11_right)
);
std_and # (
    .WIDTH(1)
) idx_between_11_min_depth_4_plus_11_comb (
    .left(idx_between_11_min_depth_4_plus_11_comb_left),
    .out(idx_between_11_min_depth_4_plus_11_comb_out),
    .right(idx_between_11_min_depth_4_plus_11_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_13_depth_plus_14_reg (
    .clk(idx_between_depth_plus_13_depth_plus_14_reg_clk),
    .done(idx_between_depth_plus_13_depth_plus_14_reg_done),
    .in(idx_between_depth_plus_13_depth_plus_14_reg_in),
    .out(idx_between_depth_plus_13_depth_plus_14_reg_out),
    .reset(idx_between_depth_plus_13_depth_plus_14_reg_reset),
    .write_en(idx_between_depth_plus_13_depth_plus_14_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_14 (
    .left(index_lt_depth_plus_14_left),
    .out(index_lt_depth_plus_14_out),
    .right(index_lt_depth_plus_14_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_13 (
    .left(index_ge_depth_plus_13_left),
    .out(index_ge_depth_plus_13_out),
    .right(index_ge_depth_plus_13_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_13_depth_plus_14_comb (
    .left(idx_between_depth_plus_13_depth_plus_14_comb_left),
    .out(idx_between_depth_plus_13_depth_plus_14_comb_out),
    .right(idx_between_depth_plus_13_depth_plus_14_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_7_depth_plus_7_reg (
    .clk(idx_between_7_depth_plus_7_reg_clk),
    .done(idx_between_7_depth_plus_7_reg_done),
    .in(idx_between_7_depth_plus_7_reg_in),
    .out(idx_between_7_depth_plus_7_reg_out),
    .reset(idx_between_7_depth_plus_7_reg_reset),
    .write_en(idx_between_7_depth_plus_7_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_7 (
    .left(index_lt_depth_plus_7_left),
    .out(index_lt_depth_plus_7_out),
    .right(index_lt_depth_plus_7_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_7 (
    .left(index_ge_7_left),
    .out(index_ge_7_out),
    .right(index_ge_7_right)
);
std_and # (
    .WIDTH(1)
) idx_between_7_depth_plus_7_comb (
    .left(idx_between_7_depth_plus_7_comb_left),
    .out(idx_between_7_depth_plus_7_comb_out),
    .right(idx_between_7_depth_plus_7_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_7_min_depth_4_plus_7_reg (
    .clk(idx_between_7_min_depth_4_plus_7_reg_clk),
    .done(idx_between_7_min_depth_4_plus_7_reg_done),
    .in(idx_between_7_min_depth_4_plus_7_reg_in),
    .out(idx_between_7_min_depth_4_plus_7_reg_out),
    .reset(idx_between_7_min_depth_4_plus_7_reg_reset),
    .write_en(idx_between_7_min_depth_4_plus_7_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_7 (
    .left(index_lt_min_depth_4_plus_7_left),
    .out(index_lt_min_depth_4_plus_7_out),
    .right(index_lt_min_depth_4_plus_7_right)
);
std_and # (
    .WIDTH(1)
) idx_between_7_min_depth_4_plus_7_comb (
    .left(idx_between_7_min_depth_4_plus_7_comb_left),
    .out(idx_between_7_min_depth_4_plus_7_comb_out),
    .right(idx_between_7_min_depth_4_plus_7_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_16_depth_plus_16_reg (
    .clk(idx_between_16_depth_plus_16_reg_clk),
    .done(idx_between_16_depth_plus_16_reg_done),
    .in(idx_between_16_depth_plus_16_reg_in),
    .out(idx_between_16_depth_plus_16_reg_out),
    .reset(idx_between_16_depth_plus_16_reg_reset),
    .write_en(idx_between_16_depth_plus_16_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_16 (
    .left(index_lt_depth_plus_16_left),
    .out(index_lt_depth_plus_16_out),
    .right(index_lt_depth_plus_16_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_16 (
    .left(index_ge_16_left),
    .out(index_ge_16_out),
    .right(index_ge_16_right)
);
std_and # (
    .WIDTH(1)
) idx_between_16_depth_plus_16_comb (
    .left(idx_between_16_depth_plus_16_comb_left),
    .out(idx_between_16_depth_plus_16_comb_out),
    .right(idx_between_16_depth_plus_16_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_18_depth_plus_19_reg (
    .clk(idx_between_depth_plus_18_depth_plus_19_reg_clk),
    .done(idx_between_depth_plus_18_depth_plus_19_reg_done),
    .in(idx_between_depth_plus_18_depth_plus_19_reg_in),
    .out(idx_between_depth_plus_18_depth_plus_19_reg_out),
    .reset(idx_between_depth_plus_18_depth_plus_19_reg_reset),
    .write_en(idx_between_depth_plus_18_depth_plus_19_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_19 (
    .left(index_lt_depth_plus_19_left),
    .out(index_lt_depth_plus_19_out),
    .right(index_lt_depth_plus_19_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_18 (
    .left(index_ge_depth_plus_18_left),
    .out(index_ge_depth_plus_18_out),
    .right(index_ge_depth_plus_18_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_18_depth_plus_19_comb (
    .left(idx_between_depth_plus_18_depth_plus_19_comb_left),
    .out(idx_between_depth_plus_18_depth_plus_19_comb_out),
    .right(idx_between_depth_plus_18_depth_plus_19_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_3_depth_plus_3_reg (
    .clk(idx_between_3_depth_plus_3_reg_clk),
    .done(idx_between_3_depth_plus_3_reg_done),
    .in(idx_between_3_depth_plus_3_reg_in),
    .out(idx_between_3_depth_plus_3_reg_out),
    .reset(idx_between_3_depth_plus_3_reg_reset),
    .write_en(idx_between_3_depth_plus_3_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_3 (
    .left(index_lt_depth_plus_3_left),
    .out(index_lt_depth_plus_3_out),
    .right(index_lt_depth_plus_3_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_3 (
    .left(index_ge_3_left),
    .out(index_ge_3_out),
    .right(index_ge_3_right)
);
std_and # (
    .WIDTH(1)
) idx_between_3_depth_plus_3_comb (
    .left(idx_between_3_depth_plus_3_comb_left),
    .out(idx_between_3_depth_plus_3_comb_out),
    .right(idx_between_3_depth_plus_3_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_12_depth_plus_12_reg (
    .clk(idx_between_12_depth_plus_12_reg_clk),
    .done(idx_between_12_depth_plus_12_reg_done),
    .in(idx_between_12_depth_plus_12_reg_in),
    .out(idx_between_12_depth_plus_12_reg_out),
    .reset(idx_between_12_depth_plus_12_reg_reset),
    .write_en(idx_between_12_depth_plus_12_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_12 (
    .left(index_lt_depth_plus_12_left),
    .out(index_lt_depth_plus_12_out),
    .right(index_lt_depth_plus_12_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_12 (
    .left(index_ge_12_left),
    .out(index_ge_12_out),
    .right(index_ge_12_right)
);
std_and # (
    .WIDTH(1)
) idx_between_12_depth_plus_12_comb (
    .left(idx_between_12_depth_plus_12_comb_left),
    .out(idx_between_12_depth_plus_12_comb_out),
    .right(idx_between_12_depth_plus_12_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_3_min_depth_4_plus_3_reg (
    .clk(idx_between_3_min_depth_4_plus_3_reg_clk),
    .done(idx_between_3_min_depth_4_plus_3_reg_done),
    .in(idx_between_3_min_depth_4_plus_3_reg_in),
    .out(idx_between_3_min_depth_4_plus_3_reg_out),
    .reset(idx_between_3_min_depth_4_plus_3_reg_reset),
    .write_en(idx_between_3_min_depth_4_plus_3_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_3 (
    .left(index_lt_min_depth_4_plus_3_left),
    .out(index_lt_min_depth_4_plus_3_out),
    .right(index_lt_min_depth_4_plus_3_right)
);
std_and # (
    .WIDTH(1)
) idx_between_3_min_depth_4_plus_3_comb (
    .left(idx_between_3_min_depth_4_plus_3_comb_left),
    .out(idx_between_3_min_depth_4_plus_3_comb_out),
    .right(idx_between_3_min_depth_4_plus_3_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_12_min_depth_4_plus_12_reg (
    .clk(idx_between_12_min_depth_4_plus_12_reg_clk),
    .done(idx_between_12_min_depth_4_plus_12_reg_done),
    .in(idx_between_12_min_depth_4_plus_12_reg_in),
    .out(idx_between_12_min_depth_4_plus_12_reg_out),
    .reset(idx_between_12_min_depth_4_plus_12_reg_reset),
    .write_en(idx_between_12_min_depth_4_plus_12_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_12 (
    .left(index_lt_min_depth_4_plus_12_left),
    .out(index_lt_min_depth_4_plus_12_out),
    .right(index_lt_min_depth_4_plus_12_right)
);
std_and # (
    .WIDTH(1)
) idx_between_12_min_depth_4_plus_12_comb (
    .left(idx_between_12_min_depth_4_plus_12_comb_left),
    .out(idx_between_12_min_depth_4_plus_12_comb_out),
    .right(idx_between_12_min_depth_4_plus_12_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_5_depth_plus_6_reg (
    .clk(idx_between_depth_plus_5_depth_plus_6_reg_clk),
    .done(idx_between_depth_plus_5_depth_plus_6_reg_done),
    .in(idx_between_depth_plus_5_depth_plus_6_reg_in),
    .out(idx_between_depth_plus_5_depth_plus_6_reg_out),
    .reset(idx_between_depth_plus_5_depth_plus_6_reg_reset),
    .write_en(idx_between_depth_plus_5_depth_plus_6_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_6 (
    .left(index_lt_depth_plus_6_left),
    .out(index_lt_depth_plus_6_out),
    .right(index_lt_depth_plus_6_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_5 (
    .left(index_ge_depth_plus_5_left),
    .out(index_ge_depth_plus_5_out),
    .right(index_ge_depth_plus_5_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_5_depth_plus_6_comb (
    .left(idx_between_depth_plus_5_depth_plus_6_comb_left),
    .out(idx_between_depth_plus_5_depth_plus_6_comb_out),
    .right(idx_between_depth_plus_5_depth_plus_6_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_14_depth_plus_15_reg (
    .clk(idx_between_depth_plus_14_depth_plus_15_reg_clk),
    .done(idx_between_depth_plus_14_depth_plus_15_reg_done),
    .in(idx_between_depth_plus_14_depth_plus_15_reg_in),
    .out(idx_between_depth_plus_14_depth_plus_15_reg_out),
    .reset(idx_between_depth_plus_14_depth_plus_15_reg_reset),
    .write_en(idx_between_depth_plus_14_depth_plus_15_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_15 (
    .left(index_lt_depth_plus_15_left),
    .out(index_lt_depth_plus_15_out),
    .right(index_lt_depth_plus_15_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_14 (
    .left(index_ge_depth_plus_14_left),
    .out(index_ge_depth_plus_14_out),
    .right(index_ge_depth_plus_14_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_14_depth_plus_15_comb (
    .left(idx_between_depth_plus_14_depth_plus_15_comb_left),
    .out(idx_between_depth_plus_14_depth_plus_15_comb_out),
    .right(idx_between_depth_plus_14_depth_plus_15_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_9_depth_plus_10_reg (
    .clk(idx_between_depth_plus_9_depth_plus_10_reg_clk),
    .done(idx_between_depth_plus_9_depth_plus_10_reg_done),
    .in(idx_between_depth_plus_9_depth_plus_10_reg_in),
    .out(idx_between_depth_plus_9_depth_plus_10_reg_out),
    .reset(idx_between_depth_plus_9_depth_plus_10_reg_reset),
    .write_en(idx_between_depth_plus_9_depth_plus_10_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_10 (
    .left(index_lt_depth_plus_10_left),
    .out(index_lt_depth_plus_10_out),
    .right(index_lt_depth_plus_10_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_9 (
    .left(index_ge_depth_plus_9_left),
    .out(index_ge_depth_plus_9_out),
    .right(index_ge_depth_plus_9_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_9_depth_plus_10_comb (
    .left(idx_between_depth_plus_9_depth_plus_10_comb_left),
    .out(idx_between_depth_plus_9_depth_plus_10_comb_out),
    .right(idx_between_depth_plus_9_depth_plus_10_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_8_depth_plus_8_reg (
    .clk(idx_between_8_depth_plus_8_reg_clk),
    .done(idx_between_8_depth_plus_8_reg_done),
    .in(idx_between_8_depth_plus_8_reg_in),
    .out(idx_between_8_depth_plus_8_reg_out),
    .reset(idx_between_8_depth_plus_8_reg_reset),
    .write_en(idx_between_8_depth_plus_8_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_8 (
    .left(index_lt_depth_plus_8_left),
    .out(index_lt_depth_plus_8_out),
    .right(index_lt_depth_plus_8_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_8 (
    .left(index_ge_8_left),
    .out(index_ge_8_out),
    .right(index_ge_8_right)
);
std_and # (
    .WIDTH(1)
) idx_between_8_depth_plus_8_comb (
    .left(idx_between_8_depth_plus_8_comb_left),
    .out(idx_between_8_depth_plus_8_comb_out),
    .right(idx_between_8_depth_plus_8_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_8_min_depth_4_plus_8_reg (
    .clk(idx_between_8_min_depth_4_plus_8_reg_clk),
    .done(idx_between_8_min_depth_4_plus_8_reg_done),
    .in(idx_between_8_min_depth_4_plus_8_reg_in),
    .out(idx_between_8_min_depth_4_plus_8_reg_out),
    .reset(idx_between_8_min_depth_4_plus_8_reg_reset),
    .write_en(idx_between_8_min_depth_4_plus_8_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_8 (
    .left(index_lt_min_depth_4_plus_8_left),
    .out(index_lt_min_depth_4_plus_8_out),
    .right(index_lt_min_depth_4_plus_8_right)
);
std_and # (
    .WIDTH(1)
) idx_between_8_min_depth_4_plus_8_comb (
    .left(idx_between_8_min_depth_4_plus_8_comb_left),
    .out(idx_between_8_min_depth_4_plus_8_comb_out),
    .right(idx_between_8_min_depth_4_plus_8_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_17_depth_plus_17_reg (
    .clk(idx_between_17_depth_plus_17_reg_clk),
    .done(idx_between_17_depth_plus_17_reg_done),
    .in(idx_between_17_depth_plus_17_reg_in),
    .out(idx_between_17_depth_plus_17_reg_out),
    .reset(idx_between_17_depth_plus_17_reg_reset),
    .write_en(idx_between_17_depth_plus_17_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_17 (
    .left(index_ge_17_left),
    .out(index_ge_17_out),
    .right(index_ge_17_right)
);
std_and # (
    .WIDTH(1)
) idx_between_17_depth_plus_17_comb (
    .left(idx_between_17_depth_plus_17_comb_left),
    .out(idx_between_17_depth_plus_17_comb_out),
    .right(idx_between_17_depth_plus_17_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_10_depth_plus_11_reg (
    .clk(idx_between_depth_plus_10_depth_plus_11_reg_clk),
    .done(idx_between_depth_plus_10_depth_plus_11_reg_done),
    .in(idx_between_depth_plus_10_depth_plus_11_reg_in),
    .out(idx_between_depth_plus_10_depth_plus_11_reg_out),
    .reset(idx_between_depth_plus_10_depth_plus_11_reg_reset),
    .write_en(idx_between_depth_plus_10_depth_plus_11_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_10 (
    .left(index_ge_depth_plus_10_left),
    .out(index_ge_depth_plus_10_out),
    .right(index_ge_depth_plus_10_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_10_depth_plus_11_comb (
    .left(idx_between_depth_plus_10_depth_plus_11_comb_left),
    .out(idx_between_depth_plus_10_depth_plus_11_comb_out),
    .right(idx_between_depth_plus_10_depth_plus_11_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_19_depth_plus_20_reg (
    .clk(idx_between_depth_plus_19_depth_plus_20_reg_clk),
    .done(idx_between_depth_plus_19_depth_plus_20_reg_done),
    .in(idx_between_depth_plus_19_depth_plus_20_reg_in),
    .out(idx_between_depth_plus_19_depth_plus_20_reg_out),
    .reset(idx_between_depth_plus_19_depth_plus_20_reg_reset),
    .write_en(idx_between_depth_plus_19_depth_plus_20_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_20 (
    .left(index_lt_depth_plus_20_left),
    .out(index_lt_depth_plus_20_out),
    .right(index_lt_depth_plus_20_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_19 (
    .left(index_ge_depth_plus_19_left),
    .out(index_ge_depth_plus_19_out),
    .right(index_ge_depth_plus_19_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_19_depth_plus_20_comb (
    .left(idx_between_depth_plus_19_depth_plus_20_comb_left),
    .out(idx_between_depth_plus_19_depth_plus_20_comb_out),
    .right(idx_between_depth_plus_19_depth_plus_20_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_6_min_depth_4_plus_6_reg (
    .clk(idx_between_6_min_depth_4_plus_6_reg_clk),
    .done(idx_between_6_min_depth_4_plus_6_reg_done),
    .in(idx_between_6_min_depth_4_plus_6_reg_in),
    .out(idx_between_6_min_depth_4_plus_6_reg_out),
    .reset(idx_between_6_min_depth_4_plus_6_reg_reset),
    .write_en(idx_between_6_min_depth_4_plus_6_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_6 (
    .left(index_lt_min_depth_4_plus_6_left),
    .out(index_lt_min_depth_4_plus_6_out),
    .right(index_lt_min_depth_4_plus_6_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_6 (
    .left(index_ge_6_left),
    .out(index_ge_6_out),
    .right(index_ge_6_right)
);
std_and # (
    .WIDTH(1)
) idx_between_6_min_depth_4_plus_6_comb (
    .left(idx_between_6_min_depth_4_plus_6_comb_left),
    .out(idx_between_6_min_depth_4_plus_6_comb_out),
    .right(idx_between_6_min_depth_4_plus_6_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_13_depth_plus_13_reg (
    .clk(idx_between_13_depth_plus_13_reg_clk),
    .done(idx_between_13_depth_plus_13_reg_done),
    .in(idx_between_13_depth_plus_13_reg_in),
    .out(idx_between_13_depth_plus_13_reg_out),
    .reset(idx_between_13_depth_plus_13_reg_reset),
    .write_en(idx_between_13_depth_plus_13_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_13 (
    .left(index_ge_13_left),
    .out(index_ge_13_out),
    .right(index_ge_13_right)
);
std_and # (
    .WIDTH(1)
) idx_between_13_depth_plus_13_comb (
    .left(idx_between_13_depth_plus_13_comb_left),
    .out(idx_between_13_depth_plus_13_comb_out),
    .right(idx_between_13_depth_plus_13_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_13_min_depth_4_plus_13_reg (
    .clk(idx_between_13_min_depth_4_plus_13_reg_clk),
    .done(idx_between_13_min_depth_4_plus_13_reg_done),
    .in(idx_between_13_min_depth_4_plus_13_reg_in),
    .out(idx_between_13_min_depth_4_plus_13_reg_out),
    .reset(idx_between_13_min_depth_4_plus_13_reg_reset),
    .write_en(idx_between_13_min_depth_4_plus_13_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_13 (
    .left(index_lt_min_depth_4_plus_13_left),
    .out(index_lt_min_depth_4_plus_13_out),
    .right(index_lt_min_depth_4_plus_13_right)
);
std_and # (
    .WIDTH(1)
) idx_between_13_min_depth_4_plus_13_comb (
    .left(idx_between_13_min_depth_4_plus_13_comb_left),
    .out(idx_between_13_min_depth_4_plus_13_comb_out),
    .right(idx_between_13_min_depth_4_plus_13_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_6_depth_plus_7_reg (
    .clk(idx_between_depth_plus_6_depth_plus_7_reg_clk),
    .done(idx_between_depth_plus_6_depth_plus_7_reg_done),
    .in(idx_between_depth_plus_6_depth_plus_7_reg_in),
    .out(idx_between_depth_plus_6_depth_plus_7_reg_out),
    .reset(idx_between_depth_plus_6_depth_plus_7_reg_reset),
    .write_en(idx_between_depth_plus_6_depth_plus_7_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_6 (
    .left(index_ge_depth_plus_6_left),
    .out(index_ge_depth_plus_6_out),
    .right(index_ge_depth_plus_6_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_6_depth_plus_7_comb (
    .left(idx_between_depth_plus_6_depth_plus_7_comb_left),
    .out(idx_between_depth_plus_6_depth_plus_7_comb_out),
    .right(idx_between_depth_plus_6_depth_plus_7_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_15_depth_plus_16_reg (
    .clk(idx_between_depth_plus_15_depth_plus_16_reg_clk),
    .done(idx_between_depth_plus_15_depth_plus_16_reg_done),
    .in(idx_between_depth_plus_15_depth_plus_16_reg_in),
    .out(idx_between_depth_plus_15_depth_plus_16_reg_out),
    .reset(idx_between_depth_plus_15_depth_plus_16_reg_reset),
    .write_en(idx_between_depth_plus_15_depth_plus_16_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_15 (
    .left(index_ge_depth_plus_15_left),
    .out(index_ge_depth_plus_15_out),
    .right(index_ge_depth_plus_15_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_15_depth_plus_16_comb (
    .left(idx_between_depth_plus_15_depth_plus_16_comb_left),
    .out(idx_between_depth_plus_15_depth_plus_16_comb_out),
    .right(idx_between_depth_plus_15_depth_plus_16_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_18_depth_plus_18_reg (
    .clk(idx_between_18_depth_plus_18_reg_clk),
    .done(idx_between_18_depth_plus_18_reg_done),
    .in(idx_between_18_depth_plus_18_reg_in),
    .out(idx_between_18_depth_plus_18_reg_out),
    .reset(idx_between_18_depth_plus_18_reg_reset),
    .write_en(idx_between_18_depth_plus_18_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_18 (
    .left(index_ge_18_left),
    .out(index_ge_18_out),
    .right(index_ge_18_right)
);
std_and # (
    .WIDTH(1)
) idx_between_18_depth_plus_18_comb (
    .left(idx_between_18_depth_plus_18_comb_left),
    .out(idx_between_18_depth_plus_18_comb_out),
    .right(idx_between_18_depth_plus_18_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_15_depth_plus_15_reg (
    .clk(idx_between_15_depth_plus_15_reg_clk),
    .done(idx_between_15_depth_plus_15_reg_done),
    .in(idx_between_15_depth_plus_15_reg_in),
    .out(idx_between_15_depth_plus_15_reg_out),
    .reset(idx_between_15_depth_plus_15_reg_reset),
    .write_en(idx_between_15_depth_plus_15_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_15 (
    .left(index_ge_15_left),
    .out(index_ge_15_out),
    .right(index_ge_15_right)
);
std_and # (
    .WIDTH(1)
) idx_between_15_depth_plus_15_comb (
    .left(idx_between_15_depth_plus_15_comb_left),
    .out(idx_between_15_depth_plus_15_comb_out),
    .right(idx_between_15_depth_plus_15_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_4_depth_plus_4_reg (
    .clk(idx_between_4_depth_plus_4_reg_clk),
    .done(idx_between_4_depth_plus_4_reg_done),
    .in(idx_between_4_depth_plus_4_reg_in),
    .out(idx_between_4_depth_plus_4_reg_out),
    .reset(idx_between_4_depth_plus_4_reg_reset),
    .write_en(idx_between_4_depth_plus_4_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_4 (
    .left(index_lt_depth_plus_4_left),
    .out(index_lt_depth_plus_4_out),
    .right(index_lt_depth_plus_4_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_4 (
    .left(index_ge_4_left),
    .out(index_ge_4_out),
    .right(index_ge_4_right)
);
std_and # (
    .WIDTH(1)
) idx_between_4_depth_plus_4_comb (
    .left(idx_between_4_depth_plus_4_comb_left),
    .out(idx_between_4_depth_plus_4_comb_out),
    .right(idx_between_4_depth_plus_4_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_4_min_depth_4_plus_4_reg (
    .clk(idx_between_4_min_depth_4_plus_4_reg_clk),
    .done(idx_between_4_min_depth_4_plus_4_reg_done),
    .in(idx_between_4_min_depth_4_plus_4_reg_in),
    .out(idx_between_4_min_depth_4_plus_4_reg_out),
    .reset(idx_between_4_min_depth_4_plus_4_reg_reset),
    .write_en(idx_between_4_min_depth_4_plus_4_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_4 (
    .left(index_lt_min_depth_4_plus_4_left),
    .out(index_lt_min_depth_4_plus_4_out),
    .right(index_lt_min_depth_4_plus_4_right)
);
std_and # (
    .WIDTH(1)
) idx_between_4_min_depth_4_plus_4_comb (
    .left(idx_between_4_min_depth_4_plus_4_comb_left),
    .out(idx_between_4_min_depth_4_plus_4_comb_out),
    .right(idx_between_4_min_depth_4_plus_4_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_5_depth_plus_5_reg (
    .clk(idx_between_5_depth_plus_5_reg_clk),
    .done(idx_between_5_depth_plus_5_reg_done),
    .in(idx_between_5_depth_plus_5_reg_in),
    .out(idx_between_5_depth_plus_5_reg_out),
    .reset(idx_between_5_depth_plus_5_reg_reset),
    .write_en(idx_between_5_depth_plus_5_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_5 (
    .left(index_lt_depth_plus_5_left),
    .out(index_lt_depth_plus_5_out),
    .right(index_lt_depth_plus_5_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_5 (
    .left(index_ge_5_left),
    .out(index_ge_5_out),
    .right(index_ge_5_right)
);
std_and # (
    .WIDTH(1)
) idx_between_5_depth_plus_5_comb (
    .left(idx_between_5_depth_plus_5_comb_left),
    .out(idx_between_5_depth_plus_5_comb_out),
    .right(idx_between_5_depth_plus_5_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_14_depth_plus_14_reg (
    .clk(idx_between_14_depth_plus_14_reg_clk),
    .done(idx_between_14_depth_plus_14_reg_done),
    .in(idx_between_14_depth_plus_14_reg_in),
    .out(idx_between_14_depth_plus_14_reg_out),
    .reset(idx_between_14_depth_plus_14_reg_reset),
    .write_en(idx_between_14_depth_plus_14_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_14 (
    .left(index_ge_14_left),
    .out(index_ge_14_out),
    .right(index_ge_14_right)
);
std_and # (
    .WIDTH(1)
) idx_between_14_depth_plus_14_comb (
    .left(idx_between_14_depth_plus_14_comb_left),
    .out(idx_between_14_depth_plus_14_comb_out),
    .right(idx_between_14_depth_plus_14_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_5_min_depth_4_plus_5_reg (
    .clk(idx_between_5_min_depth_4_plus_5_reg_clk),
    .done(idx_between_5_min_depth_4_plus_5_reg_done),
    .in(idx_between_5_min_depth_4_plus_5_reg_in),
    .out(idx_between_5_min_depth_4_plus_5_reg_out),
    .reset(idx_between_5_min_depth_4_plus_5_reg_reset),
    .write_en(idx_between_5_min_depth_4_plus_5_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_5 (
    .left(index_lt_min_depth_4_plus_5_left),
    .out(index_lt_min_depth_4_plus_5_out),
    .right(index_lt_min_depth_4_plus_5_right)
);
std_and # (
    .WIDTH(1)
) idx_between_5_min_depth_4_plus_5_comb (
    .left(idx_between_5_min_depth_4_plus_5_comb_left),
    .out(idx_between_5_min_depth_4_plus_5_comb_out),
    .right(idx_between_5_min_depth_4_plus_5_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_14_min_depth_4_plus_14_reg (
    .clk(idx_between_14_min_depth_4_plus_14_reg_clk),
    .done(idx_between_14_min_depth_4_plus_14_reg_done),
    .in(idx_between_14_min_depth_4_plus_14_reg_in),
    .out(idx_between_14_min_depth_4_plus_14_reg_out),
    .reset(idx_between_14_min_depth_4_plus_14_reg_reset),
    .write_en(idx_between_14_min_depth_4_plus_14_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_14 (
    .left(index_lt_min_depth_4_plus_14_left),
    .out(index_lt_min_depth_4_plus_14_out),
    .right(index_lt_min_depth_4_plus_14_right)
);
std_and # (
    .WIDTH(1)
) idx_between_14_min_depth_4_plus_14_comb (
    .left(idx_between_14_min_depth_4_plus_14_comb_left),
    .out(idx_between_14_min_depth_4_plus_14_comb_out),
    .right(idx_between_14_min_depth_4_plus_14_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_0_depth_plus_0_reg (
    .clk(idx_between_0_depth_plus_0_reg_clk),
    .done(idx_between_0_depth_plus_0_reg_done),
    .in(idx_between_0_depth_plus_0_reg_in),
    .out(idx_between_0_depth_plus_0_reg_out),
    .reset(idx_between_0_depth_plus_0_reg_reset),
    .write_en(idx_between_0_depth_plus_0_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_0 (
    .left(index_lt_depth_plus_0_left),
    .out(index_lt_depth_plus_0_out),
    .right(index_lt_depth_plus_0_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_9_depth_plus_9_reg (
    .clk(idx_between_9_depth_plus_9_reg_clk),
    .done(idx_between_9_depth_plus_9_reg_done),
    .in(idx_between_9_depth_plus_9_reg_in),
    .out(idx_between_9_depth_plus_9_reg_out),
    .reset(idx_between_9_depth_plus_9_reg_reset),
    .write_en(idx_between_9_depth_plus_9_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_9 (
    .left(index_ge_9_left),
    .out(index_ge_9_out),
    .right(index_ge_9_right)
);
std_and # (
    .WIDTH(1)
) idx_between_9_depth_plus_9_comb (
    .left(idx_between_9_depth_plus_9_comb_left),
    .out(idx_between_9_depth_plus_9_comb_out),
    .right(idx_between_9_depth_plus_9_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_9_min_depth_4_plus_9_reg (
    .clk(idx_between_9_min_depth_4_plus_9_reg_clk),
    .done(idx_between_9_min_depth_4_plus_9_reg_done),
    .in(idx_between_9_min_depth_4_plus_9_reg_in),
    .out(idx_between_9_min_depth_4_plus_9_reg_out),
    .reset(idx_between_9_min_depth_4_plus_9_reg_reset),
    .write_en(idx_between_9_min_depth_4_plus_9_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_9 (
    .left(index_lt_min_depth_4_plus_9_left),
    .out(index_lt_min_depth_4_plus_9_out),
    .right(index_lt_min_depth_4_plus_9_right)
);
std_and # (
    .WIDTH(1)
) idx_between_9_min_depth_4_plus_9_comb (
    .left(idx_between_9_min_depth_4_plus_9_comb_left),
    .out(idx_between_9_min_depth_4_plus_9_comb_out),
    .right(idx_between_9_min_depth_4_plus_9_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_1_depth_plus_1_reg (
    .clk(idx_between_1_depth_plus_1_reg_clk),
    .done(idx_between_1_depth_plus_1_reg_done),
    .in(idx_between_1_depth_plus_1_reg_in),
    .out(idx_between_1_depth_plus_1_reg_out),
    .reset(idx_between_1_depth_plus_1_reg_reset),
    .write_en(idx_between_1_depth_plus_1_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_1 (
    .left(index_lt_depth_plus_1_left),
    .out(index_lt_depth_plus_1_out),
    .right(index_lt_depth_plus_1_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_1 (
    .left(index_ge_1_left),
    .out(index_ge_1_out),
    .right(index_ge_1_right)
);
std_and # (
    .WIDTH(1)
) idx_between_1_depth_plus_1_comb (
    .left(idx_between_1_depth_plus_1_comb_left),
    .out(idx_between_1_depth_plus_1_comb_out),
    .right(idx_between_1_depth_plus_1_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_1_min_depth_4_plus_1_reg (
    .clk(idx_between_1_min_depth_4_plus_1_reg_clk),
    .done(idx_between_1_min_depth_4_plus_1_reg_done),
    .in(idx_between_1_min_depth_4_plus_1_reg_in),
    .out(idx_between_1_min_depth_4_plus_1_reg_out),
    .reset(idx_between_1_min_depth_4_plus_1_reg_reset),
    .write_en(idx_between_1_min_depth_4_plus_1_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_1 (
    .left(index_lt_min_depth_4_plus_1_left),
    .out(index_lt_min_depth_4_plus_1_out),
    .right(index_lt_min_depth_4_plus_1_right)
);
std_and # (
    .WIDTH(1)
) idx_between_1_min_depth_4_plus_1_comb (
    .left(idx_between_1_min_depth_4_plus_1_comb_left),
    .out(idx_between_1_min_depth_4_plus_1_comb_out),
    .right(idx_between_1_min_depth_4_plus_1_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_11_depth_plus_12_reg (
    .clk(idx_between_depth_plus_11_depth_plus_12_reg_clk),
    .done(idx_between_depth_plus_11_depth_plus_12_reg_done),
    .in(idx_between_depth_plus_11_depth_plus_12_reg_in),
    .out(idx_between_depth_plus_11_depth_plus_12_reg_out),
    .reset(idx_between_depth_plus_11_depth_plus_12_reg_reset),
    .write_en(idx_between_depth_plus_11_depth_plus_12_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_11 (
    .left(index_ge_depth_plus_11_left),
    .out(index_ge_depth_plus_11_out),
    .right(index_ge_depth_plus_11_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_11_depth_plus_12_comb (
    .left(idx_between_depth_plus_11_depth_plus_12_comb_left),
    .out(idx_between_depth_plus_11_depth_plus_12_comb_out),
    .right(idx_between_depth_plus_11_depth_plus_12_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_10_depth_plus_10_reg (
    .clk(idx_between_10_depth_plus_10_reg_clk),
    .done(idx_between_10_depth_plus_10_reg_done),
    .in(idx_between_10_depth_plus_10_reg_in),
    .out(idx_between_10_depth_plus_10_reg_out),
    .reset(idx_between_10_depth_plus_10_reg_reset),
    .write_en(idx_between_10_depth_plus_10_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_10 (
    .left(index_ge_10_left),
    .out(index_ge_10_out),
    .right(index_ge_10_right)
);
std_and # (
    .WIDTH(1)
) idx_between_10_depth_plus_10_comb (
    .left(idx_between_10_depth_plus_10_comb_left),
    .out(idx_between_10_depth_plus_10_comb_out),
    .right(idx_between_10_depth_plus_10_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_10_min_depth_4_plus_10_reg (
    .clk(idx_between_10_min_depth_4_plus_10_reg_clk),
    .done(idx_between_10_min_depth_4_plus_10_reg_done),
    .in(idx_between_10_min_depth_4_plus_10_reg_in),
    .out(idx_between_10_min_depth_4_plus_10_reg_out),
    .reset(idx_between_10_min_depth_4_plus_10_reg_reset),
    .write_en(idx_between_10_min_depth_4_plus_10_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_10 (
    .left(index_lt_min_depth_4_plus_10_left),
    .out(index_lt_min_depth_4_plus_10_out),
    .right(index_lt_min_depth_4_plus_10_right)
);
std_and # (
    .WIDTH(1)
) idx_between_10_min_depth_4_plus_10_comb (
    .left(idx_between_10_min_depth_4_plus_10_comb_left),
    .out(idx_between_10_min_depth_4_plus_10_comb_out),
    .right(idx_between_10_min_depth_4_plus_10_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_19_depth_plus_19_reg (
    .clk(idx_between_19_depth_plus_19_reg_clk),
    .done(idx_between_19_depth_plus_19_reg_done),
    .in(idx_between_19_depth_plus_19_reg_in),
    .out(idx_between_19_depth_plus_19_reg_out),
    .reset(idx_between_19_depth_plus_19_reg_reset),
    .write_en(idx_between_19_depth_plus_19_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_19 (
    .left(index_ge_19_left),
    .out(index_ge_19_out),
    .right(index_ge_19_right)
);
std_and # (
    .WIDTH(1)
) idx_between_19_depth_plus_19_comb (
    .left(idx_between_19_depth_plus_19_comb_left),
    .out(idx_between_19_depth_plus_19_comb_out),
    .right(idx_between_19_depth_plus_19_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_6_depth_plus_6_reg (
    .clk(idx_between_6_depth_plus_6_reg_clk),
    .done(idx_between_6_depth_plus_6_reg_done),
    .in(idx_between_6_depth_plus_6_reg_in),
    .out(idx_between_6_depth_plus_6_reg_out),
    .reset(idx_between_6_depth_plus_6_reg_reset),
    .write_en(idx_between_6_depth_plus_6_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_6_depth_plus_6_comb (
    .left(idx_between_6_depth_plus_6_comb_left),
    .out(idx_between_6_depth_plus_6_comb_out),
    .right(idx_between_6_depth_plus_6_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_7_depth_plus_8_reg (
    .clk(idx_between_depth_plus_7_depth_plus_8_reg_clk),
    .done(idx_between_depth_plus_7_depth_plus_8_reg_done),
    .in(idx_between_depth_plus_7_depth_plus_8_reg_in),
    .out(idx_between_depth_plus_7_depth_plus_8_reg_out),
    .reset(idx_between_depth_plus_7_depth_plus_8_reg_reset),
    .write_en(idx_between_depth_plus_7_depth_plus_8_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_7 (
    .left(index_ge_depth_plus_7_left),
    .out(index_ge_depth_plus_7_out),
    .right(index_ge_depth_plus_7_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_7_depth_plus_8_comb (
    .left(idx_between_depth_plus_7_depth_plus_8_comb_left),
    .out(idx_between_depth_plus_7_depth_plus_8_comb_out),
    .right(idx_between_depth_plus_7_depth_plus_8_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_15_min_depth_4_plus_15_reg (
    .clk(idx_between_15_min_depth_4_plus_15_reg_clk),
    .done(idx_between_15_min_depth_4_plus_15_reg_done),
    .in(idx_between_15_min_depth_4_plus_15_reg_in),
    .out(idx_between_15_min_depth_4_plus_15_reg_out),
    .reset(idx_between_15_min_depth_4_plus_15_reg_reset),
    .write_en(idx_between_15_min_depth_4_plus_15_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_15 (
    .left(index_lt_min_depth_4_plus_15_left),
    .out(index_lt_min_depth_4_plus_15_out),
    .right(index_lt_min_depth_4_plus_15_right)
);
std_and # (
    .WIDTH(1)
) idx_between_15_min_depth_4_plus_15_comb (
    .left(idx_between_15_min_depth_4_plus_15_comb_left),
    .out(idx_between_15_min_depth_4_plus_15_comb_out),
    .right(idx_between_15_min_depth_4_plus_15_comb_right)
);
std_reg # (
    .WIDTH(1)
) cond (
    .clk(cond_clk),
    .done(cond_done),
    .in(cond_in),
    .out(cond_out),
    .reset(cond_reset),
    .write_en(cond_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire (
    .in(cond_wire_in),
    .out(cond_wire_out)
);
std_reg # (
    .WIDTH(1)
) cond0 (
    .clk(cond0_clk),
    .done(cond0_done),
    .in(cond0_in),
    .out(cond0_out),
    .reset(cond0_reset),
    .write_en(cond0_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire0 (
    .in(cond_wire0_in),
    .out(cond_wire0_out)
);
std_reg # (
    .WIDTH(1)
) cond1 (
    .clk(cond1_clk),
    .done(cond1_done),
    .in(cond1_in),
    .out(cond1_out),
    .reset(cond1_reset),
    .write_en(cond1_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1 (
    .in(cond_wire1_in),
    .out(cond_wire1_out)
);
std_reg # (
    .WIDTH(1)
) cond2 (
    .clk(cond2_clk),
    .done(cond2_done),
    .in(cond2_in),
    .out(cond2_out),
    .reset(cond2_reset),
    .write_en(cond2_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire2 (
    .in(cond_wire2_in),
    .out(cond_wire2_out)
);
std_reg # (
    .WIDTH(1)
) cond3 (
    .clk(cond3_clk),
    .done(cond3_done),
    .in(cond3_in),
    .out(cond3_out),
    .reset(cond3_reset),
    .write_en(cond3_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire3 (
    .in(cond_wire3_in),
    .out(cond_wire3_out)
);
std_reg # (
    .WIDTH(1)
) cond4 (
    .clk(cond4_clk),
    .done(cond4_done),
    .in(cond4_in),
    .out(cond4_out),
    .reset(cond4_reset),
    .write_en(cond4_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire4 (
    .in(cond_wire4_in),
    .out(cond_wire4_out)
);
std_reg # (
    .WIDTH(1)
) cond5 (
    .clk(cond5_clk),
    .done(cond5_done),
    .in(cond5_in),
    .out(cond5_out),
    .reset(cond5_reset),
    .write_en(cond5_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire5 (
    .in(cond_wire5_in),
    .out(cond_wire5_out)
);
std_reg # (
    .WIDTH(1)
) cond6 (
    .clk(cond6_clk),
    .done(cond6_done),
    .in(cond6_in),
    .out(cond6_out),
    .reset(cond6_reset),
    .write_en(cond6_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire6 (
    .in(cond_wire6_in),
    .out(cond_wire6_out)
);
std_reg # (
    .WIDTH(1)
) cond7 (
    .clk(cond7_clk),
    .done(cond7_done),
    .in(cond7_in),
    .out(cond7_out),
    .reset(cond7_reset),
    .write_en(cond7_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire7 (
    .in(cond_wire7_in),
    .out(cond_wire7_out)
);
std_reg # (
    .WIDTH(1)
) cond8 (
    .clk(cond8_clk),
    .done(cond8_done),
    .in(cond8_in),
    .out(cond8_out),
    .reset(cond8_reset),
    .write_en(cond8_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire8 (
    .in(cond_wire8_in),
    .out(cond_wire8_out)
);
std_reg # (
    .WIDTH(1)
) cond9 (
    .clk(cond9_clk),
    .done(cond9_done),
    .in(cond9_in),
    .out(cond9_out),
    .reset(cond9_reset),
    .write_en(cond9_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire9 (
    .in(cond_wire9_in),
    .out(cond_wire9_out)
);
std_reg # (
    .WIDTH(1)
) cond10 (
    .clk(cond10_clk),
    .done(cond10_done),
    .in(cond10_in),
    .out(cond10_out),
    .reset(cond10_reset),
    .write_en(cond10_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire10 (
    .in(cond_wire10_in),
    .out(cond_wire10_out)
);
std_reg # (
    .WIDTH(1)
) cond11 (
    .clk(cond11_clk),
    .done(cond11_done),
    .in(cond11_in),
    .out(cond11_out),
    .reset(cond11_reset),
    .write_en(cond11_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire11 (
    .in(cond_wire11_in),
    .out(cond_wire11_out)
);
std_reg # (
    .WIDTH(1)
) cond12 (
    .clk(cond12_clk),
    .done(cond12_done),
    .in(cond12_in),
    .out(cond12_out),
    .reset(cond12_reset),
    .write_en(cond12_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire12 (
    .in(cond_wire12_in),
    .out(cond_wire12_out)
);
std_reg # (
    .WIDTH(1)
) cond13 (
    .clk(cond13_clk),
    .done(cond13_done),
    .in(cond13_in),
    .out(cond13_out),
    .reset(cond13_reset),
    .write_en(cond13_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire13 (
    .in(cond_wire13_in),
    .out(cond_wire13_out)
);
std_reg # (
    .WIDTH(1)
) cond14 (
    .clk(cond14_clk),
    .done(cond14_done),
    .in(cond14_in),
    .out(cond14_out),
    .reset(cond14_reset),
    .write_en(cond14_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire14 (
    .in(cond_wire14_in),
    .out(cond_wire14_out)
);
std_reg # (
    .WIDTH(1)
) cond15 (
    .clk(cond15_clk),
    .done(cond15_done),
    .in(cond15_in),
    .out(cond15_out),
    .reset(cond15_reset),
    .write_en(cond15_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire15 (
    .in(cond_wire15_in),
    .out(cond_wire15_out)
);
std_reg # (
    .WIDTH(1)
) cond16 (
    .clk(cond16_clk),
    .done(cond16_done),
    .in(cond16_in),
    .out(cond16_out),
    .reset(cond16_reset),
    .write_en(cond16_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire16 (
    .in(cond_wire16_in),
    .out(cond_wire16_out)
);
std_reg # (
    .WIDTH(1)
) cond17 (
    .clk(cond17_clk),
    .done(cond17_done),
    .in(cond17_in),
    .out(cond17_out),
    .reset(cond17_reset),
    .write_en(cond17_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire17 (
    .in(cond_wire17_in),
    .out(cond_wire17_out)
);
std_reg # (
    .WIDTH(1)
) cond18 (
    .clk(cond18_clk),
    .done(cond18_done),
    .in(cond18_in),
    .out(cond18_out),
    .reset(cond18_reset),
    .write_en(cond18_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire18 (
    .in(cond_wire18_in),
    .out(cond_wire18_out)
);
std_reg # (
    .WIDTH(1)
) cond19 (
    .clk(cond19_clk),
    .done(cond19_done),
    .in(cond19_in),
    .out(cond19_out),
    .reset(cond19_reset),
    .write_en(cond19_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire19 (
    .in(cond_wire19_in),
    .out(cond_wire19_out)
);
std_reg # (
    .WIDTH(1)
) cond20 (
    .clk(cond20_clk),
    .done(cond20_done),
    .in(cond20_in),
    .out(cond20_out),
    .reset(cond20_reset),
    .write_en(cond20_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire20 (
    .in(cond_wire20_in),
    .out(cond_wire20_out)
);
std_reg # (
    .WIDTH(1)
) cond21 (
    .clk(cond21_clk),
    .done(cond21_done),
    .in(cond21_in),
    .out(cond21_out),
    .reset(cond21_reset),
    .write_en(cond21_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire21 (
    .in(cond_wire21_in),
    .out(cond_wire21_out)
);
std_reg # (
    .WIDTH(1)
) cond22 (
    .clk(cond22_clk),
    .done(cond22_done),
    .in(cond22_in),
    .out(cond22_out),
    .reset(cond22_reset),
    .write_en(cond22_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire22 (
    .in(cond_wire22_in),
    .out(cond_wire22_out)
);
std_reg # (
    .WIDTH(1)
) cond23 (
    .clk(cond23_clk),
    .done(cond23_done),
    .in(cond23_in),
    .out(cond23_out),
    .reset(cond23_reset),
    .write_en(cond23_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire23 (
    .in(cond_wire23_in),
    .out(cond_wire23_out)
);
std_reg # (
    .WIDTH(1)
) cond24 (
    .clk(cond24_clk),
    .done(cond24_done),
    .in(cond24_in),
    .out(cond24_out),
    .reset(cond24_reset),
    .write_en(cond24_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire24 (
    .in(cond_wire24_in),
    .out(cond_wire24_out)
);
std_reg # (
    .WIDTH(1)
) cond25 (
    .clk(cond25_clk),
    .done(cond25_done),
    .in(cond25_in),
    .out(cond25_out),
    .reset(cond25_reset),
    .write_en(cond25_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire25 (
    .in(cond_wire25_in),
    .out(cond_wire25_out)
);
std_reg # (
    .WIDTH(1)
) cond26 (
    .clk(cond26_clk),
    .done(cond26_done),
    .in(cond26_in),
    .out(cond26_out),
    .reset(cond26_reset),
    .write_en(cond26_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire26 (
    .in(cond_wire26_in),
    .out(cond_wire26_out)
);
std_reg # (
    .WIDTH(1)
) cond27 (
    .clk(cond27_clk),
    .done(cond27_done),
    .in(cond27_in),
    .out(cond27_out),
    .reset(cond27_reset),
    .write_en(cond27_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire27 (
    .in(cond_wire27_in),
    .out(cond_wire27_out)
);
std_reg # (
    .WIDTH(1)
) cond28 (
    .clk(cond28_clk),
    .done(cond28_done),
    .in(cond28_in),
    .out(cond28_out),
    .reset(cond28_reset),
    .write_en(cond28_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire28 (
    .in(cond_wire28_in),
    .out(cond_wire28_out)
);
std_reg # (
    .WIDTH(1)
) cond29 (
    .clk(cond29_clk),
    .done(cond29_done),
    .in(cond29_in),
    .out(cond29_out),
    .reset(cond29_reset),
    .write_en(cond29_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire29 (
    .in(cond_wire29_in),
    .out(cond_wire29_out)
);
std_reg # (
    .WIDTH(1)
) cond30 (
    .clk(cond30_clk),
    .done(cond30_done),
    .in(cond30_in),
    .out(cond30_out),
    .reset(cond30_reset),
    .write_en(cond30_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire30 (
    .in(cond_wire30_in),
    .out(cond_wire30_out)
);
std_reg # (
    .WIDTH(1)
) cond31 (
    .clk(cond31_clk),
    .done(cond31_done),
    .in(cond31_in),
    .out(cond31_out),
    .reset(cond31_reset),
    .write_en(cond31_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire31 (
    .in(cond_wire31_in),
    .out(cond_wire31_out)
);
std_reg # (
    .WIDTH(1)
) cond32 (
    .clk(cond32_clk),
    .done(cond32_done),
    .in(cond32_in),
    .out(cond32_out),
    .reset(cond32_reset),
    .write_en(cond32_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire32 (
    .in(cond_wire32_in),
    .out(cond_wire32_out)
);
std_reg # (
    .WIDTH(1)
) cond33 (
    .clk(cond33_clk),
    .done(cond33_done),
    .in(cond33_in),
    .out(cond33_out),
    .reset(cond33_reset),
    .write_en(cond33_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire33 (
    .in(cond_wire33_in),
    .out(cond_wire33_out)
);
std_reg # (
    .WIDTH(1)
) cond34 (
    .clk(cond34_clk),
    .done(cond34_done),
    .in(cond34_in),
    .out(cond34_out),
    .reset(cond34_reset),
    .write_en(cond34_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire34 (
    .in(cond_wire34_in),
    .out(cond_wire34_out)
);
std_reg # (
    .WIDTH(1)
) cond35 (
    .clk(cond35_clk),
    .done(cond35_done),
    .in(cond35_in),
    .out(cond35_out),
    .reset(cond35_reset),
    .write_en(cond35_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire35 (
    .in(cond_wire35_in),
    .out(cond_wire35_out)
);
std_reg # (
    .WIDTH(1)
) cond36 (
    .clk(cond36_clk),
    .done(cond36_done),
    .in(cond36_in),
    .out(cond36_out),
    .reset(cond36_reset),
    .write_en(cond36_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire36 (
    .in(cond_wire36_in),
    .out(cond_wire36_out)
);
std_reg # (
    .WIDTH(1)
) cond37 (
    .clk(cond37_clk),
    .done(cond37_done),
    .in(cond37_in),
    .out(cond37_out),
    .reset(cond37_reset),
    .write_en(cond37_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire37 (
    .in(cond_wire37_in),
    .out(cond_wire37_out)
);
std_reg # (
    .WIDTH(1)
) cond38 (
    .clk(cond38_clk),
    .done(cond38_done),
    .in(cond38_in),
    .out(cond38_out),
    .reset(cond38_reset),
    .write_en(cond38_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire38 (
    .in(cond_wire38_in),
    .out(cond_wire38_out)
);
std_reg # (
    .WIDTH(1)
) cond39 (
    .clk(cond39_clk),
    .done(cond39_done),
    .in(cond39_in),
    .out(cond39_out),
    .reset(cond39_reset),
    .write_en(cond39_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire39 (
    .in(cond_wire39_in),
    .out(cond_wire39_out)
);
std_reg # (
    .WIDTH(1)
) cond40 (
    .clk(cond40_clk),
    .done(cond40_done),
    .in(cond40_in),
    .out(cond40_out),
    .reset(cond40_reset),
    .write_en(cond40_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire40 (
    .in(cond_wire40_in),
    .out(cond_wire40_out)
);
std_reg # (
    .WIDTH(1)
) cond41 (
    .clk(cond41_clk),
    .done(cond41_done),
    .in(cond41_in),
    .out(cond41_out),
    .reset(cond41_reset),
    .write_en(cond41_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire41 (
    .in(cond_wire41_in),
    .out(cond_wire41_out)
);
std_reg # (
    .WIDTH(1)
) cond42 (
    .clk(cond42_clk),
    .done(cond42_done),
    .in(cond42_in),
    .out(cond42_out),
    .reset(cond42_reset),
    .write_en(cond42_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire42 (
    .in(cond_wire42_in),
    .out(cond_wire42_out)
);
std_reg # (
    .WIDTH(1)
) cond43 (
    .clk(cond43_clk),
    .done(cond43_done),
    .in(cond43_in),
    .out(cond43_out),
    .reset(cond43_reset),
    .write_en(cond43_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire43 (
    .in(cond_wire43_in),
    .out(cond_wire43_out)
);
std_reg # (
    .WIDTH(1)
) cond44 (
    .clk(cond44_clk),
    .done(cond44_done),
    .in(cond44_in),
    .out(cond44_out),
    .reset(cond44_reset),
    .write_en(cond44_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire44 (
    .in(cond_wire44_in),
    .out(cond_wire44_out)
);
std_reg # (
    .WIDTH(1)
) cond45 (
    .clk(cond45_clk),
    .done(cond45_done),
    .in(cond45_in),
    .out(cond45_out),
    .reset(cond45_reset),
    .write_en(cond45_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire45 (
    .in(cond_wire45_in),
    .out(cond_wire45_out)
);
std_reg # (
    .WIDTH(1)
) cond46 (
    .clk(cond46_clk),
    .done(cond46_done),
    .in(cond46_in),
    .out(cond46_out),
    .reset(cond46_reset),
    .write_en(cond46_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire46 (
    .in(cond_wire46_in),
    .out(cond_wire46_out)
);
std_reg # (
    .WIDTH(1)
) cond47 (
    .clk(cond47_clk),
    .done(cond47_done),
    .in(cond47_in),
    .out(cond47_out),
    .reset(cond47_reset),
    .write_en(cond47_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire47 (
    .in(cond_wire47_in),
    .out(cond_wire47_out)
);
std_reg # (
    .WIDTH(1)
) cond48 (
    .clk(cond48_clk),
    .done(cond48_done),
    .in(cond48_in),
    .out(cond48_out),
    .reset(cond48_reset),
    .write_en(cond48_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire48 (
    .in(cond_wire48_in),
    .out(cond_wire48_out)
);
std_reg # (
    .WIDTH(1)
) cond49 (
    .clk(cond49_clk),
    .done(cond49_done),
    .in(cond49_in),
    .out(cond49_out),
    .reset(cond49_reset),
    .write_en(cond49_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire49 (
    .in(cond_wire49_in),
    .out(cond_wire49_out)
);
std_reg # (
    .WIDTH(1)
) cond50 (
    .clk(cond50_clk),
    .done(cond50_done),
    .in(cond50_in),
    .out(cond50_out),
    .reset(cond50_reset),
    .write_en(cond50_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire50 (
    .in(cond_wire50_in),
    .out(cond_wire50_out)
);
std_reg # (
    .WIDTH(1)
) cond51 (
    .clk(cond51_clk),
    .done(cond51_done),
    .in(cond51_in),
    .out(cond51_out),
    .reset(cond51_reset),
    .write_en(cond51_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire51 (
    .in(cond_wire51_in),
    .out(cond_wire51_out)
);
std_reg # (
    .WIDTH(1)
) cond52 (
    .clk(cond52_clk),
    .done(cond52_done),
    .in(cond52_in),
    .out(cond52_out),
    .reset(cond52_reset),
    .write_en(cond52_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire52 (
    .in(cond_wire52_in),
    .out(cond_wire52_out)
);
std_reg # (
    .WIDTH(1)
) cond53 (
    .clk(cond53_clk),
    .done(cond53_done),
    .in(cond53_in),
    .out(cond53_out),
    .reset(cond53_reset),
    .write_en(cond53_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire53 (
    .in(cond_wire53_in),
    .out(cond_wire53_out)
);
std_reg # (
    .WIDTH(1)
) cond54 (
    .clk(cond54_clk),
    .done(cond54_done),
    .in(cond54_in),
    .out(cond54_out),
    .reset(cond54_reset),
    .write_en(cond54_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire54 (
    .in(cond_wire54_in),
    .out(cond_wire54_out)
);
std_reg # (
    .WIDTH(1)
) cond55 (
    .clk(cond55_clk),
    .done(cond55_done),
    .in(cond55_in),
    .out(cond55_out),
    .reset(cond55_reset),
    .write_en(cond55_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire55 (
    .in(cond_wire55_in),
    .out(cond_wire55_out)
);
std_reg # (
    .WIDTH(1)
) cond56 (
    .clk(cond56_clk),
    .done(cond56_done),
    .in(cond56_in),
    .out(cond56_out),
    .reset(cond56_reset),
    .write_en(cond56_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire56 (
    .in(cond_wire56_in),
    .out(cond_wire56_out)
);
std_reg # (
    .WIDTH(1)
) cond57 (
    .clk(cond57_clk),
    .done(cond57_done),
    .in(cond57_in),
    .out(cond57_out),
    .reset(cond57_reset),
    .write_en(cond57_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire57 (
    .in(cond_wire57_in),
    .out(cond_wire57_out)
);
std_reg # (
    .WIDTH(1)
) cond58 (
    .clk(cond58_clk),
    .done(cond58_done),
    .in(cond58_in),
    .out(cond58_out),
    .reset(cond58_reset),
    .write_en(cond58_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire58 (
    .in(cond_wire58_in),
    .out(cond_wire58_out)
);
std_reg # (
    .WIDTH(1)
) cond59 (
    .clk(cond59_clk),
    .done(cond59_done),
    .in(cond59_in),
    .out(cond59_out),
    .reset(cond59_reset),
    .write_en(cond59_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire59 (
    .in(cond_wire59_in),
    .out(cond_wire59_out)
);
std_reg # (
    .WIDTH(1)
) cond60 (
    .clk(cond60_clk),
    .done(cond60_done),
    .in(cond60_in),
    .out(cond60_out),
    .reset(cond60_reset),
    .write_en(cond60_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire60 (
    .in(cond_wire60_in),
    .out(cond_wire60_out)
);
std_reg # (
    .WIDTH(1)
) cond61 (
    .clk(cond61_clk),
    .done(cond61_done),
    .in(cond61_in),
    .out(cond61_out),
    .reset(cond61_reset),
    .write_en(cond61_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire61 (
    .in(cond_wire61_in),
    .out(cond_wire61_out)
);
std_reg # (
    .WIDTH(1)
) cond62 (
    .clk(cond62_clk),
    .done(cond62_done),
    .in(cond62_in),
    .out(cond62_out),
    .reset(cond62_reset),
    .write_en(cond62_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire62 (
    .in(cond_wire62_in),
    .out(cond_wire62_out)
);
std_reg # (
    .WIDTH(1)
) cond63 (
    .clk(cond63_clk),
    .done(cond63_done),
    .in(cond63_in),
    .out(cond63_out),
    .reset(cond63_reset),
    .write_en(cond63_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire63 (
    .in(cond_wire63_in),
    .out(cond_wire63_out)
);
std_reg # (
    .WIDTH(1)
) cond64 (
    .clk(cond64_clk),
    .done(cond64_done),
    .in(cond64_in),
    .out(cond64_out),
    .reset(cond64_reset),
    .write_en(cond64_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire64 (
    .in(cond_wire64_in),
    .out(cond_wire64_out)
);
std_reg # (
    .WIDTH(1)
) cond65 (
    .clk(cond65_clk),
    .done(cond65_done),
    .in(cond65_in),
    .out(cond65_out),
    .reset(cond65_reset),
    .write_en(cond65_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire65 (
    .in(cond_wire65_in),
    .out(cond_wire65_out)
);
std_reg # (
    .WIDTH(1)
) cond66 (
    .clk(cond66_clk),
    .done(cond66_done),
    .in(cond66_in),
    .out(cond66_out),
    .reset(cond66_reset),
    .write_en(cond66_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire66 (
    .in(cond_wire66_in),
    .out(cond_wire66_out)
);
std_reg # (
    .WIDTH(1)
) cond67 (
    .clk(cond67_clk),
    .done(cond67_done),
    .in(cond67_in),
    .out(cond67_out),
    .reset(cond67_reset),
    .write_en(cond67_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire67 (
    .in(cond_wire67_in),
    .out(cond_wire67_out)
);
std_reg # (
    .WIDTH(1)
) cond68 (
    .clk(cond68_clk),
    .done(cond68_done),
    .in(cond68_in),
    .out(cond68_out),
    .reset(cond68_reset),
    .write_en(cond68_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire68 (
    .in(cond_wire68_in),
    .out(cond_wire68_out)
);
std_reg # (
    .WIDTH(1)
) cond69 (
    .clk(cond69_clk),
    .done(cond69_done),
    .in(cond69_in),
    .out(cond69_out),
    .reset(cond69_reset),
    .write_en(cond69_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire69 (
    .in(cond_wire69_in),
    .out(cond_wire69_out)
);
std_reg # (
    .WIDTH(1)
) cond70 (
    .clk(cond70_clk),
    .done(cond70_done),
    .in(cond70_in),
    .out(cond70_out),
    .reset(cond70_reset),
    .write_en(cond70_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire70 (
    .in(cond_wire70_in),
    .out(cond_wire70_out)
);
std_reg # (
    .WIDTH(1)
) cond71 (
    .clk(cond71_clk),
    .done(cond71_done),
    .in(cond71_in),
    .out(cond71_out),
    .reset(cond71_reset),
    .write_en(cond71_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire71 (
    .in(cond_wire71_in),
    .out(cond_wire71_out)
);
std_reg # (
    .WIDTH(1)
) cond72 (
    .clk(cond72_clk),
    .done(cond72_done),
    .in(cond72_in),
    .out(cond72_out),
    .reset(cond72_reset),
    .write_en(cond72_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire72 (
    .in(cond_wire72_in),
    .out(cond_wire72_out)
);
std_reg # (
    .WIDTH(1)
) cond73 (
    .clk(cond73_clk),
    .done(cond73_done),
    .in(cond73_in),
    .out(cond73_out),
    .reset(cond73_reset),
    .write_en(cond73_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire73 (
    .in(cond_wire73_in),
    .out(cond_wire73_out)
);
std_reg # (
    .WIDTH(1)
) cond74 (
    .clk(cond74_clk),
    .done(cond74_done),
    .in(cond74_in),
    .out(cond74_out),
    .reset(cond74_reset),
    .write_en(cond74_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire74 (
    .in(cond_wire74_in),
    .out(cond_wire74_out)
);
std_reg # (
    .WIDTH(1)
) cond75 (
    .clk(cond75_clk),
    .done(cond75_done),
    .in(cond75_in),
    .out(cond75_out),
    .reset(cond75_reset),
    .write_en(cond75_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire75 (
    .in(cond_wire75_in),
    .out(cond_wire75_out)
);
std_reg # (
    .WIDTH(1)
) cond76 (
    .clk(cond76_clk),
    .done(cond76_done),
    .in(cond76_in),
    .out(cond76_out),
    .reset(cond76_reset),
    .write_en(cond76_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire76 (
    .in(cond_wire76_in),
    .out(cond_wire76_out)
);
std_reg # (
    .WIDTH(1)
) cond77 (
    .clk(cond77_clk),
    .done(cond77_done),
    .in(cond77_in),
    .out(cond77_out),
    .reset(cond77_reset),
    .write_en(cond77_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire77 (
    .in(cond_wire77_in),
    .out(cond_wire77_out)
);
std_reg # (
    .WIDTH(1)
) cond78 (
    .clk(cond78_clk),
    .done(cond78_done),
    .in(cond78_in),
    .out(cond78_out),
    .reset(cond78_reset),
    .write_en(cond78_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire78 (
    .in(cond_wire78_in),
    .out(cond_wire78_out)
);
std_reg # (
    .WIDTH(1)
) cond79 (
    .clk(cond79_clk),
    .done(cond79_done),
    .in(cond79_in),
    .out(cond79_out),
    .reset(cond79_reset),
    .write_en(cond79_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire79 (
    .in(cond_wire79_in),
    .out(cond_wire79_out)
);
std_reg # (
    .WIDTH(1)
) cond80 (
    .clk(cond80_clk),
    .done(cond80_done),
    .in(cond80_in),
    .out(cond80_out),
    .reset(cond80_reset),
    .write_en(cond80_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire80 (
    .in(cond_wire80_in),
    .out(cond_wire80_out)
);
std_reg # (
    .WIDTH(1)
) cond81 (
    .clk(cond81_clk),
    .done(cond81_done),
    .in(cond81_in),
    .out(cond81_out),
    .reset(cond81_reset),
    .write_en(cond81_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire81 (
    .in(cond_wire81_in),
    .out(cond_wire81_out)
);
std_reg # (
    .WIDTH(1)
) cond82 (
    .clk(cond82_clk),
    .done(cond82_done),
    .in(cond82_in),
    .out(cond82_out),
    .reset(cond82_reset),
    .write_en(cond82_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire82 (
    .in(cond_wire82_in),
    .out(cond_wire82_out)
);
std_reg # (
    .WIDTH(1)
) cond83 (
    .clk(cond83_clk),
    .done(cond83_done),
    .in(cond83_in),
    .out(cond83_out),
    .reset(cond83_reset),
    .write_en(cond83_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire83 (
    .in(cond_wire83_in),
    .out(cond_wire83_out)
);
std_reg # (
    .WIDTH(1)
) cond84 (
    .clk(cond84_clk),
    .done(cond84_done),
    .in(cond84_in),
    .out(cond84_out),
    .reset(cond84_reset),
    .write_en(cond84_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire84 (
    .in(cond_wire84_in),
    .out(cond_wire84_out)
);
std_reg # (
    .WIDTH(1)
) cond85 (
    .clk(cond85_clk),
    .done(cond85_done),
    .in(cond85_in),
    .out(cond85_out),
    .reset(cond85_reset),
    .write_en(cond85_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire85 (
    .in(cond_wire85_in),
    .out(cond_wire85_out)
);
std_reg # (
    .WIDTH(1)
) cond86 (
    .clk(cond86_clk),
    .done(cond86_done),
    .in(cond86_in),
    .out(cond86_out),
    .reset(cond86_reset),
    .write_en(cond86_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire86 (
    .in(cond_wire86_in),
    .out(cond_wire86_out)
);
std_reg # (
    .WIDTH(1)
) cond87 (
    .clk(cond87_clk),
    .done(cond87_done),
    .in(cond87_in),
    .out(cond87_out),
    .reset(cond87_reset),
    .write_en(cond87_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire87 (
    .in(cond_wire87_in),
    .out(cond_wire87_out)
);
std_reg # (
    .WIDTH(1)
) cond88 (
    .clk(cond88_clk),
    .done(cond88_done),
    .in(cond88_in),
    .out(cond88_out),
    .reset(cond88_reset),
    .write_en(cond88_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire88 (
    .in(cond_wire88_in),
    .out(cond_wire88_out)
);
std_reg # (
    .WIDTH(1)
) cond89 (
    .clk(cond89_clk),
    .done(cond89_done),
    .in(cond89_in),
    .out(cond89_out),
    .reset(cond89_reset),
    .write_en(cond89_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire89 (
    .in(cond_wire89_in),
    .out(cond_wire89_out)
);
std_reg # (
    .WIDTH(1)
) cond90 (
    .clk(cond90_clk),
    .done(cond90_done),
    .in(cond90_in),
    .out(cond90_out),
    .reset(cond90_reset),
    .write_en(cond90_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire90 (
    .in(cond_wire90_in),
    .out(cond_wire90_out)
);
std_reg # (
    .WIDTH(1)
) cond91 (
    .clk(cond91_clk),
    .done(cond91_done),
    .in(cond91_in),
    .out(cond91_out),
    .reset(cond91_reset),
    .write_en(cond91_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire91 (
    .in(cond_wire91_in),
    .out(cond_wire91_out)
);
std_reg # (
    .WIDTH(1)
) cond92 (
    .clk(cond92_clk),
    .done(cond92_done),
    .in(cond92_in),
    .out(cond92_out),
    .reset(cond92_reset),
    .write_en(cond92_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire92 (
    .in(cond_wire92_in),
    .out(cond_wire92_out)
);
std_reg # (
    .WIDTH(1)
) cond93 (
    .clk(cond93_clk),
    .done(cond93_done),
    .in(cond93_in),
    .out(cond93_out),
    .reset(cond93_reset),
    .write_en(cond93_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire93 (
    .in(cond_wire93_in),
    .out(cond_wire93_out)
);
std_reg # (
    .WIDTH(1)
) cond94 (
    .clk(cond94_clk),
    .done(cond94_done),
    .in(cond94_in),
    .out(cond94_out),
    .reset(cond94_reset),
    .write_en(cond94_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire94 (
    .in(cond_wire94_in),
    .out(cond_wire94_out)
);
std_reg # (
    .WIDTH(1)
) cond95 (
    .clk(cond95_clk),
    .done(cond95_done),
    .in(cond95_in),
    .out(cond95_out),
    .reset(cond95_reset),
    .write_en(cond95_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire95 (
    .in(cond_wire95_in),
    .out(cond_wire95_out)
);
std_reg # (
    .WIDTH(1)
) cond96 (
    .clk(cond96_clk),
    .done(cond96_done),
    .in(cond96_in),
    .out(cond96_out),
    .reset(cond96_reset),
    .write_en(cond96_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire96 (
    .in(cond_wire96_in),
    .out(cond_wire96_out)
);
std_reg # (
    .WIDTH(1)
) cond97 (
    .clk(cond97_clk),
    .done(cond97_done),
    .in(cond97_in),
    .out(cond97_out),
    .reset(cond97_reset),
    .write_en(cond97_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire97 (
    .in(cond_wire97_in),
    .out(cond_wire97_out)
);
std_reg # (
    .WIDTH(1)
) cond98 (
    .clk(cond98_clk),
    .done(cond98_done),
    .in(cond98_in),
    .out(cond98_out),
    .reset(cond98_reset),
    .write_en(cond98_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire98 (
    .in(cond_wire98_in),
    .out(cond_wire98_out)
);
std_reg # (
    .WIDTH(1)
) cond99 (
    .clk(cond99_clk),
    .done(cond99_done),
    .in(cond99_in),
    .out(cond99_out),
    .reset(cond99_reset),
    .write_en(cond99_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire99 (
    .in(cond_wire99_in),
    .out(cond_wire99_out)
);
std_reg # (
    .WIDTH(1)
) cond100 (
    .clk(cond100_clk),
    .done(cond100_done),
    .in(cond100_in),
    .out(cond100_out),
    .reset(cond100_reset),
    .write_en(cond100_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire100 (
    .in(cond_wire100_in),
    .out(cond_wire100_out)
);
std_reg # (
    .WIDTH(1)
) cond101 (
    .clk(cond101_clk),
    .done(cond101_done),
    .in(cond101_in),
    .out(cond101_out),
    .reset(cond101_reset),
    .write_en(cond101_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire101 (
    .in(cond_wire101_in),
    .out(cond_wire101_out)
);
std_reg # (
    .WIDTH(1)
) cond102 (
    .clk(cond102_clk),
    .done(cond102_done),
    .in(cond102_in),
    .out(cond102_out),
    .reset(cond102_reset),
    .write_en(cond102_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire102 (
    .in(cond_wire102_in),
    .out(cond_wire102_out)
);
std_reg # (
    .WIDTH(1)
) cond103 (
    .clk(cond103_clk),
    .done(cond103_done),
    .in(cond103_in),
    .out(cond103_out),
    .reset(cond103_reset),
    .write_en(cond103_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire103 (
    .in(cond_wire103_in),
    .out(cond_wire103_out)
);
std_reg # (
    .WIDTH(1)
) cond104 (
    .clk(cond104_clk),
    .done(cond104_done),
    .in(cond104_in),
    .out(cond104_out),
    .reset(cond104_reset),
    .write_en(cond104_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire104 (
    .in(cond_wire104_in),
    .out(cond_wire104_out)
);
std_reg # (
    .WIDTH(1)
) cond105 (
    .clk(cond105_clk),
    .done(cond105_done),
    .in(cond105_in),
    .out(cond105_out),
    .reset(cond105_reset),
    .write_en(cond105_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire105 (
    .in(cond_wire105_in),
    .out(cond_wire105_out)
);
std_reg # (
    .WIDTH(1)
) cond106 (
    .clk(cond106_clk),
    .done(cond106_done),
    .in(cond106_in),
    .out(cond106_out),
    .reset(cond106_reset),
    .write_en(cond106_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire106 (
    .in(cond_wire106_in),
    .out(cond_wire106_out)
);
std_reg # (
    .WIDTH(1)
) cond107 (
    .clk(cond107_clk),
    .done(cond107_done),
    .in(cond107_in),
    .out(cond107_out),
    .reset(cond107_reset),
    .write_en(cond107_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire107 (
    .in(cond_wire107_in),
    .out(cond_wire107_out)
);
std_reg # (
    .WIDTH(1)
) cond108 (
    .clk(cond108_clk),
    .done(cond108_done),
    .in(cond108_in),
    .out(cond108_out),
    .reset(cond108_reset),
    .write_en(cond108_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire108 (
    .in(cond_wire108_in),
    .out(cond_wire108_out)
);
std_reg # (
    .WIDTH(1)
) cond109 (
    .clk(cond109_clk),
    .done(cond109_done),
    .in(cond109_in),
    .out(cond109_out),
    .reset(cond109_reset),
    .write_en(cond109_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire109 (
    .in(cond_wire109_in),
    .out(cond_wire109_out)
);
std_reg # (
    .WIDTH(1)
) cond110 (
    .clk(cond110_clk),
    .done(cond110_done),
    .in(cond110_in),
    .out(cond110_out),
    .reset(cond110_reset),
    .write_en(cond110_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire110 (
    .in(cond_wire110_in),
    .out(cond_wire110_out)
);
std_reg # (
    .WIDTH(1)
) cond111 (
    .clk(cond111_clk),
    .done(cond111_done),
    .in(cond111_in),
    .out(cond111_out),
    .reset(cond111_reset),
    .write_en(cond111_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire111 (
    .in(cond_wire111_in),
    .out(cond_wire111_out)
);
std_reg # (
    .WIDTH(1)
) cond112 (
    .clk(cond112_clk),
    .done(cond112_done),
    .in(cond112_in),
    .out(cond112_out),
    .reset(cond112_reset),
    .write_en(cond112_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire112 (
    .in(cond_wire112_in),
    .out(cond_wire112_out)
);
std_reg # (
    .WIDTH(1)
) cond113 (
    .clk(cond113_clk),
    .done(cond113_done),
    .in(cond113_in),
    .out(cond113_out),
    .reset(cond113_reset),
    .write_en(cond113_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire113 (
    .in(cond_wire113_in),
    .out(cond_wire113_out)
);
std_reg # (
    .WIDTH(1)
) cond114 (
    .clk(cond114_clk),
    .done(cond114_done),
    .in(cond114_in),
    .out(cond114_out),
    .reset(cond114_reset),
    .write_en(cond114_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire114 (
    .in(cond_wire114_in),
    .out(cond_wire114_out)
);
std_reg # (
    .WIDTH(1)
) cond115 (
    .clk(cond115_clk),
    .done(cond115_done),
    .in(cond115_in),
    .out(cond115_out),
    .reset(cond115_reset),
    .write_en(cond115_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire115 (
    .in(cond_wire115_in),
    .out(cond_wire115_out)
);
std_reg # (
    .WIDTH(1)
) cond116 (
    .clk(cond116_clk),
    .done(cond116_done),
    .in(cond116_in),
    .out(cond116_out),
    .reset(cond116_reset),
    .write_en(cond116_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire116 (
    .in(cond_wire116_in),
    .out(cond_wire116_out)
);
std_reg # (
    .WIDTH(1)
) cond117 (
    .clk(cond117_clk),
    .done(cond117_done),
    .in(cond117_in),
    .out(cond117_out),
    .reset(cond117_reset),
    .write_en(cond117_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire117 (
    .in(cond_wire117_in),
    .out(cond_wire117_out)
);
std_reg # (
    .WIDTH(1)
) cond118 (
    .clk(cond118_clk),
    .done(cond118_done),
    .in(cond118_in),
    .out(cond118_out),
    .reset(cond118_reset),
    .write_en(cond118_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire118 (
    .in(cond_wire118_in),
    .out(cond_wire118_out)
);
std_reg # (
    .WIDTH(1)
) cond119 (
    .clk(cond119_clk),
    .done(cond119_done),
    .in(cond119_in),
    .out(cond119_out),
    .reset(cond119_reset),
    .write_en(cond119_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire119 (
    .in(cond_wire119_in),
    .out(cond_wire119_out)
);
std_reg # (
    .WIDTH(1)
) cond120 (
    .clk(cond120_clk),
    .done(cond120_done),
    .in(cond120_in),
    .out(cond120_out),
    .reset(cond120_reset),
    .write_en(cond120_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire120 (
    .in(cond_wire120_in),
    .out(cond_wire120_out)
);
std_reg # (
    .WIDTH(1)
) cond121 (
    .clk(cond121_clk),
    .done(cond121_done),
    .in(cond121_in),
    .out(cond121_out),
    .reset(cond121_reset),
    .write_en(cond121_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire121 (
    .in(cond_wire121_in),
    .out(cond_wire121_out)
);
std_reg # (
    .WIDTH(1)
) cond122 (
    .clk(cond122_clk),
    .done(cond122_done),
    .in(cond122_in),
    .out(cond122_out),
    .reset(cond122_reset),
    .write_en(cond122_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire122 (
    .in(cond_wire122_in),
    .out(cond_wire122_out)
);
std_reg # (
    .WIDTH(1)
) cond123 (
    .clk(cond123_clk),
    .done(cond123_done),
    .in(cond123_in),
    .out(cond123_out),
    .reset(cond123_reset),
    .write_en(cond123_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire123 (
    .in(cond_wire123_in),
    .out(cond_wire123_out)
);
std_reg # (
    .WIDTH(1)
) cond124 (
    .clk(cond124_clk),
    .done(cond124_done),
    .in(cond124_in),
    .out(cond124_out),
    .reset(cond124_reset),
    .write_en(cond124_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire124 (
    .in(cond_wire124_in),
    .out(cond_wire124_out)
);
std_reg # (
    .WIDTH(1)
) cond125 (
    .clk(cond125_clk),
    .done(cond125_done),
    .in(cond125_in),
    .out(cond125_out),
    .reset(cond125_reset),
    .write_en(cond125_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire125 (
    .in(cond_wire125_in),
    .out(cond_wire125_out)
);
std_reg # (
    .WIDTH(1)
) cond126 (
    .clk(cond126_clk),
    .done(cond126_done),
    .in(cond126_in),
    .out(cond126_out),
    .reset(cond126_reset),
    .write_en(cond126_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire126 (
    .in(cond_wire126_in),
    .out(cond_wire126_out)
);
std_reg # (
    .WIDTH(1)
) cond127 (
    .clk(cond127_clk),
    .done(cond127_done),
    .in(cond127_in),
    .out(cond127_out),
    .reset(cond127_reset),
    .write_en(cond127_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire127 (
    .in(cond_wire127_in),
    .out(cond_wire127_out)
);
std_reg # (
    .WIDTH(1)
) cond128 (
    .clk(cond128_clk),
    .done(cond128_done),
    .in(cond128_in),
    .out(cond128_out),
    .reset(cond128_reset),
    .write_en(cond128_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire128 (
    .in(cond_wire128_in),
    .out(cond_wire128_out)
);
std_reg # (
    .WIDTH(1)
) cond129 (
    .clk(cond129_clk),
    .done(cond129_done),
    .in(cond129_in),
    .out(cond129_out),
    .reset(cond129_reset),
    .write_en(cond129_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire129 (
    .in(cond_wire129_in),
    .out(cond_wire129_out)
);
std_reg # (
    .WIDTH(1)
) cond130 (
    .clk(cond130_clk),
    .done(cond130_done),
    .in(cond130_in),
    .out(cond130_out),
    .reset(cond130_reset),
    .write_en(cond130_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire130 (
    .in(cond_wire130_in),
    .out(cond_wire130_out)
);
std_reg # (
    .WIDTH(1)
) cond131 (
    .clk(cond131_clk),
    .done(cond131_done),
    .in(cond131_in),
    .out(cond131_out),
    .reset(cond131_reset),
    .write_en(cond131_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire131 (
    .in(cond_wire131_in),
    .out(cond_wire131_out)
);
std_reg # (
    .WIDTH(1)
) cond132 (
    .clk(cond132_clk),
    .done(cond132_done),
    .in(cond132_in),
    .out(cond132_out),
    .reset(cond132_reset),
    .write_en(cond132_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire132 (
    .in(cond_wire132_in),
    .out(cond_wire132_out)
);
std_reg # (
    .WIDTH(1)
) cond133 (
    .clk(cond133_clk),
    .done(cond133_done),
    .in(cond133_in),
    .out(cond133_out),
    .reset(cond133_reset),
    .write_en(cond133_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire133 (
    .in(cond_wire133_in),
    .out(cond_wire133_out)
);
std_reg # (
    .WIDTH(1)
) cond134 (
    .clk(cond134_clk),
    .done(cond134_done),
    .in(cond134_in),
    .out(cond134_out),
    .reset(cond134_reset),
    .write_en(cond134_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire134 (
    .in(cond_wire134_in),
    .out(cond_wire134_out)
);
std_reg # (
    .WIDTH(1)
) cond135 (
    .clk(cond135_clk),
    .done(cond135_done),
    .in(cond135_in),
    .out(cond135_out),
    .reset(cond135_reset),
    .write_en(cond135_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire135 (
    .in(cond_wire135_in),
    .out(cond_wire135_out)
);
std_reg # (
    .WIDTH(1)
) cond136 (
    .clk(cond136_clk),
    .done(cond136_done),
    .in(cond136_in),
    .out(cond136_out),
    .reset(cond136_reset),
    .write_en(cond136_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire136 (
    .in(cond_wire136_in),
    .out(cond_wire136_out)
);
std_reg # (
    .WIDTH(1)
) cond137 (
    .clk(cond137_clk),
    .done(cond137_done),
    .in(cond137_in),
    .out(cond137_out),
    .reset(cond137_reset),
    .write_en(cond137_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire137 (
    .in(cond_wire137_in),
    .out(cond_wire137_out)
);
std_reg # (
    .WIDTH(1)
) cond138 (
    .clk(cond138_clk),
    .done(cond138_done),
    .in(cond138_in),
    .out(cond138_out),
    .reset(cond138_reset),
    .write_en(cond138_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire138 (
    .in(cond_wire138_in),
    .out(cond_wire138_out)
);
std_reg # (
    .WIDTH(1)
) cond139 (
    .clk(cond139_clk),
    .done(cond139_done),
    .in(cond139_in),
    .out(cond139_out),
    .reset(cond139_reset),
    .write_en(cond139_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire139 (
    .in(cond_wire139_in),
    .out(cond_wire139_out)
);
std_reg # (
    .WIDTH(1)
) cond140 (
    .clk(cond140_clk),
    .done(cond140_done),
    .in(cond140_in),
    .out(cond140_out),
    .reset(cond140_reset),
    .write_en(cond140_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire140 (
    .in(cond_wire140_in),
    .out(cond_wire140_out)
);
std_reg # (
    .WIDTH(1)
) cond141 (
    .clk(cond141_clk),
    .done(cond141_done),
    .in(cond141_in),
    .out(cond141_out),
    .reset(cond141_reset),
    .write_en(cond141_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire141 (
    .in(cond_wire141_in),
    .out(cond_wire141_out)
);
std_reg # (
    .WIDTH(1)
) cond142 (
    .clk(cond142_clk),
    .done(cond142_done),
    .in(cond142_in),
    .out(cond142_out),
    .reset(cond142_reset),
    .write_en(cond142_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire142 (
    .in(cond_wire142_in),
    .out(cond_wire142_out)
);
std_reg # (
    .WIDTH(1)
) cond143 (
    .clk(cond143_clk),
    .done(cond143_done),
    .in(cond143_in),
    .out(cond143_out),
    .reset(cond143_reset),
    .write_en(cond143_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire143 (
    .in(cond_wire143_in),
    .out(cond_wire143_out)
);
std_reg # (
    .WIDTH(1)
) cond144 (
    .clk(cond144_clk),
    .done(cond144_done),
    .in(cond144_in),
    .out(cond144_out),
    .reset(cond144_reset),
    .write_en(cond144_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire144 (
    .in(cond_wire144_in),
    .out(cond_wire144_out)
);
std_reg # (
    .WIDTH(1)
) cond145 (
    .clk(cond145_clk),
    .done(cond145_done),
    .in(cond145_in),
    .out(cond145_out),
    .reset(cond145_reset),
    .write_en(cond145_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire145 (
    .in(cond_wire145_in),
    .out(cond_wire145_out)
);
std_reg # (
    .WIDTH(1)
) cond146 (
    .clk(cond146_clk),
    .done(cond146_done),
    .in(cond146_in),
    .out(cond146_out),
    .reset(cond146_reset),
    .write_en(cond146_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire146 (
    .in(cond_wire146_in),
    .out(cond_wire146_out)
);
std_reg # (
    .WIDTH(1)
) cond147 (
    .clk(cond147_clk),
    .done(cond147_done),
    .in(cond147_in),
    .out(cond147_out),
    .reset(cond147_reset),
    .write_en(cond147_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire147 (
    .in(cond_wire147_in),
    .out(cond_wire147_out)
);
std_reg # (
    .WIDTH(1)
) cond148 (
    .clk(cond148_clk),
    .done(cond148_done),
    .in(cond148_in),
    .out(cond148_out),
    .reset(cond148_reset),
    .write_en(cond148_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire148 (
    .in(cond_wire148_in),
    .out(cond_wire148_out)
);
std_reg # (
    .WIDTH(1)
) cond149 (
    .clk(cond149_clk),
    .done(cond149_done),
    .in(cond149_in),
    .out(cond149_out),
    .reset(cond149_reset),
    .write_en(cond149_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire149 (
    .in(cond_wire149_in),
    .out(cond_wire149_out)
);
std_reg # (
    .WIDTH(1)
) cond150 (
    .clk(cond150_clk),
    .done(cond150_done),
    .in(cond150_in),
    .out(cond150_out),
    .reset(cond150_reset),
    .write_en(cond150_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire150 (
    .in(cond_wire150_in),
    .out(cond_wire150_out)
);
std_reg # (
    .WIDTH(1)
) cond151 (
    .clk(cond151_clk),
    .done(cond151_done),
    .in(cond151_in),
    .out(cond151_out),
    .reset(cond151_reset),
    .write_en(cond151_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire151 (
    .in(cond_wire151_in),
    .out(cond_wire151_out)
);
std_reg # (
    .WIDTH(1)
) cond152 (
    .clk(cond152_clk),
    .done(cond152_done),
    .in(cond152_in),
    .out(cond152_out),
    .reset(cond152_reset),
    .write_en(cond152_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire152 (
    .in(cond_wire152_in),
    .out(cond_wire152_out)
);
std_reg # (
    .WIDTH(1)
) cond153 (
    .clk(cond153_clk),
    .done(cond153_done),
    .in(cond153_in),
    .out(cond153_out),
    .reset(cond153_reset),
    .write_en(cond153_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire153 (
    .in(cond_wire153_in),
    .out(cond_wire153_out)
);
std_reg # (
    .WIDTH(1)
) cond154 (
    .clk(cond154_clk),
    .done(cond154_done),
    .in(cond154_in),
    .out(cond154_out),
    .reset(cond154_reset),
    .write_en(cond154_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire154 (
    .in(cond_wire154_in),
    .out(cond_wire154_out)
);
std_reg # (
    .WIDTH(1)
) cond155 (
    .clk(cond155_clk),
    .done(cond155_done),
    .in(cond155_in),
    .out(cond155_out),
    .reset(cond155_reset),
    .write_en(cond155_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire155 (
    .in(cond_wire155_in),
    .out(cond_wire155_out)
);
std_reg # (
    .WIDTH(1)
) cond156 (
    .clk(cond156_clk),
    .done(cond156_done),
    .in(cond156_in),
    .out(cond156_out),
    .reset(cond156_reset),
    .write_en(cond156_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire156 (
    .in(cond_wire156_in),
    .out(cond_wire156_out)
);
std_reg # (
    .WIDTH(1)
) cond157 (
    .clk(cond157_clk),
    .done(cond157_done),
    .in(cond157_in),
    .out(cond157_out),
    .reset(cond157_reset),
    .write_en(cond157_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire157 (
    .in(cond_wire157_in),
    .out(cond_wire157_out)
);
std_reg # (
    .WIDTH(1)
) cond158 (
    .clk(cond158_clk),
    .done(cond158_done),
    .in(cond158_in),
    .out(cond158_out),
    .reset(cond158_reset),
    .write_en(cond158_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire158 (
    .in(cond_wire158_in),
    .out(cond_wire158_out)
);
std_reg # (
    .WIDTH(1)
) cond159 (
    .clk(cond159_clk),
    .done(cond159_done),
    .in(cond159_in),
    .out(cond159_out),
    .reset(cond159_reset),
    .write_en(cond159_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire159 (
    .in(cond_wire159_in),
    .out(cond_wire159_out)
);
std_reg # (
    .WIDTH(1)
) cond160 (
    .clk(cond160_clk),
    .done(cond160_done),
    .in(cond160_in),
    .out(cond160_out),
    .reset(cond160_reset),
    .write_en(cond160_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire160 (
    .in(cond_wire160_in),
    .out(cond_wire160_out)
);
std_reg # (
    .WIDTH(1)
) cond161 (
    .clk(cond161_clk),
    .done(cond161_done),
    .in(cond161_in),
    .out(cond161_out),
    .reset(cond161_reset),
    .write_en(cond161_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire161 (
    .in(cond_wire161_in),
    .out(cond_wire161_out)
);
std_reg # (
    .WIDTH(1)
) cond162 (
    .clk(cond162_clk),
    .done(cond162_done),
    .in(cond162_in),
    .out(cond162_out),
    .reset(cond162_reset),
    .write_en(cond162_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire162 (
    .in(cond_wire162_in),
    .out(cond_wire162_out)
);
std_reg # (
    .WIDTH(1)
) cond163 (
    .clk(cond163_clk),
    .done(cond163_done),
    .in(cond163_in),
    .out(cond163_out),
    .reset(cond163_reset),
    .write_en(cond163_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire163 (
    .in(cond_wire163_in),
    .out(cond_wire163_out)
);
std_reg # (
    .WIDTH(1)
) cond164 (
    .clk(cond164_clk),
    .done(cond164_done),
    .in(cond164_in),
    .out(cond164_out),
    .reset(cond164_reset),
    .write_en(cond164_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire164 (
    .in(cond_wire164_in),
    .out(cond_wire164_out)
);
std_reg # (
    .WIDTH(1)
) cond165 (
    .clk(cond165_clk),
    .done(cond165_done),
    .in(cond165_in),
    .out(cond165_out),
    .reset(cond165_reset),
    .write_en(cond165_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire165 (
    .in(cond_wire165_in),
    .out(cond_wire165_out)
);
std_reg # (
    .WIDTH(1)
) cond166 (
    .clk(cond166_clk),
    .done(cond166_done),
    .in(cond166_in),
    .out(cond166_out),
    .reset(cond166_reset),
    .write_en(cond166_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire166 (
    .in(cond_wire166_in),
    .out(cond_wire166_out)
);
std_reg # (
    .WIDTH(1)
) cond167 (
    .clk(cond167_clk),
    .done(cond167_done),
    .in(cond167_in),
    .out(cond167_out),
    .reset(cond167_reset),
    .write_en(cond167_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire167 (
    .in(cond_wire167_in),
    .out(cond_wire167_out)
);
std_reg # (
    .WIDTH(1)
) cond168 (
    .clk(cond168_clk),
    .done(cond168_done),
    .in(cond168_in),
    .out(cond168_out),
    .reset(cond168_reset),
    .write_en(cond168_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire168 (
    .in(cond_wire168_in),
    .out(cond_wire168_out)
);
std_reg # (
    .WIDTH(1)
) cond169 (
    .clk(cond169_clk),
    .done(cond169_done),
    .in(cond169_in),
    .out(cond169_out),
    .reset(cond169_reset),
    .write_en(cond169_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire169 (
    .in(cond_wire169_in),
    .out(cond_wire169_out)
);
std_reg # (
    .WIDTH(1)
) cond170 (
    .clk(cond170_clk),
    .done(cond170_done),
    .in(cond170_in),
    .out(cond170_out),
    .reset(cond170_reset),
    .write_en(cond170_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire170 (
    .in(cond_wire170_in),
    .out(cond_wire170_out)
);
std_reg # (
    .WIDTH(1)
) cond171 (
    .clk(cond171_clk),
    .done(cond171_done),
    .in(cond171_in),
    .out(cond171_out),
    .reset(cond171_reset),
    .write_en(cond171_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire171 (
    .in(cond_wire171_in),
    .out(cond_wire171_out)
);
std_reg # (
    .WIDTH(1)
) cond172 (
    .clk(cond172_clk),
    .done(cond172_done),
    .in(cond172_in),
    .out(cond172_out),
    .reset(cond172_reset),
    .write_en(cond172_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire172 (
    .in(cond_wire172_in),
    .out(cond_wire172_out)
);
std_reg # (
    .WIDTH(1)
) cond173 (
    .clk(cond173_clk),
    .done(cond173_done),
    .in(cond173_in),
    .out(cond173_out),
    .reset(cond173_reset),
    .write_en(cond173_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire173 (
    .in(cond_wire173_in),
    .out(cond_wire173_out)
);
std_reg # (
    .WIDTH(1)
) cond174 (
    .clk(cond174_clk),
    .done(cond174_done),
    .in(cond174_in),
    .out(cond174_out),
    .reset(cond174_reset),
    .write_en(cond174_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire174 (
    .in(cond_wire174_in),
    .out(cond_wire174_out)
);
std_reg # (
    .WIDTH(1)
) cond175 (
    .clk(cond175_clk),
    .done(cond175_done),
    .in(cond175_in),
    .out(cond175_out),
    .reset(cond175_reset),
    .write_en(cond175_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire175 (
    .in(cond_wire175_in),
    .out(cond_wire175_out)
);
std_reg # (
    .WIDTH(1)
) cond176 (
    .clk(cond176_clk),
    .done(cond176_done),
    .in(cond176_in),
    .out(cond176_out),
    .reset(cond176_reset),
    .write_en(cond176_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire176 (
    .in(cond_wire176_in),
    .out(cond_wire176_out)
);
std_reg # (
    .WIDTH(1)
) cond177 (
    .clk(cond177_clk),
    .done(cond177_done),
    .in(cond177_in),
    .out(cond177_out),
    .reset(cond177_reset),
    .write_en(cond177_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire177 (
    .in(cond_wire177_in),
    .out(cond_wire177_out)
);
std_reg # (
    .WIDTH(1)
) cond178 (
    .clk(cond178_clk),
    .done(cond178_done),
    .in(cond178_in),
    .out(cond178_out),
    .reset(cond178_reset),
    .write_en(cond178_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire178 (
    .in(cond_wire178_in),
    .out(cond_wire178_out)
);
std_reg # (
    .WIDTH(1)
) cond179 (
    .clk(cond179_clk),
    .done(cond179_done),
    .in(cond179_in),
    .out(cond179_out),
    .reset(cond179_reset),
    .write_en(cond179_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire179 (
    .in(cond_wire179_in),
    .out(cond_wire179_out)
);
std_reg # (
    .WIDTH(1)
) cond180 (
    .clk(cond180_clk),
    .done(cond180_done),
    .in(cond180_in),
    .out(cond180_out),
    .reset(cond180_reset),
    .write_en(cond180_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire180 (
    .in(cond_wire180_in),
    .out(cond_wire180_out)
);
std_reg # (
    .WIDTH(1)
) cond181 (
    .clk(cond181_clk),
    .done(cond181_done),
    .in(cond181_in),
    .out(cond181_out),
    .reset(cond181_reset),
    .write_en(cond181_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire181 (
    .in(cond_wire181_in),
    .out(cond_wire181_out)
);
std_reg # (
    .WIDTH(1)
) cond182 (
    .clk(cond182_clk),
    .done(cond182_done),
    .in(cond182_in),
    .out(cond182_out),
    .reset(cond182_reset),
    .write_en(cond182_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire182 (
    .in(cond_wire182_in),
    .out(cond_wire182_out)
);
std_reg # (
    .WIDTH(1)
) cond183 (
    .clk(cond183_clk),
    .done(cond183_done),
    .in(cond183_in),
    .out(cond183_out),
    .reset(cond183_reset),
    .write_en(cond183_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire183 (
    .in(cond_wire183_in),
    .out(cond_wire183_out)
);
std_reg # (
    .WIDTH(1)
) cond184 (
    .clk(cond184_clk),
    .done(cond184_done),
    .in(cond184_in),
    .out(cond184_out),
    .reset(cond184_reset),
    .write_en(cond184_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire184 (
    .in(cond_wire184_in),
    .out(cond_wire184_out)
);
std_reg # (
    .WIDTH(1)
) cond185 (
    .clk(cond185_clk),
    .done(cond185_done),
    .in(cond185_in),
    .out(cond185_out),
    .reset(cond185_reset),
    .write_en(cond185_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire185 (
    .in(cond_wire185_in),
    .out(cond_wire185_out)
);
std_reg # (
    .WIDTH(1)
) cond186 (
    .clk(cond186_clk),
    .done(cond186_done),
    .in(cond186_in),
    .out(cond186_out),
    .reset(cond186_reset),
    .write_en(cond186_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire186 (
    .in(cond_wire186_in),
    .out(cond_wire186_out)
);
std_reg # (
    .WIDTH(1)
) cond187 (
    .clk(cond187_clk),
    .done(cond187_done),
    .in(cond187_in),
    .out(cond187_out),
    .reset(cond187_reset),
    .write_en(cond187_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire187 (
    .in(cond_wire187_in),
    .out(cond_wire187_out)
);
std_reg # (
    .WIDTH(1)
) cond188 (
    .clk(cond188_clk),
    .done(cond188_done),
    .in(cond188_in),
    .out(cond188_out),
    .reset(cond188_reset),
    .write_en(cond188_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire188 (
    .in(cond_wire188_in),
    .out(cond_wire188_out)
);
std_reg # (
    .WIDTH(1)
) cond189 (
    .clk(cond189_clk),
    .done(cond189_done),
    .in(cond189_in),
    .out(cond189_out),
    .reset(cond189_reset),
    .write_en(cond189_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire189 (
    .in(cond_wire189_in),
    .out(cond_wire189_out)
);
std_reg # (
    .WIDTH(1)
) cond190 (
    .clk(cond190_clk),
    .done(cond190_done),
    .in(cond190_in),
    .out(cond190_out),
    .reset(cond190_reset),
    .write_en(cond190_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire190 (
    .in(cond_wire190_in),
    .out(cond_wire190_out)
);
std_reg # (
    .WIDTH(1)
) cond191 (
    .clk(cond191_clk),
    .done(cond191_done),
    .in(cond191_in),
    .out(cond191_out),
    .reset(cond191_reset),
    .write_en(cond191_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire191 (
    .in(cond_wire191_in),
    .out(cond_wire191_out)
);
std_reg # (
    .WIDTH(1)
) cond192 (
    .clk(cond192_clk),
    .done(cond192_done),
    .in(cond192_in),
    .out(cond192_out),
    .reset(cond192_reset),
    .write_en(cond192_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire192 (
    .in(cond_wire192_in),
    .out(cond_wire192_out)
);
std_reg # (
    .WIDTH(1)
) cond193 (
    .clk(cond193_clk),
    .done(cond193_done),
    .in(cond193_in),
    .out(cond193_out),
    .reset(cond193_reset),
    .write_en(cond193_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire193 (
    .in(cond_wire193_in),
    .out(cond_wire193_out)
);
std_reg # (
    .WIDTH(1)
) cond194 (
    .clk(cond194_clk),
    .done(cond194_done),
    .in(cond194_in),
    .out(cond194_out),
    .reset(cond194_reset),
    .write_en(cond194_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire194 (
    .in(cond_wire194_in),
    .out(cond_wire194_out)
);
std_reg # (
    .WIDTH(1)
) cond195 (
    .clk(cond195_clk),
    .done(cond195_done),
    .in(cond195_in),
    .out(cond195_out),
    .reset(cond195_reset),
    .write_en(cond195_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire195 (
    .in(cond_wire195_in),
    .out(cond_wire195_out)
);
std_reg # (
    .WIDTH(1)
) cond196 (
    .clk(cond196_clk),
    .done(cond196_done),
    .in(cond196_in),
    .out(cond196_out),
    .reset(cond196_reset),
    .write_en(cond196_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire196 (
    .in(cond_wire196_in),
    .out(cond_wire196_out)
);
std_reg # (
    .WIDTH(1)
) cond197 (
    .clk(cond197_clk),
    .done(cond197_done),
    .in(cond197_in),
    .out(cond197_out),
    .reset(cond197_reset),
    .write_en(cond197_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire197 (
    .in(cond_wire197_in),
    .out(cond_wire197_out)
);
std_reg # (
    .WIDTH(1)
) cond198 (
    .clk(cond198_clk),
    .done(cond198_done),
    .in(cond198_in),
    .out(cond198_out),
    .reset(cond198_reset),
    .write_en(cond198_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire198 (
    .in(cond_wire198_in),
    .out(cond_wire198_out)
);
std_reg # (
    .WIDTH(1)
) cond199 (
    .clk(cond199_clk),
    .done(cond199_done),
    .in(cond199_in),
    .out(cond199_out),
    .reset(cond199_reset),
    .write_en(cond199_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire199 (
    .in(cond_wire199_in),
    .out(cond_wire199_out)
);
std_reg # (
    .WIDTH(1)
) cond200 (
    .clk(cond200_clk),
    .done(cond200_done),
    .in(cond200_in),
    .out(cond200_out),
    .reset(cond200_reset),
    .write_en(cond200_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire200 (
    .in(cond_wire200_in),
    .out(cond_wire200_out)
);
std_reg # (
    .WIDTH(1)
) cond201 (
    .clk(cond201_clk),
    .done(cond201_done),
    .in(cond201_in),
    .out(cond201_out),
    .reset(cond201_reset),
    .write_en(cond201_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire201 (
    .in(cond_wire201_in),
    .out(cond_wire201_out)
);
std_reg # (
    .WIDTH(1)
) cond202 (
    .clk(cond202_clk),
    .done(cond202_done),
    .in(cond202_in),
    .out(cond202_out),
    .reset(cond202_reset),
    .write_en(cond202_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire202 (
    .in(cond_wire202_in),
    .out(cond_wire202_out)
);
std_reg # (
    .WIDTH(1)
) cond203 (
    .clk(cond203_clk),
    .done(cond203_done),
    .in(cond203_in),
    .out(cond203_out),
    .reset(cond203_reset),
    .write_en(cond203_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire203 (
    .in(cond_wire203_in),
    .out(cond_wire203_out)
);
std_reg # (
    .WIDTH(1)
) cond204 (
    .clk(cond204_clk),
    .done(cond204_done),
    .in(cond204_in),
    .out(cond204_out),
    .reset(cond204_reset),
    .write_en(cond204_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire204 (
    .in(cond_wire204_in),
    .out(cond_wire204_out)
);
std_reg # (
    .WIDTH(1)
) cond205 (
    .clk(cond205_clk),
    .done(cond205_done),
    .in(cond205_in),
    .out(cond205_out),
    .reset(cond205_reset),
    .write_en(cond205_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire205 (
    .in(cond_wire205_in),
    .out(cond_wire205_out)
);
std_reg # (
    .WIDTH(1)
) cond206 (
    .clk(cond206_clk),
    .done(cond206_done),
    .in(cond206_in),
    .out(cond206_out),
    .reset(cond206_reset),
    .write_en(cond206_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire206 (
    .in(cond_wire206_in),
    .out(cond_wire206_out)
);
std_reg # (
    .WIDTH(1)
) cond207 (
    .clk(cond207_clk),
    .done(cond207_done),
    .in(cond207_in),
    .out(cond207_out),
    .reset(cond207_reset),
    .write_en(cond207_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire207 (
    .in(cond_wire207_in),
    .out(cond_wire207_out)
);
std_reg # (
    .WIDTH(1)
) cond208 (
    .clk(cond208_clk),
    .done(cond208_done),
    .in(cond208_in),
    .out(cond208_out),
    .reset(cond208_reset),
    .write_en(cond208_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire208 (
    .in(cond_wire208_in),
    .out(cond_wire208_out)
);
std_reg # (
    .WIDTH(1)
) cond209 (
    .clk(cond209_clk),
    .done(cond209_done),
    .in(cond209_in),
    .out(cond209_out),
    .reset(cond209_reset),
    .write_en(cond209_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire209 (
    .in(cond_wire209_in),
    .out(cond_wire209_out)
);
std_reg # (
    .WIDTH(1)
) cond210 (
    .clk(cond210_clk),
    .done(cond210_done),
    .in(cond210_in),
    .out(cond210_out),
    .reset(cond210_reset),
    .write_en(cond210_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire210 (
    .in(cond_wire210_in),
    .out(cond_wire210_out)
);
std_reg # (
    .WIDTH(1)
) cond211 (
    .clk(cond211_clk),
    .done(cond211_done),
    .in(cond211_in),
    .out(cond211_out),
    .reset(cond211_reset),
    .write_en(cond211_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire211 (
    .in(cond_wire211_in),
    .out(cond_wire211_out)
);
std_reg # (
    .WIDTH(1)
) cond212 (
    .clk(cond212_clk),
    .done(cond212_done),
    .in(cond212_in),
    .out(cond212_out),
    .reset(cond212_reset),
    .write_en(cond212_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire212 (
    .in(cond_wire212_in),
    .out(cond_wire212_out)
);
std_reg # (
    .WIDTH(1)
) cond213 (
    .clk(cond213_clk),
    .done(cond213_done),
    .in(cond213_in),
    .out(cond213_out),
    .reset(cond213_reset),
    .write_en(cond213_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire213 (
    .in(cond_wire213_in),
    .out(cond_wire213_out)
);
std_reg # (
    .WIDTH(1)
) cond214 (
    .clk(cond214_clk),
    .done(cond214_done),
    .in(cond214_in),
    .out(cond214_out),
    .reset(cond214_reset),
    .write_en(cond214_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire214 (
    .in(cond_wire214_in),
    .out(cond_wire214_out)
);
std_reg # (
    .WIDTH(1)
) cond215 (
    .clk(cond215_clk),
    .done(cond215_done),
    .in(cond215_in),
    .out(cond215_out),
    .reset(cond215_reset),
    .write_en(cond215_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire215 (
    .in(cond_wire215_in),
    .out(cond_wire215_out)
);
std_reg # (
    .WIDTH(1)
) cond216 (
    .clk(cond216_clk),
    .done(cond216_done),
    .in(cond216_in),
    .out(cond216_out),
    .reset(cond216_reset),
    .write_en(cond216_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire216 (
    .in(cond_wire216_in),
    .out(cond_wire216_out)
);
std_reg # (
    .WIDTH(1)
) cond217 (
    .clk(cond217_clk),
    .done(cond217_done),
    .in(cond217_in),
    .out(cond217_out),
    .reset(cond217_reset),
    .write_en(cond217_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire217 (
    .in(cond_wire217_in),
    .out(cond_wire217_out)
);
std_reg # (
    .WIDTH(1)
) cond218 (
    .clk(cond218_clk),
    .done(cond218_done),
    .in(cond218_in),
    .out(cond218_out),
    .reset(cond218_reset),
    .write_en(cond218_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire218 (
    .in(cond_wire218_in),
    .out(cond_wire218_out)
);
std_reg # (
    .WIDTH(1)
) cond219 (
    .clk(cond219_clk),
    .done(cond219_done),
    .in(cond219_in),
    .out(cond219_out),
    .reset(cond219_reset),
    .write_en(cond219_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire219 (
    .in(cond_wire219_in),
    .out(cond_wire219_out)
);
std_reg # (
    .WIDTH(1)
) cond220 (
    .clk(cond220_clk),
    .done(cond220_done),
    .in(cond220_in),
    .out(cond220_out),
    .reset(cond220_reset),
    .write_en(cond220_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire220 (
    .in(cond_wire220_in),
    .out(cond_wire220_out)
);
std_reg # (
    .WIDTH(1)
) cond221 (
    .clk(cond221_clk),
    .done(cond221_done),
    .in(cond221_in),
    .out(cond221_out),
    .reset(cond221_reset),
    .write_en(cond221_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire221 (
    .in(cond_wire221_in),
    .out(cond_wire221_out)
);
std_reg # (
    .WIDTH(1)
) cond222 (
    .clk(cond222_clk),
    .done(cond222_done),
    .in(cond222_in),
    .out(cond222_out),
    .reset(cond222_reset),
    .write_en(cond222_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire222 (
    .in(cond_wire222_in),
    .out(cond_wire222_out)
);
std_reg # (
    .WIDTH(1)
) cond223 (
    .clk(cond223_clk),
    .done(cond223_done),
    .in(cond223_in),
    .out(cond223_out),
    .reset(cond223_reset),
    .write_en(cond223_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire223 (
    .in(cond_wire223_in),
    .out(cond_wire223_out)
);
std_reg # (
    .WIDTH(1)
) cond224 (
    .clk(cond224_clk),
    .done(cond224_done),
    .in(cond224_in),
    .out(cond224_out),
    .reset(cond224_reset),
    .write_en(cond224_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire224 (
    .in(cond_wire224_in),
    .out(cond_wire224_out)
);
std_reg # (
    .WIDTH(1)
) cond225 (
    .clk(cond225_clk),
    .done(cond225_done),
    .in(cond225_in),
    .out(cond225_out),
    .reset(cond225_reset),
    .write_en(cond225_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire225 (
    .in(cond_wire225_in),
    .out(cond_wire225_out)
);
std_reg # (
    .WIDTH(1)
) cond226 (
    .clk(cond226_clk),
    .done(cond226_done),
    .in(cond226_in),
    .out(cond226_out),
    .reset(cond226_reset),
    .write_en(cond226_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire226 (
    .in(cond_wire226_in),
    .out(cond_wire226_out)
);
std_reg # (
    .WIDTH(1)
) cond227 (
    .clk(cond227_clk),
    .done(cond227_done),
    .in(cond227_in),
    .out(cond227_out),
    .reset(cond227_reset),
    .write_en(cond227_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire227 (
    .in(cond_wire227_in),
    .out(cond_wire227_out)
);
std_reg # (
    .WIDTH(1)
) cond228 (
    .clk(cond228_clk),
    .done(cond228_done),
    .in(cond228_in),
    .out(cond228_out),
    .reset(cond228_reset),
    .write_en(cond228_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire228 (
    .in(cond_wire228_in),
    .out(cond_wire228_out)
);
std_reg # (
    .WIDTH(1)
) cond229 (
    .clk(cond229_clk),
    .done(cond229_done),
    .in(cond229_in),
    .out(cond229_out),
    .reset(cond229_reset),
    .write_en(cond229_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire229 (
    .in(cond_wire229_in),
    .out(cond_wire229_out)
);
std_reg # (
    .WIDTH(1)
) cond230 (
    .clk(cond230_clk),
    .done(cond230_done),
    .in(cond230_in),
    .out(cond230_out),
    .reset(cond230_reset),
    .write_en(cond230_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire230 (
    .in(cond_wire230_in),
    .out(cond_wire230_out)
);
std_reg # (
    .WIDTH(1)
) cond231 (
    .clk(cond231_clk),
    .done(cond231_done),
    .in(cond231_in),
    .out(cond231_out),
    .reset(cond231_reset),
    .write_en(cond231_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire231 (
    .in(cond_wire231_in),
    .out(cond_wire231_out)
);
std_reg # (
    .WIDTH(1)
) cond232 (
    .clk(cond232_clk),
    .done(cond232_done),
    .in(cond232_in),
    .out(cond232_out),
    .reset(cond232_reset),
    .write_en(cond232_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire232 (
    .in(cond_wire232_in),
    .out(cond_wire232_out)
);
std_reg # (
    .WIDTH(1)
) cond233 (
    .clk(cond233_clk),
    .done(cond233_done),
    .in(cond233_in),
    .out(cond233_out),
    .reset(cond233_reset),
    .write_en(cond233_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire233 (
    .in(cond_wire233_in),
    .out(cond_wire233_out)
);
std_reg # (
    .WIDTH(1)
) cond234 (
    .clk(cond234_clk),
    .done(cond234_done),
    .in(cond234_in),
    .out(cond234_out),
    .reset(cond234_reset),
    .write_en(cond234_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire234 (
    .in(cond_wire234_in),
    .out(cond_wire234_out)
);
std_reg # (
    .WIDTH(1)
) cond235 (
    .clk(cond235_clk),
    .done(cond235_done),
    .in(cond235_in),
    .out(cond235_out),
    .reset(cond235_reset),
    .write_en(cond235_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire235 (
    .in(cond_wire235_in),
    .out(cond_wire235_out)
);
std_reg # (
    .WIDTH(1)
) cond236 (
    .clk(cond236_clk),
    .done(cond236_done),
    .in(cond236_in),
    .out(cond236_out),
    .reset(cond236_reset),
    .write_en(cond236_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire236 (
    .in(cond_wire236_in),
    .out(cond_wire236_out)
);
std_reg # (
    .WIDTH(1)
) cond237 (
    .clk(cond237_clk),
    .done(cond237_done),
    .in(cond237_in),
    .out(cond237_out),
    .reset(cond237_reset),
    .write_en(cond237_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire237 (
    .in(cond_wire237_in),
    .out(cond_wire237_out)
);
std_reg # (
    .WIDTH(1)
) cond238 (
    .clk(cond238_clk),
    .done(cond238_done),
    .in(cond238_in),
    .out(cond238_out),
    .reset(cond238_reset),
    .write_en(cond238_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire238 (
    .in(cond_wire238_in),
    .out(cond_wire238_out)
);
std_reg # (
    .WIDTH(1)
) cond239 (
    .clk(cond239_clk),
    .done(cond239_done),
    .in(cond239_in),
    .out(cond239_out),
    .reset(cond239_reset),
    .write_en(cond239_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire239 (
    .in(cond_wire239_in),
    .out(cond_wire239_out)
);
std_reg # (
    .WIDTH(1)
) cond240 (
    .clk(cond240_clk),
    .done(cond240_done),
    .in(cond240_in),
    .out(cond240_out),
    .reset(cond240_reset),
    .write_en(cond240_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire240 (
    .in(cond_wire240_in),
    .out(cond_wire240_out)
);
std_reg # (
    .WIDTH(1)
) cond241 (
    .clk(cond241_clk),
    .done(cond241_done),
    .in(cond241_in),
    .out(cond241_out),
    .reset(cond241_reset),
    .write_en(cond241_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire241 (
    .in(cond_wire241_in),
    .out(cond_wire241_out)
);
std_reg # (
    .WIDTH(1)
) cond242 (
    .clk(cond242_clk),
    .done(cond242_done),
    .in(cond242_in),
    .out(cond242_out),
    .reset(cond242_reset),
    .write_en(cond242_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire242 (
    .in(cond_wire242_in),
    .out(cond_wire242_out)
);
std_reg # (
    .WIDTH(1)
) cond243 (
    .clk(cond243_clk),
    .done(cond243_done),
    .in(cond243_in),
    .out(cond243_out),
    .reset(cond243_reset),
    .write_en(cond243_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire243 (
    .in(cond_wire243_in),
    .out(cond_wire243_out)
);
std_reg # (
    .WIDTH(1)
) cond244 (
    .clk(cond244_clk),
    .done(cond244_done),
    .in(cond244_in),
    .out(cond244_out),
    .reset(cond244_reset),
    .write_en(cond244_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire244 (
    .in(cond_wire244_in),
    .out(cond_wire244_out)
);
std_reg # (
    .WIDTH(1)
) cond245 (
    .clk(cond245_clk),
    .done(cond245_done),
    .in(cond245_in),
    .out(cond245_out),
    .reset(cond245_reset),
    .write_en(cond245_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire245 (
    .in(cond_wire245_in),
    .out(cond_wire245_out)
);
std_reg # (
    .WIDTH(1)
) cond246 (
    .clk(cond246_clk),
    .done(cond246_done),
    .in(cond246_in),
    .out(cond246_out),
    .reset(cond246_reset),
    .write_en(cond246_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire246 (
    .in(cond_wire246_in),
    .out(cond_wire246_out)
);
std_reg # (
    .WIDTH(1)
) cond247 (
    .clk(cond247_clk),
    .done(cond247_done),
    .in(cond247_in),
    .out(cond247_out),
    .reset(cond247_reset),
    .write_en(cond247_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire247 (
    .in(cond_wire247_in),
    .out(cond_wire247_out)
);
std_reg # (
    .WIDTH(1)
) cond248 (
    .clk(cond248_clk),
    .done(cond248_done),
    .in(cond248_in),
    .out(cond248_out),
    .reset(cond248_reset),
    .write_en(cond248_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire248 (
    .in(cond_wire248_in),
    .out(cond_wire248_out)
);
std_reg # (
    .WIDTH(1)
) cond249 (
    .clk(cond249_clk),
    .done(cond249_done),
    .in(cond249_in),
    .out(cond249_out),
    .reset(cond249_reset),
    .write_en(cond249_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire249 (
    .in(cond_wire249_in),
    .out(cond_wire249_out)
);
std_reg # (
    .WIDTH(1)
) cond250 (
    .clk(cond250_clk),
    .done(cond250_done),
    .in(cond250_in),
    .out(cond250_out),
    .reset(cond250_reset),
    .write_en(cond250_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire250 (
    .in(cond_wire250_in),
    .out(cond_wire250_out)
);
std_reg # (
    .WIDTH(1)
) cond251 (
    .clk(cond251_clk),
    .done(cond251_done),
    .in(cond251_in),
    .out(cond251_out),
    .reset(cond251_reset),
    .write_en(cond251_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire251 (
    .in(cond_wire251_in),
    .out(cond_wire251_out)
);
std_reg # (
    .WIDTH(1)
) cond252 (
    .clk(cond252_clk),
    .done(cond252_done),
    .in(cond252_in),
    .out(cond252_out),
    .reset(cond252_reset),
    .write_en(cond252_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire252 (
    .in(cond_wire252_in),
    .out(cond_wire252_out)
);
std_reg # (
    .WIDTH(1)
) cond253 (
    .clk(cond253_clk),
    .done(cond253_done),
    .in(cond253_in),
    .out(cond253_out),
    .reset(cond253_reset),
    .write_en(cond253_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire253 (
    .in(cond_wire253_in),
    .out(cond_wire253_out)
);
std_reg # (
    .WIDTH(1)
) cond254 (
    .clk(cond254_clk),
    .done(cond254_done),
    .in(cond254_in),
    .out(cond254_out),
    .reset(cond254_reset),
    .write_en(cond254_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire254 (
    .in(cond_wire254_in),
    .out(cond_wire254_out)
);
std_reg # (
    .WIDTH(1)
) cond255 (
    .clk(cond255_clk),
    .done(cond255_done),
    .in(cond255_in),
    .out(cond255_out),
    .reset(cond255_reset),
    .write_en(cond255_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire255 (
    .in(cond_wire255_in),
    .out(cond_wire255_out)
);
std_reg # (
    .WIDTH(1)
) cond256 (
    .clk(cond256_clk),
    .done(cond256_done),
    .in(cond256_in),
    .out(cond256_out),
    .reset(cond256_reset),
    .write_en(cond256_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire256 (
    .in(cond_wire256_in),
    .out(cond_wire256_out)
);
std_reg # (
    .WIDTH(1)
) cond257 (
    .clk(cond257_clk),
    .done(cond257_done),
    .in(cond257_in),
    .out(cond257_out),
    .reset(cond257_reset),
    .write_en(cond257_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire257 (
    .in(cond_wire257_in),
    .out(cond_wire257_out)
);
std_reg # (
    .WIDTH(1)
) cond258 (
    .clk(cond258_clk),
    .done(cond258_done),
    .in(cond258_in),
    .out(cond258_out),
    .reset(cond258_reset),
    .write_en(cond258_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire258 (
    .in(cond_wire258_in),
    .out(cond_wire258_out)
);
std_reg # (
    .WIDTH(1)
) cond259 (
    .clk(cond259_clk),
    .done(cond259_done),
    .in(cond259_in),
    .out(cond259_out),
    .reset(cond259_reset),
    .write_en(cond259_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire259 (
    .in(cond_wire259_in),
    .out(cond_wire259_out)
);
std_reg # (
    .WIDTH(1)
) cond260 (
    .clk(cond260_clk),
    .done(cond260_done),
    .in(cond260_in),
    .out(cond260_out),
    .reset(cond260_reset),
    .write_en(cond260_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire260 (
    .in(cond_wire260_in),
    .out(cond_wire260_out)
);
std_reg # (
    .WIDTH(1)
) cond261 (
    .clk(cond261_clk),
    .done(cond261_done),
    .in(cond261_in),
    .out(cond261_out),
    .reset(cond261_reset),
    .write_en(cond261_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire261 (
    .in(cond_wire261_in),
    .out(cond_wire261_out)
);
std_reg # (
    .WIDTH(1)
) cond262 (
    .clk(cond262_clk),
    .done(cond262_done),
    .in(cond262_in),
    .out(cond262_out),
    .reset(cond262_reset),
    .write_en(cond262_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire262 (
    .in(cond_wire262_in),
    .out(cond_wire262_out)
);
std_reg # (
    .WIDTH(1)
) cond263 (
    .clk(cond263_clk),
    .done(cond263_done),
    .in(cond263_in),
    .out(cond263_out),
    .reset(cond263_reset),
    .write_en(cond263_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire263 (
    .in(cond_wire263_in),
    .out(cond_wire263_out)
);
std_reg # (
    .WIDTH(1)
) cond264 (
    .clk(cond264_clk),
    .done(cond264_done),
    .in(cond264_in),
    .out(cond264_out),
    .reset(cond264_reset),
    .write_en(cond264_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire264 (
    .in(cond_wire264_in),
    .out(cond_wire264_out)
);
std_reg # (
    .WIDTH(1)
) cond265 (
    .clk(cond265_clk),
    .done(cond265_done),
    .in(cond265_in),
    .out(cond265_out),
    .reset(cond265_reset),
    .write_en(cond265_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire265 (
    .in(cond_wire265_in),
    .out(cond_wire265_out)
);
std_reg # (
    .WIDTH(1)
) cond266 (
    .clk(cond266_clk),
    .done(cond266_done),
    .in(cond266_in),
    .out(cond266_out),
    .reset(cond266_reset),
    .write_en(cond266_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire266 (
    .in(cond_wire266_in),
    .out(cond_wire266_out)
);
std_reg # (
    .WIDTH(1)
) cond267 (
    .clk(cond267_clk),
    .done(cond267_done),
    .in(cond267_in),
    .out(cond267_out),
    .reset(cond267_reset),
    .write_en(cond267_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire267 (
    .in(cond_wire267_in),
    .out(cond_wire267_out)
);
std_reg # (
    .WIDTH(1)
) cond268 (
    .clk(cond268_clk),
    .done(cond268_done),
    .in(cond268_in),
    .out(cond268_out),
    .reset(cond268_reset),
    .write_en(cond268_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire268 (
    .in(cond_wire268_in),
    .out(cond_wire268_out)
);
std_reg # (
    .WIDTH(1)
) fsm (
    .clk(fsm_clk),
    .done(fsm_done),
    .in(fsm_in),
    .out(fsm_out),
    .reset(fsm_reset),
    .write_en(fsm_write_en)
);
undef # (
    .WIDTH(1)
) ud (
    .out(ud_out)
);
std_add # (
    .WIDTH(1)
) adder (
    .left(adder_left),
    .out(adder_out),
    .right(adder_right)
);
undef # (
    .WIDTH(1)
) ud0 (
    .out(ud0_out)
);
std_add # (
    .WIDTH(1)
) adder0 (
    .left(adder0_left),
    .out(adder0_out),
    .right(adder0_right)
);
std_reg # (
    .WIDTH(1)
) signal_reg (
    .clk(signal_reg_clk),
    .done(signal_reg_done),
    .in(signal_reg_in),
    .out(signal_reg_out),
    .reset(signal_reg_reset),
    .write_en(signal_reg_write_en)
);
std_reg # (
    .WIDTH(2)
) fsm0 (
    .clk(fsm0_clk),
    .done(fsm0_done),
    .in(fsm0_in),
    .out(fsm0_out),
    .reset(fsm0_reset),
    .write_en(fsm0_write_en)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_go (
    .in(early_reset_static_par_go_in),
    .out(early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_done (
    .in(early_reset_static_par_done_in),
    .out(early_reset_static_par_done_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par0_go (
    .in(early_reset_static_par0_go_in),
    .out(early_reset_static_par0_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par0_done (
    .in(early_reset_static_par0_done_in),
    .out(early_reset_static_par0_done_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_go (
    .in(wrapper_early_reset_static_par_go_in),
    .out(wrapper_early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_done (
    .in(wrapper_early_reset_static_par_done_in),
    .out(wrapper_early_reset_static_par_done_out)
);
std_wire # (
    .WIDTH(1)
) while_wrapper_early_reset_static_par0_go (
    .in(while_wrapper_early_reset_static_par0_go_in),
    .out(while_wrapper_early_reset_static_par0_go_out)
);
std_wire # (
    .WIDTH(1)
) while_wrapper_early_reset_static_par0_done (
    .in(while_wrapper_early_reset_static_par0_done_in),
    .out(while_wrapper_early_reset_static_par0_done_out)
);
std_wire # (
    .WIDTH(1)
) tdcc_go (
    .in(tdcc_go_in),
    .out(tdcc_go_out)
);
std_wire # (
    .WIDTH(1)
) tdcc_done (
    .in(tdcc_done_in),
    .out(tdcc_done_out)
);
wire _guard0 = 1;
wire _guard1 = early_reset_static_par0_go_out;
wire _guard2 = early_reset_static_par0_go_out;
wire _guard3 = early_reset_static_par0_go_out;
wire _guard4 = early_reset_static_par0_go_out;
wire _guard5 = cond_wire58_out;
wire _guard6 = early_reset_static_par0_go_out;
wire _guard7 = _guard5 & _guard6;
wire _guard8 = cond_wire56_out;
wire _guard9 = early_reset_static_par0_go_out;
wire _guard10 = _guard8 & _guard9;
wire _guard11 = fsm_out == 1'd0;
wire _guard12 = cond_wire56_out;
wire _guard13 = _guard11 & _guard12;
wire _guard14 = fsm_out == 1'd0;
wire _guard15 = _guard13 & _guard14;
wire _guard16 = fsm_out == 1'd0;
wire _guard17 = cond_wire58_out;
wire _guard18 = _guard16 & _guard17;
wire _guard19 = fsm_out == 1'd0;
wire _guard20 = _guard18 & _guard19;
wire _guard21 = _guard15 | _guard20;
wire _guard22 = early_reset_static_par0_go_out;
wire _guard23 = _guard21 & _guard22;
wire _guard24 = fsm_out == 1'd0;
wire _guard25 = cond_wire56_out;
wire _guard26 = _guard24 & _guard25;
wire _guard27 = fsm_out == 1'd0;
wire _guard28 = _guard26 & _guard27;
wire _guard29 = fsm_out == 1'd0;
wire _guard30 = cond_wire58_out;
wire _guard31 = _guard29 & _guard30;
wire _guard32 = fsm_out == 1'd0;
wire _guard33 = _guard31 & _guard32;
wire _guard34 = _guard28 | _guard33;
wire _guard35 = early_reset_static_par0_go_out;
wire _guard36 = _guard34 & _guard35;
wire _guard37 = fsm_out == 1'd0;
wire _guard38 = cond_wire56_out;
wire _guard39 = _guard37 & _guard38;
wire _guard40 = fsm_out == 1'd0;
wire _guard41 = _guard39 & _guard40;
wire _guard42 = fsm_out == 1'd0;
wire _guard43 = cond_wire58_out;
wire _guard44 = _guard42 & _guard43;
wire _guard45 = fsm_out == 1'd0;
wire _guard46 = _guard44 & _guard45;
wire _guard47 = _guard41 | _guard46;
wire _guard48 = early_reset_static_par0_go_out;
wire _guard49 = _guard47 & _guard48;
wire _guard50 = cond_wire70_out;
wire _guard51 = early_reset_static_par0_go_out;
wire _guard52 = _guard50 & _guard51;
wire _guard53 = cond_wire68_out;
wire _guard54 = early_reset_static_par0_go_out;
wire _guard55 = _guard53 & _guard54;
wire _guard56 = fsm_out == 1'd0;
wire _guard57 = cond_wire68_out;
wire _guard58 = _guard56 & _guard57;
wire _guard59 = fsm_out == 1'd0;
wire _guard60 = _guard58 & _guard59;
wire _guard61 = fsm_out == 1'd0;
wire _guard62 = cond_wire70_out;
wire _guard63 = _guard61 & _guard62;
wire _guard64 = fsm_out == 1'd0;
wire _guard65 = _guard63 & _guard64;
wire _guard66 = _guard60 | _guard65;
wire _guard67 = early_reset_static_par0_go_out;
wire _guard68 = _guard66 & _guard67;
wire _guard69 = fsm_out == 1'd0;
wire _guard70 = cond_wire68_out;
wire _guard71 = _guard69 & _guard70;
wire _guard72 = fsm_out == 1'd0;
wire _guard73 = _guard71 & _guard72;
wire _guard74 = fsm_out == 1'd0;
wire _guard75 = cond_wire70_out;
wire _guard76 = _guard74 & _guard75;
wire _guard77 = fsm_out == 1'd0;
wire _guard78 = _guard76 & _guard77;
wire _guard79 = _guard73 | _guard78;
wire _guard80 = early_reset_static_par0_go_out;
wire _guard81 = _guard79 & _guard80;
wire _guard82 = fsm_out == 1'd0;
wire _guard83 = cond_wire68_out;
wire _guard84 = _guard82 & _guard83;
wire _guard85 = fsm_out == 1'd0;
wire _guard86 = _guard84 & _guard85;
wire _guard87 = fsm_out == 1'd0;
wire _guard88 = cond_wire70_out;
wire _guard89 = _guard87 & _guard88;
wire _guard90 = fsm_out == 1'd0;
wire _guard91 = _guard89 & _guard90;
wire _guard92 = _guard86 | _guard91;
wire _guard93 = early_reset_static_par0_go_out;
wire _guard94 = _guard92 & _guard93;
wire _guard95 = cond_wire57_out;
wire _guard96 = early_reset_static_par0_go_out;
wire _guard97 = _guard95 & _guard96;
wire _guard98 = cond_wire57_out;
wire _guard99 = early_reset_static_par0_go_out;
wire _guard100 = _guard98 & _guard99;
wire _guard101 = cond_wire86_out;
wire _guard102 = early_reset_static_par0_go_out;
wire _guard103 = _guard101 & _guard102;
wire _guard104 = cond_wire86_out;
wire _guard105 = early_reset_static_par0_go_out;
wire _guard106 = _guard104 & _guard105;
wire _guard107 = cond_wire94_out;
wire _guard108 = early_reset_static_par0_go_out;
wire _guard109 = _guard107 & _guard108;
wire _guard110 = cond_wire94_out;
wire _guard111 = early_reset_static_par0_go_out;
wire _guard112 = _guard110 & _guard111;
wire _guard113 = cond_wire98_out;
wire _guard114 = early_reset_static_par0_go_out;
wire _guard115 = _guard113 & _guard114;
wire _guard116 = cond_wire98_out;
wire _guard117 = early_reset_static_par0_go_out;
wire _guard118 = _guard116 & _guard117;
wire _guard119 = cond_wire138_out;
wire _guard120 = early_reset_static_par0_go_out;
wire _guard121 = _guard119 & _guard120;
wire _guard122 = cond_wire138_out;
wire _guard123 = early_reset_static_par0_go_out;
wire _guard124 = _guard122 & _guard123;
wire _guard125 = cond_wire123_out;
wire _guard126 = early_reset_static_par0_go_out;
wire _guard127 = _guard125 & _guard126;
wire _guard128 = cond_wire123_out;
wire _guard129 = early_reset_static_par0_go_out;
wire _guard130 = _guard128 & _guard129;
wire _guard131 = cond_wire182_out;
wire _guard132 = early_reset_static_par0_go_out;
wire _guard133 = _guard131 & _guard132;
wire _guard134 = cond_wire180_out;
wire _guard135 = early_reset_static_par0_go_out;
wire _guard136 = _guard134 & _guard135;
wire _guard137 = fsm_out == 1'd0;
wire _guard138 = cond_wire180_out;
wire _guard139 = _guard137 & _guard138;
wire _guard140 = fsm_out == 1'd0;
wire _guard141 = _guard139 & _guard140;
wire _guard142 = fsm_out == 1'd0;
wire _guard143 = cond_wire182_out;
wire _guard144 = _guard142 & _guard143;
wire _guard145 = fsm_out == 1'd0;
wire _guard146 = _guard144 & _guard145;
wire _guard147 = _guard141 | _guard146;
wire _guard148 = early_reset_static_par0_go_out;
wire _guard149 = _guard147 & _guard148;
wire _guard150 = fsm_out == 1'd0;
wire _guard151 = cond_wire180_out;
wire _guard152 = _guard150 & _guard151;
wire _guard153 = fsm_out == 1'd0;
wire _guard154 = _guard152 & _guard153;
wire _guard155 = fsm_out == 1'd0;
wire _guard156 = cond_wire182_out;
wire _guard157 = _guard155 & _guard156;
wire _guard158 = fsm_out == 1'd0;
wire _guard159 = _guard157 & _guard158;
wire _guard160 = _guard154 | _guard159;
wire _guard161 = early_reset_static_par0_go_out;
wire _guard162 = _guard160 & _guard161;
wire _guard163 = fsm_out == 1'd0;
wire _guard164 = cond_wire180_out;
wire _guard165 = _guard163 & _guard164;
wire _guard166 = fsm_out == 1'd0;
wire _guard167 = _guard165 & _guard166;
wire _guard168 = fsm_out == 1'd0;
wire _guard169 = cond_wire182_out;
wire _guard170 = _guard168 & _guard169;
wire _guard171 = fsm_out == 1'd0;
wire _guard172 = _guard170 & _guard171;
wire _guard173 = _guard167 | _guard172;
wire _guard174 = early_reset_static_par0_go_out;
wire _guard175 = _guard173 & _guard174;
wire _guard176 = cond_wire177_out;
wire _guard177 = early_reset_static_par0_go_out;
wire _guard178 = _guard176 & _guard177;
wire _guard179 = cond_wire177_out;
wire _guard180 = early_reset_static_par0_go_out;
wire _guard181 = _guard179 & _guard180;
wire _guard182 = cond_wire210_out;
wire _guard183 = early_reset_static_par0_go_out;
wire _guard184 = _guard182 & _guard183;
wire _guard185 = cond_wire210_out;
wire _guard186 = early_reset_static_par0_go_out;
wire _guard187 = _guard185 & _guard186;
wire _guard188 = cond_wire185_out;
wire _guard189 = early_reset_static_par0_go_out;
wire _guard190 = _guard188 & _guard189;
wire _guard191 = cond_wire185_out;
wire _guard192 = early_reset_static_par0_go_out;
wire _guard193 = _guard191 & _guard192;
wire _guard194 = cond_wire218_out;
wire _guard195 = early_reset_static_par0_go_out;
wire _guard196 = _guard194 & _guard195;
wire _guard197 = cond_wire218_out;
wire _guard198 = early_reset_static_par0_go_out;
wire _guard199 = _guard197 & _guard198;
wire _guard200 = cond_wire206_out;
wire _guard201 = early_reset_static_par0_go_out;
wire _guard202 = _guard200 & _guard201;
wire _guard203 = cond_wire206_out;
wire _guard204 = early_reset_static_par0_go_out;
wire _guard205 = _guard203 & _guard204;
wire _guard206 = cond_wire14_out;
wire _guard207 = early_reset_static_par0_go_out;
wire _guard208 = _guard206 & _guard207;
wire _guard209 = cond_wire14_out;
wire _guard210 = early_reset_static_par0_go_out;
wire _guard211 = _guard209 & _guard210;
wire _guard212 = cond_wire39_out;
wire _guard213 = early_reset_static_par0_go_out;
wire _guard214 = _guard212 & _guard213;
wire _guard215 = cond_wire39_out;
wire _guard216 = early_reset_static_par0_go_out;
wire _guard217 = _guard215 & _guard216;
wire _guard218 = early_reset_static_par_go_out;
wire _guard219 = early_reset_static_par0_go_out;
wire _guard220 = _guard218 | _guard219;
wire _guard221 = early_reset_static_par0_go_out;
wire _guard222 = early_reset_static_par_go_out;
wire _guard223 = early_reset_static_par_go_out;
wire _guard224 = early_reset_static_par0_go_out;
wire _guard225 = _guard223 | _guard224;
wire _guard226 = early_reset_static_par0_go_out;
wire _guard227 = early_reset_static_par_go_out;
wire _guard228 = early_reset_static_par0_go_out;
wire _guard229 = early_reset_static_par0_go_out;
wire _guard230 = early_reset_static_par0_go_out;
wire _guard231 = early_reset_static_par0_go_out;
wire _guard232 = early_reset_static_par0_go_out;
wire _guard233 = early_reset_static_par0_go_out;
wire _guard234 = early_reset_static_par0_go_out;
wire _guard235 = ~_guard0;
wire _guard236 = early_reset_static_par0_go_out;
wire _guard237 = _guard235 & _guard236;
wire _guard238 = ~_guard0;
wire _guard239 = early_reset_static_par0_go_out;
wire _guard240 = _guard238 & _guard239;
wire _guard241 = early_reset_static_par0_go_out;
wire _guard242 = early_reset_static_par0_go_out;
wire _guard243 = ~_guard0;
wire _guard244 = early_reset_static_par0_go_out;
wire _guard245 = _guard243 & _guard244;
wire _guard246 = early_reset_static_par0_go_out;
wire _guard247 = ~_guard0;
wire _guard248 = early_reset_static_par0_go_out;
wire _guard249 = _guard247 & _guard248;
wire _guard250 = early_reset_static_par0_go_out;
wire _guard251 = ~_guard0;
wire _guard252 = early_reset_static_par0_go_out;
wire _guard253 = _guard251 & _guard252;
wire _guard254 = early_reset_static_par0_go_out;
wire _guard255 = early_reset_static_par0_go_out;
wire _guard256 = ~_guard0;
wire _guard257 = early_reset_static_par0_go_out;
wire _guard258 = _guard256 & _guard257;
wire _guard259 = early_reset_static_par0_go_out;
wire _guard260 = early_reset_static_par0_go_out;
wire _guard261 = early_reset_static_par0_go_out;
wire _guard262 = early_reset_static_par0_go_out;
wire _guard263 = early_reset_static_par0_go_out;
wire _guard264 = early_reset_static_par0_go_out;
wire _guard265 = early_reset_static_par0_go_out;
wire _guard266 = early_reset_static_par0_go_out;
wire _guard267 = ~_guard0;
wire _guard268 = early_reset_static_par0_go_out;
wire _guard269 = _guard267 & _guard268;
wire _guard270 = early_reset_static_par0_go_out;
wire _guard271 = ~_guard0;
wire _guard272 = early_reset_static_par0_go_out;
wire _guard273 = _guard271 & _guard272;
wire _guard274 = ~_guard0;
wire _guard275 = early_reset_static_par0_go_out;
wire _guard276 = _guard274 & _guard275;
wire _guard277 = early_reset_static_par0_go_out;
wire _guard278 = ~_guard0;
wire _guard279 = early_reset_static_par0_go_out;
wire _guard280 = _guard278 & _guard279;
wire _guard281 = early_reset_static_par0_go_out;
wire _guard282 = early_reset_static_par0_go_out;
wire _guard283 = ~_guard0;
wire _guard284 = early_reset_static_par0_go_out;
wire _guard285 = _guard283 & _guard284;
wire _guard286 = early_reset_static_par0_go_out;
wire _guard287 = early_reset_static_par0_go_out;
wire _guard288 = early_reset_static_par0_go_out;
wire _guard289 = early_reset_static_par0_go_out;
wire _guard290 = early_reset_static_par0_go_out;
wire _guard291 = ~_guard0;
wire _guard292 = early_reset_static_par0_go_out;
wire _guard293 = _guard291 & _guard292;
wire _guard294 = early_reset_static_par0_go_out;
wire _guard295 = ~_guard0;
wire _guard296 = early_reset_static_par0_go_out;
wire _guard297 = _guard295 & _guard296;
wire _guard298 = early_reset_static_par0_go_out;
wire _guard299 = early_reset_static_par0_go_out;
wire _guard300 = ~_guard0;
wire _guard301 = early_reset_static_par0_go_out;
wire _guard302 = _guard300 & _guard301;
wire _guard303 = early_reset_static_par0_go_out;
wire _guard304 = ~_guard0;
wire _guard305 = early_reset_static_par0_go_out;
wire _guard306 = _guard304 & _guard305;
wire _guard307 = early_reset_static_par0_go_out;
wire _guard308 = early_reset_static_par0_go_out;
wire _guard309 = early_reset_static_par0_go_out;
wire _guard310 = early_reset_static_par0_go_out;
wire _guard311 = early_reset_static_par0_go_out;
wire _guard312 = early_reset_static_par0_go_out;
wire _guard313 = ~_guard0;
wire _guard314 = early_reset_static_par0_go_out;
wire _guard315 = _guard313 & _guard314;
wire _guard316 = early_reset_static_par0_go_out;
wire _guard317 = early_reset_static_par0_go_out;
wire _guard318 = ~_guard0;
wire _guard319 = early_reset_static_par0_go_out;
wire _guard320 = _guard318 & _guard319;
wire _guard321 = early_reset_static_par0_go_out;
wire _guard322 = early_reset_static_par0_go_out;
wire _guard323 = early_reset_static_par0_go_out;
wire _guard324 = early_reset_static_par0_go_out;
wire _guard325 = early_reset_static_par_go_out;
wire _guard326 = early_reset_static_par_go_out;
wire _guard327 = early_reset_static_par0_go_out;
wire _guard328 = early_reset_static_par0_go_out;
wire _guard329 = early_reset_static_par0_go_out;
wire _guard330 = cond_wire11_out;
wire _guard331 = early_reset_static_par0_go_out;
wire _guard332 = _guard330 & _guard331;
wire _guard333 = cond_wire11_out;
wire _guard334 = early_reset_static_par0_go_out;
wire _guard335 = _guard333 & _guard334;
wire _guard336 = cond_wire16_out;
wire _guard337 = early_reset_static_par0_go_out;
wire _guard338 = _guard336 & _guard337;
wire _guard339 = cond_wire16_out;
wire _guard340 = early_reset_static_par0_go_out;
wire _guard341 = _guard339 & _guard340;
wire _guard342 = cond_wire1_out;
wire _guard343 = early_reset_static_par0_go_out;
wire _guard344 = _guard342 & _guard343;
wire _guard345 = cond_wire1_out;
wire _guard346 = early_reset_static_par0_go_out;
wire _guard347 = _guard345 & _guard346;
wire _guard348 = cond_wire50_out;
wire _guard349 = early_reset_static_par0_go_out;
wire _guard350 = _guard348 & _guard349;
wire _guard351 = cond_wire48_out;
wire _guard352 = early_reset_static_par0_go_out;
wire _guard353 = _guard351 & _guard352;
wire _guard354 = fsm_out == 1'd0;
wire _guard355 = cond_wire48_out;
wire _guard356 = _guard354 & _guard355;
wire _guard357 = fsm_out == 1'd0;
wire _guard358 = _guard356 & _guard357;
wire _guard359 = fsm_out == 1'd0;
wire _guard360 = cond_wire50_out;
wire _guard361 = _guard359 & _guard360;
wire _guard362 = fsm_out == 1'd0;
wire _guard363 = _guard361 & _guard362;
wire _guard364 = _guard358 | _guard363;
wire _guard365 = early_reset_static_par0_go_out;
wire _guard366 = _guard364 & _guard365;
wire _guard367 = fsm_out == 1'd0;
wire _guard368 = cond_wire48_out;
wire _guard369 = _guard367 & _guard368;
wire _guard370 = fsm_out == 1'd0;
wire _guard371 = _guard369 & _guard370;
wire _guard372 = fsm_out == 1'd0;
wire _guard373 = cond_wire50_out;
wire _guard374 = _guard372 & _guard373;
wire _guard375 = fsm_out == 1'd0;
wire _guard376 = _guard374 & _guard375;
wire _guard377 = _guard371 | _guard376;
wire _guard378 = early_reset_static_par0_go_out;
wire _guard379 = _guard377 & _guard378;
wire _guard380 = fsm_out == 1'd0;
wire _guard381 = cond_wire48_out;
wire _guard382 = _guard380 & _guard381;
wire _guard383 = fsm_out == 1'd0;
wire _guard384 = _guard382 & _guard383;
wire _guard385 = fsm_out == 1'd0;
wire _guard386 = cond_wire50_out;
wire _guard387 = _guard385 & _guard386;
wire _guard388 = fsm_out == 1'd0;
wire _guard389 = _guard387 & _guard388;
wire _guard390 = _guard384 | _guard389;
wire _guard391 = early_reset_static_par0_go_out;
wire _guard392 = _guard390 & _guard391;
wire _guard393 = cond_wire54_out;
wire _guard394 = early_reset_static_par0_go_out;
wire _guard395 = _guard393 & _guard394;
wire _guard396 = cond_wire52_out;
wire _guard397 = early_reset_static_par0_go_out;
wire _guard398 = _guard396 & _guard397;
wire _guard399 = fsm_out == 1'd0;
wire _guard400 = cond_wire52_out;
wire _guard401 = _guard399 & _guard400;
wire _guard402 = fsm_out == 1'd0;
wire _guard403 = _guard401 & _guard402;
wire _guard404 = fsm_out == 1'd0;
wire _guard405 = cond_wire54_out;
wire _guard406 = _guard404 & _guard405;
wire _guard407 = fsm_out == 1'd0;
wire _guard408 = _guard406 & _guard407;
wire _guard409 = _guard403 | _guard408;
wire _guard410 = early_reset_static_par0_go_out;
wire _guard411 = _guard409 & _guard410;
wire _guard412 = fsm_out == 1'd0;
wire _guard413 = cond_wire52_out;
wire _guard414 = _guard412 & _guard413;
wire _guard415 = fsm_out == 1'd0;
wire _guard416 = _guard414 & _guard415;
wire _guard417 = fsm_out == 1'd0;
wire _guard418 = cond_wire54_out;
wire _guard419 = _guard417 & _guard418;
wire _guard420 = fsm_out == 1'd0;
wire _guard421 = _guard419 & _guard420;
wire _guard422 = _guard416 | _guard421;
wire _guard423 = early_reset_static_par0_go_out;
wire _guard424 = _guard422 & _guard423;
wire _guard425 = fsm_out == 1'd0;
wire _guard426 = cond_wire52_out;
wire _guard427 = _guard425 & _guard426;
wire _guard428 = fsm_out == 1'd0;
wire _guard429 = _guard427 & _guard428;
wire _guard430 = fsm_out == 1'd0;
wire _guard431 = cond_wire54_out;
wire _guard432 = _guard430 & _guard431;
wire _guard433 = fsm_out == 1'd0;
wire _guard434 = _guard432 & _guard433;
wire _guard435 = _guard429 | _guard434;
wire _guard436 = early_reset_static_par0_go_out;
wire _guard437 = _guard435 & _guard436;
wire _guard438 = cond_wire49_out;
wire _guard439 = early_reset_static_par0_go_out;
wire _guard440 = _guard438 & _guard439;
wire _guard441 = cond_wire49_out;
wire _guard442 = early_reset_static_par0_go_out;
wire _guard443 = _guard441 & _guard442;
wire _guard444 = cond_wire94_out;
wire _guard445 = early_reset_static_par0_go_out;
wire _guard446 = _guard444 & _guard445;
wire _guard447 = cond_wire94_out;
wire _guard448 = early_reset_static_par0_go_out;
wire _guard449 = _guard447 & _guard448;
wire _guard450 = cond_wire135_out;
wire _guard451 = early_reset_static_par0_go_out;
wire _guard452 = _guard450 & _guard451;
wire _guard453 = cond_wire135_out;
wire _guard454 = early_reset_static_par0_go_out;
wire _guard455 = _guard453 & _guard454;
wire _guard456 = cond_wire173_out;
wire _guard457 = early_reset_static_par0_go_out;
wire _guard458 = _guard456 & _guard457;
wire _guard459 = cond_wire173_out;
wire _guard460 = early_reset_static_par0_go_out;
wire _guard461 = _guard459 & _guard460;
wire _guard462 = cond_wire181_out;
wire _guard463 = early_reset_static_par0_go_out;
wire _guard464 = _guard462 & _guard463;
wire _guard465 = cond_wire181_out;
wire _guard466 = early_reset_static_par0_go_out;
wire _guard467 = _guard465 & _guard466;
wire _guard468 = cond_wire223_out;
wire _guard469 = early_reset_static_par0_go_out;
wire _guard470 = _guard468 & _guard469;
wire _guard471 = cond_wire221_out;
wire _guard472 = early_reset_static_par0_go_out;
wire _guard473 = _guard471 & _guard472;
wire _guard474 = fsm_out == 1'd0;
wire _guard475 = cond_wire221_out;
wire _guard476 = _guard474 & _guard475;
wire _guard477 = fsm_out == 1'd0;
wire _guard478 = _guard476 & _guard477;
wire _guard479 = fsm_out == 1'd0;
wire _guard480 = cond_wire223_out;
wire _guard481 = _guard479 & _guard480;
wire _guard482 = fsm_out == 1'd0;
wire _guard483 = _guard481 & _guard482;
wire _guard484 = _guard478 | _guard483;
wire _guard485 = early_reset_static_par0_go_out;
wire _guard486 = _guard484 & _guard485;
wire _guard487 = fsm_out == 1'd0;
wire _guard488 = cond_wire221_out;
wire _guard489 = _guard487 & _guard488;
wire _guard490 = fsm_out == 1'd0;
wire _guard491 = _guard489 & _guard490;
wire _guard492 = fsm_out == 1'd0;
wire _guard493 = cond_wire223_out;
wire _guard494 = _guard492 & _guard493;
wire _guard495 = fsm_out == 1'd0;
wire _guard496 = _guard494 & _guard495;
wire _guard497 = _guard491 | _guard496;
wire _guard498 = early_reset_static_par0_go_out;
wire _guard499 = _guard497 & _guard498;
wire _guard500 = fsm_out == 1'd0;
wire _guard501 = cond_wire221_out;
wire _guard502 = _guard500 & _guard501;
wire _guard503 = fsm_out == 1'd0;
wire _guard504 = _guard502 & _guard503;
wire _guard505 = fsm_out == 1'd0;
wire _guard506 = cond_wire223_out;
wire _guard507 = _guard505 & _guard506;
wire _guard508 = fsm_out == 1'd0;
wire _guard509 = _guard507 & _guard508;
wire _guard510 = _guard504 | _guard509;
wire _guard511 = early_reset_static_par0_go_out;
wire _guard512 = _guard510 & _guard511;
wire _guard513 = cond_wire201_out;
wire _guard514 = early_reset_static_par0_go_out;
wire _guard515 = _guard513 & _guard514;
wire _guard516 = cond_wire201_out;
wire _guard517 = early_reset_static_par0_go_out;
wire _guard518 = _guard516 & _guard517;
wire _guard519 = cond_wire252_out;
wire _guard520 = early_reset_static_par0_go_out;
wire _guard521 = _guard519 & _guard520;
wire _guard522 = cond_wire250_out;
wire _guard523 = early_reset_static_par0_go_out;
wire _guard524 = _guard522 & _guard523;
wire _guard525 = fsm_out == 1'd0;
wire _guard526 = cond_wire250_out;
wire _guard527 = _guard525 & _guard526;
wire _guard528 = fsm_out == 1'd0;
wire _guard529 = _guard527 & _guard528;
wire _guard530 = fsm_out == 1'd0;
wire _guard531 = cond_wire252_out;
wire _guard532 = _guard530 & _guard531;
wire _guard533 = fsm_out == 1'd0;
wire _guard534 = _guard532 & _guard533;
wire _guard535 = _guard529 | _guard534;
wire _guard536 = early_reset_static_par0_go_out;
wire _guard537 = _guard535 & _guard536;
wire _guard538 = fsm_out == 1'd0;
wire _guard539 = cond_wire250_out;
wire _guard540 = _guard538 & _guard539;
wire _guard541 = fsm_out == 1'd0;
wire _guard542 = _guard540 & _guard541;
wire _guard543 = fsm_out == 1'd0;
wire _guard544 = cond_wire252_out;
wire _guard545 = _guard543 & _guard544;
wire _guard546 = fsm_out == 1'd0;
wire _guard547 = _guard545 & _guard546;
wire _guard548 = _guard542 | _guard547;
wire _guard549 = early_reset_static_par0_go_out;
wire _guard550 = _guard548 & _guard549;
wire _guard551 = fsm_out == 1'd0;
wire _guard552 = cond_wire250_out;
wire _guard553 = _guard551 & _guard552;
wire _guard554 = fsm_out == 1'd0;
wire _guard555 = _guard553 & _guard554;
wire _guard556 = fsm_out == 1'd0;
wire _guard557 = cond_wire252_out;
wire _guard558 = _guard556 & _guard557;
wire _guard559 = fsm_out == 1'd0;
wire _guard560 = _guard558 & _guard559;
wire _guard561 = _guard555 | _guard560;
wire _guard562 = early_reset_static_par0_go_out;
wire _guard563 = _guard561 & _guard562;
wire _guard564 = cond_wire251_out;
wire _guard565 = early_reset_static_par0_go_out;
wire _guard566 = _guard564 & _guard565;
wire _guard567 = cond_wire251_out;
wire _guard568 = early_reset_static_par0_go_out;
wire _guard569 = _guard567 & _guard568;
wire _guard570 = cond_wire259_out;
wire _guard571 = early_reset_static_par0_go_out;
wire _guard572 = _guard570 & _guard571;
wire _guard573 = cond_wire259_out;
wire _guard574 = early_reset_static_par0_go_out;
wire _guard575 = _guard573 & _guard574;
wire _guard576 = cond_wire234_out;
wire _guard577 = early_reset_static_par0_go_out;
wire _guard578 = _guard576 & _guard577;
wire _guard579 = cond_wire234_out;
wire _guard580 = early_reset_static_par0_go_out;
wire _guard581 = _guard579 & _guard580;
wire _guard582 = early_reset_static_par_go_out;
wire _guard583 = cond_wire105_out;
wire _guard584 = early_reset_static_par0_go_out;
wire _guard585 = _guard583 & _guard584;
wire _guard586 = _guard582 | _guard585;
wire _guard587 = cond_wire105_out;
wire _guard588 = early_reset_static_par0_go_out;
wire _guard589 = _guard587 & _guard588;
wire _guard590 = early_reset_static_par_go_out;
wire _guard591 = early_reset_static_par_go_out;
wire _guard592 = cond_wire237_out;
wire _guard593 = early_reset_static_par0_go_out;
wire _guard594 = _guard592 & _guard593;
wire _guard595 = _guard591 | _guard594;
wire _guard596 = early_reset_static_par_go_out;
wire _guard597 = cond_wire237_out;
wire _guard598 = early_reset_static_par0_go_out;
wire _guard599 = _guard597 & _guard598;
wire _guard600 = early_reset_static_par0_go_out;
wire _guard601 = early_reset_static_par0_go_out;
wire _guard602 = early_reset_static_par0_go_out;
wire _guard603 = early_reset_static_par0_go_out;
wire _guard604 = early_reset_static_par0_go_out;
wire _guard605 = early_reset_static_par0_go_out;
wire _guard606 = early_reset_static_par0_go_out;
wire _guard607 = early_reset_static_par0_go_out;
wire _guard608 = early_reset_static_par0_go_out;
wire _guard609 = early_reset_static_par0_go_out;
wire _guard610 = early_reset_static_par0_go_out;
wire _guard611 = early_reset_static_par0_go_out;
wire _guard612 = early_reset_static_par_go_out;
wire _guard613 = early_reset_static_par0_go_out;
wire _guard614 = _guard612 | _guard613;
wire _guard615 = early_reset_static_par0_go_out;
wire _guard616 = early_reset_static_par_go_out;
wire _guard617 = early_reset_static_par0_go_out;
wire _guard618 = early_reset_static_par0_go_out;
wire _guard619 = early_reset_static_par_go_out;
wire _guard620 = early_reset_static_par0_go_out;
wire _guard621 = _guard619 | _guard620;
wire _guard622 = early_reset_static_par0_go_out;
wire _guard623 = early_reset_static_par_go_out;
wire _guard624 = early_reset_static_par0_go_out;
wire _guard625 = early_reset_static_par0_go_out;
wire _guard626 = early_reset_static_par0_go_out;
wire _guard627 = early_reset_static_par0_go_out;
wire _guard628 = cond_wire9_out;
wire _guard629 = early_reset_static_par0_go_out;
wire _guard630 = _guard628 & _guard629;
wire _guard631 = cond_wire142_out;
wire _guard632 = early_reset_static_par0_go_out;
wire _guard633 = _guard631 & _guard632;
wire _guard634 = cond_wire162_out;
wire _guard635 = early_reset_static_par0_go_out;
wire _guard636 = _guard634 & _guard635;
wire _guard637 = cond_wire166_out;
wire _guard638 = early_reset_static_par0_go_out;
wire _guard639 = _guard637 & _guard638;
wire _guard640 = cond_wire150_out;
wire _guard641 = early_reset_static_par0_go_out;
wire _guard642 = _guard640 & _guard641;
wire _guard643 = cond_wire158_out;
wire _guard644 = early_reset_static_par0_go_out;
wire _guard645 = _guard643 & _guard644;
wire _guard646 = cond_wire170_out;
wire _guard647 = early_reset_static_par0_go_out;
wire _guard648 = _guard646 & _guard647;
wire _guard649 = cond_wire154_out;
wire _guard650 = early_reset_static_par0_go_out;
wire _guard651 = _guard649 & _guard650;
wire _guard652 = cond_wire146_out;
wire _guard653 = early_reset_static_par0_go_out;
wire _guard654 = _guard652 & _guard653;
wire _guard655 = tdcc_done_out;
wire _guard656 = cond_wire171_out;
wire _guard657 = early_reset_static_par0_go_out;
wire _guard658 = _guard656 & _guard657;
wire _guard659 = cond_wire_out;
wire _guard660 = early_reset_static_par0_go_out;
wire _guard661 = _guard659 & _guard660;
wire _guard662 = cond_wire63_out;
wire _guard663 = early_reset_static_par0_go_out;
wire _guard664 = _guard662 & _guard663;
wire _guard665 = cond_wire43_out;
wire _guard666 = early_reset_static_par0_go_out;
wire _guard667 = _guard665 & _guard666;
wire _guard668 = cond_wire71_out;
wire _guard669 = early_reset_static_par0_go_out;
wire _guard670 = _guard668 & _guard669;
wire _guard671 = cond_wire67_out;
wire _guard672 = early_reset_static_par0_go_out;
wire _guard673 = _guard671 & _guard672;
wire _guard674 = cond_wire51_out;
wire _guard675 = early_reset_static_par0_go_out;
wire _guard676 = _guard674 & _guard675;
wire _guard677 = cond_wire47_out;
wire _guard678 = early_reset_static_par0_go_out;
wire _guard679 = _guard677 & _guard678;
wire _guard680 = cond_wire55_out;
wire _guard681 = early_reset_static_par0_go_out;
wire _guard682 = _guard680 & _guard681;
wire _guard683 = cond_wire59_out;
wire _guard684 = early_reset_static_par0_go_out;
wire _guard685 = _guard683 & _guard684;
wire _guard686 = cond_wire195_out;
wire _guard687 = early_reset_static_par0_go_out;
wire _guard688 = _guard686 & _guard687;
wire _guard689 = cond_wire175_out;
wire _guard690 = early_reset_static_par0_go_out;
wire _guard691 = _guard689 & _guard690;
wire _guard692 = cond_wire203_out;
wire _guard693 = early_reset_static_par0_go_out;
wire _guard694 = _guard692 & _guard693;
wire _guard695 = cond_wire199_out;
wire _guard696 = early_reset_static_par0_go_out;
wire _guard697 = _guard695 & _guard696;
wire _guard698 = cond_wire183_out;
wire _guard699 = early_reset_static_par0_go_out;
wire _guard700 = _guard698 & _guard699;
wire _guard701 = cond_wire179_out;
wire _guard702 = early_reset_static_par0_go_out;
wire _guard703 = _guard701 & _guard702;
wire _guard704 = cond_wire187_out;
wire _guard705 = early_reset_static_par0_go_out;
wire _guard706 = _guard704 & _guard705;
wire _guard707 = cond_wire191_out;
wire _guard708 = early_reset_static_par0_go_out;
wire _guard709 = _guard707 & _guard708;
wire _guard710 = cond_wire183_out;
wire _guard711 = early_reset_static_par0_go_out;
wire _guard712 = _guard710 & _guard711;
wire _guard713 = cond_wire175_out;
wire _guard714 = early_reset_static_par0_go_out;
wire _guard715 = _guard713 & _guard714;
wire _guard716 = cond_wire191_out;
wire _guard717 = early_reset_static_par0_go_out;
wire _guard718 = _guard716 & _guard717;
wire _guard719 = cond_wire179_out;
wire _guard720 = early_reset_static_par0_go_out;
wire _guard721 = _guard719 & _guard720;
wire _guard722 = cond_wire203_out;
wire _guard723 = early_reset_static_par0_go_out;
wire _guard724 = _guard722 & _guard723;
wire _guard725 = cond_wire187_out;
wire _guard726 = early_reset_static_par0_go_out;
wire _guard727 = _guard725 & _guard726;
wire _guard728 = cond_wire195_out;
wire _guard729 = early_reset_static_par0_go_out;
wire _guard730 = _guard728 & _guard729;
wire _guard731 = cond_wire199_out;
wire _guard732 = early_reset_static_par0_go_out;
wire _guard733 = _guard731 & _guard732;
wire _guard734 = cond_wire204_out;
wire _guard735 = early_reset_static_par0_go_out;
wire _guard736 = _guard734 & _guard735;
wire _guard737 = cond_wire8_out;
wire _guard738 = early_reset_static_par0_go_out;
wire _guard739 = _guard737 & _guard738;
wire _guard740 = cond_wire38_out;
wire _guard741 = early_reset_static_par0_go_out;
wire _guard742 = _guard740 & _guard741;
wire _guard743 = cond_wire18_out;
wire _guard744 = early_reset_static_par0_go_out;
wire _guard745 = _guard743 & _guard744;
wire _guard746 = cond_wire28_out;
wire _guard747 = early_reset_static_par0_go_out;
wire _guard748 = _guard746 & _guard747;
wire _guard749 = cond_wire13_out;
wire _guard750 = early_reset_static_par0_go_out;
wire _guard751 = _guard749 & _guard750;
wire _guard752 = cond_wire23_out;
wire _guard753 = early_reset_static_par0_go_out;
wire _guard754 = _guard752 & _guard753;
wire _guard755 = cond_wire3_out;
wire _guard756 = early_reset_static_par0_go_out;
wire _guard757 = _guard755 & _guard756;
wire _guard758 = cond_wire33_out;
wire _guard759 = early_reset_static_par0_go_out;
wire _guard760 = _guard758 & _guard759;
wire _guard761 = cond_wire228_out;
wire _guard762 = early_reset_static_par0_go_out;
wire _guard763 = _guard761 & _guard762;
wire _guard764 = cond_wire208_out;
wire _guard765 = early_reset_static_par0_go_out;
wire _guard766 = _guard764 & _guard765;
wire _guard767 = cond_wire236_out;
wire _guard768 = early_reset_static_par0_go_out;
wire _guard769 = _guard767 & _guard768;
wire _guard770 = cond_wire232_out;
wire _guard771 = early_reset_static_par0_go_out;
wire _guard772 = _guard770 & _guard771;
wire _guard773 = cond_wire216_out;
wire _guard774 = early_reset_static_par0_go_out;
wire _guard775 = _guard773 & _guard774;
wire _guard776 = cond_wire212_out;
wire _guard777 = early_reset_static_par0_go_out;
wire _guard778 = _guard776 & _guard777;
wire _guard779 = cond_wire220_out;
wire _guard780 = early_reset_static_par0_go_out;
wire _guard781 = _guard779 & _guard780;
wire _guard782 = cond_wire224_out;
wire _guard783 = early_reset_static_par0_go_out;
wire _guard784 = _guard782 & _guard783;
wire _guard785 = cond_wire125_out;
wire _guard786 = early_reset_static_par0_go_out;
wire _guard787 = _guard785 & _guard786;
wire _guard788 = cond_wire137_out;
wire _guard789 = early_reset_static_par0_go_out;
wire _guard790 = _guard788 & _guard789;
wire _guard791 = cond_wire117_out;
wire _guard792 = early_reset_static_par0_go_out;
wire _guard793 = _guard791 & _guard792;
wire _guard794 = cond_wire129_out;
wire _guard795 = early_reset_static_par0_go_out;
wire _guard796 = _guard794 & _guard795;
wire _guard797 = cond_wire133_out;
wire _guard798 = early_reset_static_par0_go_out;
wire _guard799 = _guard797 & _guard798;
wire _guard800 = cond_wire109_out;
wire _guard801 = early_reset_static_par0_go_out;
wire _guard802 = _guard800 & _guard801;
wire _guard803 = cond_wire113_out;
wire _guard804 = early_reset_static_par0_go_out;
wire _guard805 = _guard803 & _guard804;
wire _guard806 = cond_wire121_out;
wire _guard807 = early_reset_static_par0_go_out;
wire _guard808 = _guard806 & _guard807;
wire _guard809 = cond_wire24_out;
wire _guard810 = early_reset_static_par0_go_out;
wire _guard811 = _guard809 & _guard810;
wire _guard812 = cond_wire39_out;
wire _guard813 = early_reset_static_par0_go_out;
wire _guard814 = _guard812 & _guard813;
wire _guard815 = fsm_out == 1'd0;
wire _guard816 = cond_wire175_out;
wire _guard817 = _guard815 & _guard816;
wire _guard818 = fsm_out == 1'd0;
wire _guard819 = _guard817 & _guard818;
wire _guard820 = fsm_out == 1'd0;
wire _guard821 = cond_wire179_out;
wire _guard822 = _guard820 & _guard821;
wire _guard823 = fsm_out == 1'd0;
wire _guard824 = _guard822 & _guard823;
wire _guard825 = _guard819 | _guard824;
wire _guard826 = fsm_out == 1'd0;
wire _guard827 = cond_wire183_out;
wire _guard828 = _guard826 & _guard827;
wire _guard829 = fsm_out == 1'd0;
wire _guard830 = _guard828 & _guard829;
wire _guard831 = _guard825 | _guard830;
wire _guard832 = fsm_out == 1'd0;
wire _guard833 = cond_wire187_out;
wire _guard834 = _guard832 & _guard833;
wire _guard835 = fsm_out == 1'd0;
wire _guard836 = _guard834 & _guard835;
wire _guard837 = _guard831 | _guard836;
wire _guard838 = fsm_out == 1'd0;
wire _guard839 = cond_wire191_out;
wire _guard840 = _guard838 & _guard839;
wire _guard841 = fsm_out == 1'd0;
wire _guard842 = _guard840 & _guard841;
wire _guard843 = _guard837 | _guard842;
wire _guard844 = fsm_out == 1'd0;
wire _guard845 = cond_wire195_out;
wire _guard846 = _guard844 & _guard845;
wire _guard847 = fsm_out == 1'd0;
wire _guard848 = _guard846 & _guard847;
wire _guard849 = _guard843 | _guard848;
wire _guard850 = fsm_out == 1'd0;
wire _guard851 = cond_wire199_out;
wire _guard852 = _guard850 & _guard851;
wire _guard853 = fsm_out == 1'd0;
wire _guard854 = _guard852 & _guard853;
wire _guard855 = _guard849 | _guard854;
wire _guard856 = fsm_out == 1'd0;
wire _guard857 = cond_wire203_out;
wire _guard858 = _guard856 & _guard857;
wire _guard859 = fsm_out == 1'd0;
wire _guard860 = _guard858 & _guard859;
wire _guard861 = _guard855 | _guard860;
wire _guard862 = early_reset_static_par0_go_out;
wire _guard863 = _guard861 & _guard862;
wire _guard864 = cond_wire261_out;
wire _guard865 = early_reset_static_par0_go_out;
wire _guard866 = _guard864 & _guard865;
wire _guard867 = cond_wire241_out;
wire _guard868 = early_reset_static_par0_go_out;
wire _guard869 = _guard867 & _guard868;
wire _guard870 = cond_wire268_out;
wire _guard871 = early_reset_static_par0_go_out;
wire _guard872 = _guard870 & _guard871;
wire _guard873 = cond_wire265_out;
wire _guard874 = early_reset_static_par0_go_out;
wire _guard875 = _guard873 & _guard874;
wire _guard876 = cond_wire249_out;
wire _guard877 = early_reset_static_par0_go_out;
wire _guard878 = _guard876 & _guard877;
wire _guard879 = cond_wire245_out;
wire _guard880 = early_reset_static_par0_go_out;
wire _guard881 = _guard879 & _guard880;
wire _guard882 = cond_wire253_out;
wire _guard883 = early_reset_static_par0_go_out;
wire _guard884 = _guard882 & _guard883;
wire _guard885 = cond_wire257_out;
wire _guard886 = early_reset_static_par0_go_out;
wire _guard887 = _guard885 & _guard886;
wire _guard888 = cond_wire19_out;
wire _guard889 = early_reset_static_par0_go_out;
wire _guard890 = _guard888 & _guard889;
wire _guard891 = cond_wire29_out;
wire _guard892 = early_reset_static_par0_go_out;
wire _guard893 = _guard891 & _guard892;
wire _guard894 = fsm_out == 1'd0;
wire _guard895 = cond_wire241_out;
wire _guard896 = _guard894 & _guard895;
wire _guard897 = fsm_out == 1'd0;
wire _guard898 = _guard896 & _guard897;
wire _guard899 = fsm_out == 1'd0;
wire _guard900 = cond_wire245_out;
wire _guard901 = _guard899 & _guard900;
wire _guard902 = fsm_out == 1'd0;
wire _guard903 = _guard901 & _guard902;
wire _guard904 = _guard898 | _guard903;
wire _guard905 = fsm_out == 1'd0;
wire _guard906 = cond_wire249_out;
wire _guard907 = _guard905 & _guard906;
wire _guard908 = fsm_out == 1'd0;
wire _guard909 = _guard907 & _guard908;
wire _guard910 = _guard904 | _guard909;
wire _guard911 = fsm_out == 1'd0;
wire _guard912 = cond_wire253_out;
wire _guard913 = _guard911 & _guard912;
wire _guard914 = fsm_out == 1'd0;
wire _guard915 = _guard913 & _guard914;
wire _guard916 = _guard910 | _guard915;
wire _guard917 = fsm_out == 1'd0;
wire _guard918 = cond_wire257_out;
wire _guard919 = _guard917 & _guard918;
wire _guard920 = fsm_out == 1'd0;
wire _guard921 = _guard919 & _guard920;
wire _guard922 = _guard916 | _guard921;
wire _guard923 = fsm_out == 1'd0;
wire _guard924 = cond_wire261_out;
wire _guard925 = _guard923 & _guard924;
wire _guard926 = fsm_out == 1'd0;
wire _guard927 = _guard925 & _guard926;
wire _guard928 = _guard922 | _guard927;
wire _guard929 = fsm_out == 1'd0;
wire _guard930 = cond_wire265_out;
wire _guard931 = _guard929 & _guard930;
wire _guard932 = fsm_out == 1'd0;
wire _guard933 = _guard931 & _guard932;
wire _guard934 = _guard928 | _guard933;
wire _guard935 = fsm_out == 1'd0;
wire _guard936 = cond_wire268_out;
wire _guard937 = _guard935 & _guard936;
wire _guard938 = fsm_out == 1'd0;
wire _guard939 = _guard937 & _guard938;
wire _guard940 = _guard934 | _guard939;
wire _guard941 = early_reset_static_par0_go_out;
wire _guard942 = _guard940 & _guard941;
wire _guard943 = cond_wire162_out;
wire _guard944 = early_reset_static_par0_go_out;
wire _guard945 = _guard943 & _guard944;
wire _guard946 = cond_wire142_out;
wire _guard947 = early_reset_static_par0_go_out;
wire _guard948 = _guard946 & _guard947;
wire _guard949 = cond_wire170_out;
wire _guard950 = early_reset_static_par0_go_out;
wire _guard951 = _guard949 & _guard950;
wire _guard952 = cond_wire166_out;
wire _guard953 = early_reset_static_par0_go_out;
wire _guard954 = _guard952 & _guard953;
wire _guard955 = cond_wire150_out;
wire _guard956 = early_reset_static_par0_go_out;
wire _guard957 = _guard955 & _guard956;
wire _guard958 = cond_wire146_out;
wire _guard959 = early_reset_static_par0_go_out;
wire _guard960 = _guard958 & _guard959;
wire _guard961 = cond_wire154_out;
wire _guard962 = early_reset_static_par0_go_out;
wire _guard963 = _guard961 & _guard962;
wire _guard964 = cond_wire158_out;
wire _guard965 = early_reset_static_par0_go_out;
wire _guard966 = _guard964 & _guard965;
wire _guard967 = cond_wire105_out;
wire _guard968 = early_reset_static_par0_go_out;
wire _guard969 = _guard967 & _guard968;
wire _guard970 = cond_wire104_out;
wire _guard971 = early_reset_static_par0_go_out;
wire _guard972 = _guard970 & _guard971;
wire _guard973 = cond_wire92_out;
wire _guard974 = early_reset_static_par0_go_out;
wire _guard975 = _guard973 & _guard974;
wire _guard976 = cond_wire80_out;
wire _guard977 = early_reset_static_par0_go_out;
wire _guard978 = _guard976 & _guard977;
wire _guard979 = cond_wire88_out;
wire _guard980 = early_reset_static_par0_go_out;
wire _guard981 = _guard979 & _guard980;
wire _guard982 = cond_wire96_out;
wire _guard983 = early_reset_static_par0_go_out;
wire _guard984 = _guard982 & _guard983;
wire _guard985 = cond_wire100_out;
wire _guard986 = early_reset_static_par0_go_out;
wire _guard987 = _guard985 & _guard986;
wire _guard988 = cond_wire76_out;
wire _guard989 = early_reset_static_par0_go_out;
wire _guard990 = _guard988 & _guard989;
wire _guard991 = cond_wire84_out;
wire _guard992 = early_reset_static_par0_go_out;
wire _guard993 = _guard991 & _guard992;
wire _guard994 = cond_wire138_out;
wire _guard995 = early_reset_static_par0_go_out;
wire _guard996 = _guard994 & _guard995;
wire _guard997 = cond_wire237_out;
wire _guard998 = early_reset_static_par0_go_out;
wire _guard999 = _guard997 & _guard998;
wire _guard1000 = cond_wire59_out;
wire _guard1001 = early_reset_static_par0_go_out;
wire _guard1002 = _guard1000 & _guard1001;
wire _guard1003 = cond_wire71_out;
wire _guard1004 = early_reset_static_par0_go_out;
wire _guard1005 = _guard1003 & _guard1004;
wire _guard1006 = cond_wire51_out;
wire _guard1007 = early_reset_static_par0_go_out;
wire _guard1008 = _guard1006 & _guard1007;
wire _guard1009 = cond_wire55_out;
wire _guard1010 = early_reset_static_par0_go_out;
wire _guard1011 = _guard1009 & _guard1010;
wire _guard1012 = cond_wire43_out;
wire _guard1013 = early_reset_static_par0_go_out;
wire _guard1014 = _guard1012 & _guard1013;
wire _guard1015 = cond_wire67_out;
wire _guard1016 = early_reset_static_par0_go_out;
wire _guard1017 = _guard1015 & _guard1016;
wire _guard1018 = cond_wire63_out;
wire _guard1019 = early_reset_static_par0_go_out;
wire _guard1020 = _guard1018 & _guard1019;
wire _guard1021 = cond_wire47_out;
wire _guard1022 = early_reset_static_par0_go_out;
wire _guard1023 = _guard1021 & _guard1022;
wire _guard1024 = fsm_out == 1'd0;
wire _guard1025 = cond_wire43_out;
wire _guard1026 = _guard1024 & _guard1025;
wire _guard1027 = fsm_out == 1'd0;
wire _guard1028 = _guard1026 & _guard1027;
wire _guard1029 = fsm_out == 1'd0;
wire _guard1030 = cond_wire47_out;
wire _guard1031 = _guard1029 & _guard1030;
wire _guard1032 = fsm_out == 1'd0;
wire _guard1033 = _guard1031 & _guard1032;
wire _guard1034 = _guard1028 | _guard1033;
wire _guard1035 = fsm_out == 1'd0;
wire _guard1036 = cond_wire51_out;
wire _guard1037 = _guard1035 & _guard1036;
wire _guard1038 = fsm_out == 1'd0;
wire _guard1039 = _guard1037 & _guard1038;
wire _guard1040 = _guard1034 | _guard1039;
wire _guard1041 = fsm_out == 1'd0;
wire _guard1042 = cond_wire55_out;
wire _guard1043 = _guard1041 & _guard1042;
wire _guard1044 = fsm_out == 1'd0;
wire _guard1045 = _guard1043 & _guard1044;
wire _guard1046 = _guard1040 | _guard1045;
wire _guard1047 = fsm_out == 1'd0;
wire _guard1048 = cond_wire59_out;
wire _guard1049 = _guard1047 & _guard1048;
wire _guard1050 = fsm_out == 1'd0;
wire _guard1051 = _guard1049 & _guard1050;
wire _guard1052 = _guard1046 | _guard1051;
wire _guard1053 = fsm_out == 1'd0;
wire _guard1054 = cond_wire63_out;
wire _guard1055 = _guard1053 & _guard1054;
wire _guard1056 = fsm_out == 1'd0;
wire _guard1057 = _guard1055 & _guard1056;
wire _guard1058 = _guard1052 | _guard1057;
wire _guard1059 = fsm_out == 1'd0;
wire _guard1060 = cond_wire67_out;
wire _guard1061 = _guard1059 & _guard1060;
wire _guard1062 = fsm_out == 1'd0;
wire _guard1063 = _guard1061 & _guard1062;
wire _guard1064 = _guard1058 | _guard1063;
wire _guard1065 = fsm_out == 1'd0;
wire _guard1066 = cond_wire71_out;
wire _guard1067 = _guard1065 & _guard1066;
wire _guard1068 = fsm_out == 1'd0;
wire _guard1069 = _guard1067 & _guard1068;
wire _guard1070 = _guard1064 | _guard1069;
wire _guard1071 = early_reset_static_par0_go_out;
wire _guard1072 = _guard1070 & _guard1071;
wire _guard1073 = fsm_out == 1'd0;
wire _guard1074 = cond_wire142_out;
wire _guard1075 = _guard1073 & _guard1074;
wire _guard1076 = fsm_out == 1'd0;
wire _guard1077 = _guard1075 & _guard1076;
wire _guard1078 = fsm_out == 1'd0;
wire _guard1079 = cond_wire146_out;
wire _guard1080 = _guard1078 & _guard1079;
wire _guard1081 = fsm_out == 1'd0;
wire _guard1082 = _guard1080 & _guard1081;
wire _guard1083 = _guard1077 | _guard1082;
wire _guard1084 = fsm_out == 1'd0;
wire _guard1085 = cond_wire150_out;
wire _guard1086 = _guard1084 & _guard1085;
wire _guard1087 = fsm_out == 1'd0;
wire _guard1088 = _guard1086 & _guard1087;
wire _guard1089 = _guard1083 | _guard1088;
wire _guard1090 = fsm_out == 1'd0;
wire _guard1091 = cond_wire154_out;
wire _guard1092 = _guard1090 & _guard1091;
wire _guard1093 = fsm_out == 1'd0;
wire _guard1094 = _guard1092 & _guard1093;
wire _guard1095 = _guard1089 | _guard1094;
wire _guard1096 = fsm_out == 1'd0;
wire _guard1097 = cond_wire158_out;
wire _guard1098 = _guard1096 & _guard1097;
wire _guard1099 = fsm_out == 1'd0;
wire _guard1100 = _guard1098 & _guard1099;
wire _guard1101 = _guard1095 | _guard1100;
wire _guard1102 = fsm_out == 1'd0;
wire _guard1103 = cond_wire162_out;
wire _guard1104 = _guard1102 & _guard1103;
wire _guard1105 = fsm_out == 1'd0;
wire _guard1106 = _guard1104 & _guard1105;
wire _guard1107 = _guard1101 | _guard1106;
wire _guard1108 = fsm_out == 1'd0;
wire _guard1109 = cond_wire166_out;
wire _guard1110 = _guard1108 & _guard1109;
wire _guard1111 = fsm_out == 1'd0;
wire _guard1112 = _guard1110 & _guard1111;
wire _guard1113 = _guard1107 | _guard1112;
wire _guard1114 = fsm_out == 1'd0;
wire _guard1115 = cond_wire170_out;
wire _guard1116 = _guard1114 & _guard1115;
wire _guard1117 = fsm_out == 1'd0;
wire _guard1118 = _guard1116 & _guard1117;
wire _guard1119 = _guard1113 | _guard1118;
wire _guard1120 = early_reset_static_par0_go_out;
wire _guard1121 = _guard1119 & _guard1120;
wire _guard1122 = cond_wire_out;
wire _guard1123 = early_reset_static_par0_go_out;
wire _guard1124 = _guard1122 & _guard1123;
wire _guard1125 = cond_wire4_out;
wire _guard1126 = early_reset_static_par0_go_out;
wire _guard1127 = _guard1125 & _guard1126;
wire _guard1128 = fsm_out == 1'd0;
wire _guard1129 = cond_wire3_out;
wire _guard1130 = _guard1128 & _guard1129;
wire _guard1131 = fsm_out == 1'd0;
wire _guard1132 = _guard1130 & _guard1131;
wire _guard1133 = fsm_out == 1'd0;
wire _guard1134 = cond_wire8_out;
wire _guard1135 = _guard1133 & _guard1134;
wire _guard1136 = fsm_out == 1'd0;
wire _guard1137 = _guard1135 & _guard1136;
wire _guard1138 = _guard1132 | _guard1137;
wire _guard1139 = fsm_out == 1'd0;
wire _guard1140 = cond_wire13_out;
wire _guard1141 = _guard1139 & _guard1140;
wire _guard1142 = fsm_out == 1'd0;
wire _guard1143 = _guard1141 & _guard1142;
wire _guard1144 = _guard1138 | _guard1143;
wire _guard1145 = fsm_out == 1'd0;
wire _guard1146 = cond_wire18_out;
wire _guard1147 = _guard1145 & _guard1146;
wire _guard1148 = fsm_out == 1'd0;
wire _guard1149 = _guard1147 & _guard1148;
wire _guard1150 = _guard1144 | _guard1149;
wire _guard1151 = fsm_out == 1'd0;
wire _guard1152 = cond_wire23_out;
wire _guard1153 = _guard1151 & _guard1152;
wire _guard1154 = fsm_out == 1'd0;
wire _guard1155 = _guard1153 & _guard1154;
wire _guard1156 = _guard1150 | _guard1155;
wire _guard1157 = fsm_out == 1'd0;
wire _guard1158 = cond_wire28_out;
wire _guard1159 = _guard1157 & _guard1158;
wire _guard1160 = fsm_out == 1'd0;
wire _guard1161 = _guard1159 & _guard1160;
wire _guard1162 = _guard1156 | _guard1161;
wire _guard1163 = fsm_out == 1'd0;
wire _guard1164 = cond_wire33_out;
wire _guard1165 = _guard1163 & _guard1164;
wire _guard1166 = fsm_out == 1'd0;
wire _guard1167 = _guard1165 & _guard1166;
wire _guard1168 = _guard1162 | _guard1167;
wire _guard1169 = fsm_out == 1'd0;
wire _guard1170 = cond_wire38_out;
wire _guard1171 = _guard1169 & _guard1170;
wire _guard1172 = fsm_out == 1'd0;
wire _guard1173 = _guard1171 & _guard1172;
wire _guard1174 = _guard1168 | _guard1173;
wire _guard1175 = early_reset_static_par0_go_out;
wire _guard1176 = _guard1174 & _guard1175;
wire _guard1177 = fsm_out == 1'd0;
wire _guard1178 = cond_wire76_out;
wire _guard1179 = _guard1177 & _guard1178;
wire _guard1180 = fsm_out == 1'd0;
wire _guard1181 = _guard1179 & _guard1180;
wire _guard1182 = fsm_out == 1'd0;
wire _guard1183 = cond_wire80_out;
wire _guard1184 = _guard1182 & _guard1183;
wire _guard1185 = fsm_out == 1'd0;
wire _guard1186 = _guard1184 & _guard1185;
wire _guard1187 = _guard1181 | _guard1186;
wire _guard1188 = fsm_out == 1'd0;
wire _guard1189 = cond_wire84_out;
wire _guard1190 = _guard1188 & _guard1189;
wire _guard1191 = fsm_out == 1'd0;
wire _guard1192 = _guard1190 & _guard1191;
wire _guard1193 = _guard1187 | _guard1192;
wire _guard1194 = fsm_out == 1'd0;
wire _guard1195 = cond_wire88_out;
wire _guard1196 = _guard1194 & _guard1195;
wire _guard1197 = fsm_out == 1'd0;
wire _guard1198 = _guard1196 & _guard1197;
wire _guard1199 = _guard1193 | _guard1198;
wire _guard1200 = fsm_out == 1'd0;
wire _guard1201 = cond_wire92_out;
wire _guard1202 = _guard1200 & _guard1201;
wire _guard1203 = fsm_out == 1'd0;
wire _guard1204 = _guard1202 & _guard1203;
wire _guard1205 = _guard1199 | _guard1204;
wire _guard1206 = fsm_out == 1'd0;
wire _guard1207 = cond_wire96_out;
wire _guard1208 = _guard1206 & _guard1207;
wire _guard1209 = fsm_out == 1'd0;
wire _guard1210 = _guard1208 & _guard1209;
wire _guard1211 = _guard1205 | _guard1210;
wire _guard1212 = fsm_out == 1'd0;
wire _guard1213 = cond_wire100_out;
wire _guard1214 = _guard1212 & _guard1213;
wire _guard1215 = fsm_out == 1'd0;
wire _guard1216 = _guard1214 & _guard1215;
wire _guard1217 = _guard1211 | _guard1216;
wire _guard1218 = fsm_out == 1'd0;
wire _guard1219 = cond_wire104_out;
wire _guard1220 = _guard1218 & _guard1219;
wire _guard1221 = fsm_out == 1'd0;
wire _guard1222 = _guard1220 & _guard1221;
wire _guard1223 = _guard1217 | _guard1222;
wire _guard1224 = early_reset_static_par0_go_out;
wire _guard1225 = _guard1223 & _guard1224;
wire _guard1226 = fsm_out == 1'd0;
wire _guard1227 = cond_wire109_out;
wire _guard1228 = _guard1226 & _guard1227;
wire _guard1229 = fsm_out == 1'd0;
wire _guard1230 = _guard1228 & _guard1229;
wire _guard1231 = fsm_out == 1'd0;
wire _guard1232 = cond_wire113_out;
wire _guard1233 = _guard1231 & _guard1232;
wire _guard1234 = fsm_out == 1'd0;
wire _guard1235 = _guard1233 & _guard1234;
wire _guard1236 = _guard1230 | _guard1235;
wire _guard1237 = fsm_out == 1'd0;
wire _guard1238 = cond_wire117_out;
wire _guard1239 = _guard1237 & _guard1238;
wire _guard1240 = fsm_out == 1'd0;
wire _guard1241 = _guard1239 & _guard1240;
wire _guard1242 = _guard1236 | _guard1241;
wire _guard1243 = fsm_out == 1'd0;
wire _guard1244 = cond_wire121_out;
wire _guard1245 = _guard1243 & _guard1244;
wire _guard1246 = fsm_out == 1'd0;
wire _guard1247 = _guard1245 & _guard1246;
wire _guard1248 = _guard1242 | _guard1247;
wire _guard1249 = fsm_out == 1'd0;
wire _guard1250 = cond_wire125_out;
wire _guard1251 = _guard1249 & _guard1250;
wire _guard1252 = fsm_out == 1'd0;
wire _guard1253 = _guard1251 & _guard1252;
wire _guard1254 = _guard1248 | _guard1253;
wire _guard1255 = fsm_out == 1'd0;
wire _guard1256 = cond_wire129_out;
wire _guard1257 = _guard1255 & _guard1256;
wire _guard1258 = fsm_out == 1'd0;
wire _guard1259 = _guard1257 & _guard1258;
wire _guard1260 = _guard1254 | _guard1259;
wire _guard1261 = fsm_out == 1'd0;
wire _guard1262 = cond_wire133_out;
wire _guard1263 = _guard1261 & _guard1262;
wire _guard1264 = fsm_out == 1'd0;
wire _guard1265 = _guard1263 & _guard1264;
wire _guard1266 = _guard1260 | _guard1265;
wire _guard1267 = fsm_out == 1'd0;
wire _guard1268 = cond_wire137_out;
wire _guard1269 = _guard1267 & _guard1268;
wire _guard1270 = fsm_out == 1'd0;
wire _guard1271 = _guard1269 & _guard1270;
wire _guard1272 = _guard1266 | _guard1271;
wire _guard1273 = early_reset_static_par0_go_out;
wire _guard1274 = _guard1272 & _guard1273;
wire _guard1275 = cond_wire224_out;
wire _guard1276 = early_reset_static_par0_go_out;
wire _guard1277 = _guard1275 & _guard1276;
wire _guard1278 = cond_wire208_out;
wire _guard1279 = early_reset_static_par0_go_out;
wire _guard1280 = _guard1278 & _guard1279;
wire _guard1281 = cond_wire212_out;
wire _guard1282 = early_reset_static_par0_go_out;
wire _guard1283 = _guard1281 & _guard1282;
wire _guard1284 = cond_wire228_out;
wire _guard1285 = early_reset_static_par0_go_out;
wire _guard1286 = _guard1284 & _guard1285;
wire _guard1287 = cond_wire216_out;
wire _guard1288 = early_reset_static_par0_go_out;
wire _guard1289 = _guard1287 & _guard1288;
wire _guard1290 = cond_wire220_out;
wire _guard1291 = early_reset_static_par0_go_out;
wire _guard1292 = _guard1290 & _guard1291;
wire _guard1293 = cond_wire236_out;
wire _guard1294 = early_reset_static_par0_go_out;
wire _guard1295 = _guard1293 & _guard1294;
wire _guard1296 = cond_wire232_out;
wire _guard1297 = early_reset_static_par0_go_out;
wire _guard1298 = _guard1296 & _guard1297;
wire _guard1299 = fsm_out == 1'd0;
wire _guard1300 = cond_wire208_out;
wire _guard1301 = _guard1299 & _guard1300;
wire _guard1302 = fsm_out == 1'd0;
wire _guard1303 = _guard1301 & _guard1302;
wire _guard1304 = fsm_out == 1'd0;
wire _guard1305 = cond_wire212_out;
wire _guard1306 = _guard1304 & _guard1305;
wire _guard1307 = fsm_out == 1'd0;
wire _guard1308 = _guard1306 & _guard1307;
wire _guard1309 = _guard1303 | _guard1308;
wire _guard1310 = fsm_out == 1'd0;
wire _guard1311 = cond_wire216_out;
wire _guard1312 = _guard1310 & _guard1311;
wire _guard1313 = fsm_out == 1'd0;
wire _guard1314 = _guard1312 & _guard1313;
wire _guard1315 = _guard1309 | _guard1314;
wire _guard1316 = fsm_out == 1'd0;
wire _guard1317 = cond_wire220_out;
wire _guard1318 = _guard1316 & _guard1317;
wire _guard1319 = fsm_out == 1'd0;
wire _guard1320 = _guard1318 & _guard1319;
wire _guard1321 = _guard1315 | _guard1320;
wire _guard1322 = fsm_out == 1'd0;
wire _guard1323 = cond_wire224_out;
wire _guard1324 = _guard1322 & _guard1323;
wire _guard1325 = fsm_out == 1'd0;
wire _guard1326 = _guard1324 & _guard1325;
wire _guard1327 = _guard1321 | _guard1326;
wire _guard1328 = fsm_out == 1'd0;
wire _guard1329 = cond_wire228_out;
wire _guard1330 = _guard1328 & _guard1329;
wire _guard1331 = fsm_out == 1'd0;
wire _guard1332 = _guard1330 & _guard1331;
wire _guard1333 = _guard1327 | _guard1332;
wire _guard1334 = fsm_out == 1'd0;
wire _guard1335 = cond_wire232_out;
wire _guard1336 = _guard1334 & _guard1335;
wire _guard1337 = fsm_out == 1'd0;
wire _guard1338 = _guard1336 & _guard1337;
wire _guard1339 = _guard1333 | _guard1338;
wire _guard1340 = fsm_out == 1'd0;
wire _guard1341 = cond_wire236_out;
wire _guard1342 = _guard1340 & _guard1341;
wire _guard1343 = fsm_out == 1'd0;
wire _guard1344 = _guard1342 & _guard1343;
wire _guard1345 = _guard1339 | _guard1344;
wire _guard1346 = early_reset_static_par0_go_out;
wire _guard1347 = _guard1345 & _guard1346;
wire _guard1348 = cond_wire253_out;
wire _guard1349 = early_reset_static_par0_go_out;
wire _guard1350 = _guard1348 & _guard1349;
wire _guard1351 = cond_wire257_out;
wire _guard1352 = early_reset_static_par0_go_out;
wire _guard1353 = _guard1351 & _guard1352;
wire _guard1354 = cond_wire241_out;
wire _guard1355 = early_reset_static_par0_go_out;
wire _guard1356 = _guard1354 & _guard1355;
wire _guard1357 = cond_wire261_out;
wire _guard1358 = early_reset_static_par0_go_out;
wire _guard1359 = _guard1357 & _guard1358;
wire _guard1360 = cond_wire265_out;
wire _guard1361 = early_reset_static_par0_go_out;
wire _guard1362 = _guard1360 & _guard1361;
wire _guard1363 = cond_wire245_out;
wire _guard1364 = early_reset_static_par0_go_out;
wire _guard1365 = _guard1363 & _guard1364;
wire _guard1366 = cond_wire249_out;
wire _guard1367 = early_reset_static_par0_go_out;
wire _guard1368 = _guard1366 & _guard1367;
wire _guard1369 = cond_wire268_out;
wire _guard1370 = early_reset_static_par0_go_out;
wire _guard1371 = _guard1369 & _guard1370;
wire _guard1372 = cond_wire72_out;
wire _guard1373 = early_reset_static_par0_go_out;
wire _guard1374 = _guard1372 & _guard1373;
wire _guard1375 = cond_wire28_out;
wire _guard1376 = early_reset_static_par0_go_out;
wire _guard1377 = _guard1375 & _guard1376;
wire _guard1378 = cond_wire3_out;
wire _guard1379 = early_reset_static_par0_go_out;
wire _guard1380 = _guard1378 & _guard1379;
wire _guard1381 = cond_wire38_out;
wire _guard1382 = early_reset_static_par0_go_out;
wire _guard1383 = _guard1381 & _guard1382;
wire _guard1384 = cond_wire33_out;
wire _guard1385 = early_reset_static_par0_go_out;
wire _guard1386 = _guard1384 & _guard1385;
wire _guard1387 = cond_wire13_out;
wire _guard1388 = early_reset_static_par0_go_out;
wire _guard1389 = _guard1387 & _guard1388;
wire _guard1390 = cond_wire8_out;
wire _guard1391 = early_reset_static_par0_go_out;
wire _guard1392 = _guard1390 & _guard1391;
wire _guard1393 = cond_wire18_out;
wire _guard1394 = early_reset_static_par0_go_out;
wire _guard1395 = _guard1393 & _guard1394;
wire _guard1396 = cond_wire23_out;
wire _guard1397 = early_reset_static_par0_go_out;
wire _guard1398 = _guard1396 & _guard1397;
wire _guard1399 = cond_wire129_out;
wire _guard1400 = early_reset_static_par0_go_out;
wire _guard1401 = _guard1399 & _guard1400;
wire _guard1402 = cond_wire109_out;
wire _guard1403 = early_reset_static_par0_go_out;
wire _guard1404 = _guard1402 & _guard1403;
wire _guard1405 = cond_wire137_out;
wire _guard1406 = early_reset_static_par0_go_out;
wire _guard1407 = _guard1405 & _guard1406;
wire _guard1408 = cond_wire133_out;
wire _guard1409 = early_reset_static_par0_go_out;
wire _guard1410 = _guard1408 & _guard1409;
wire _guard1411 = cond_wire117_out;
wire _guard1412 = early_reset_static_par0_go_out;
wire _guard1413 = _guard1411 & _guard1412;
wire _guard1414 = cond_wire113_out;
wire _guard1415 = early_reset_static_par0_go_out;
wire _guard1416 = _guard1414 & _guard1415;
wire _guard1417 = cond_wire121_out;
wire _guard1418 = early_reset_static_par0_go_out;
wire _guard1419 = _guard1417 & _guard1418;
wire _guard1420 = cond_wire125_out;
wire _guard1421 = early_reset_static_par0_go_out;
wire _guard1422 = _guard1420 & _guard1421;
wire _guard1423 = cond_wire14_out;
wire _guard1424 = early_reset_static_par0_go_out;
wire _guard1425 = _guard1423 & _guard1424;
wire _guard1426 = cond_wire34_out;
wire _guard1427 = early_reset_static_par0_go_out;
wire _guard1428 = _guard1426 & _guard1427;
wire _guard1429 = cond_wire96_out;
wire _guard1430 = early_reset_static_par0_go_out;
wire _guard1431 = _guard1429 & _guard1430;
wire _guard1432 = cond_wire76_out;
wire _guard1433 = early_reset_static_par0_go_out;
wire _guard1434 = _guard1432 & _guard1433;
wire _guard1435 = cond_wire104_out;
wire _guard1436 = early_reset_static_par0_go_out;
wire _guard1437 = _guard1435 & _guard1436;
wire _guard1438 = cond_wire100_out;
wire _guard1439 = early_reset_static_par0_go_out;
wire _guard1440 = _guard1438 & _guard1439;
wire _guard1441 = cond_wire84_out;
wire _guard1442 = early_reset_static_par0_go_out;
wire _guard1443 = _guard1441 & _guard1442;
wire _guard1444 = cond_wire80_out;
wire _guard1445 = early_reset_static_par0_go_out;
wire _guard1446 = _guard1444 & _guard1445;
wire _guard1447 = cond_wire88_out;
wire _guard1448 = early_reset_static_par0_go_out;
wire _guard1449 = _guard1447 & _guard1448;
wire _guard1450 = cond_wire92_out;
wire _guard1451 = early_reset_static_par0_go_out;
wire _guard1452 = _guard1450 & _guard1451;
wire _guard1453 = early_reset_static_par0_go_out;
wire _guard1454 = ~_guard0;
wire _guard1455 = early_reset_static_par0_go_out;
wire _guard1456 = _guard1454 & _guard1455;
wire _guard1457 = ~_guard0;
wire _guard1458 = early_reset_static_par0_go_out;
wire _guard1459 = _guard1457 & _guard1458;
wire _guard1460 = early_reset_static_par0_go_out;
wire _guard1461 = early_reset_static_par0_go_out;
wire _guard1462 = early_reset_static_par0_go_out;
wire _guard1463 = ~_guard0;
wire _guard1464 = early_reset_static_par0_go_out;
wire _guard1465 = _guard1463 & _guard1464;
wire _guard1466 = early_reset_static_par0_go_out;
wire _guard1467 = ~_guard0;
wire _guard1468 = early_reset_static_par0_go_out;
wire _guard1469 = _guard1467 & _guard1468;
wire _guard1470 = early_reset_static_par0_go_out;
wire _guard1471 = early_reset_static_par0_go_out;
wire _guard1472 = early_reset_static_par0_go_out;
wire _guard1473 = early_reset_static_par0_go_out;
wire _guard1474 = ~_guard0;
wire _guard1475 = early_reset_static_par0_go_out;
wire _guard1476 = _guard1474 & _guard1475;
wire _guard1477 = ~_guard0;
wire _guard1478 = early_reset_static_par0_go_out;
wire _guard1479 = _guard1477 & _guard1478;
wire _guard1480 = early_reset_static_par0_go_out;
wire _guard1481 = early_reset_static_par0_go_out;
wire _guard1482 = early_reset_static_par0_go_out;
wire _guard1483 = early_reset_static_par0_go_out;
wire _guard1484 = early_reset_static_par0_go_out;
wire _guard1485 = ~_guard0;
wire _guard1486 = early_reset_static_par0_go_out;
wire _guard1487 = _guard1485 & _guard1486;
wire _guard1488 = early_reset_static_par0_go_out;
wire _guard1489 = early_reset_static_par0_go_out;
wire _guard1490 = early_reset_static_par0_go_out;
wire _guard1491 = early_reset_static_par0_go_out;
wire _guard1492 = early_reset_static_par0_go_out;
wire _guard1493 = early_reset_static_par0_go_out;
wire _guard1494 = early_reset_static_par0_go_out;
wire _guard1495 = early_reset_static_par0_go_out;
wire _guard1496 = ~_guard0;
wire _guard1497 = early_reset_static_par0_go_out;
wire _guard1498 = _guard1496 & _guard1497;
wire _guard1499 = early_reset_static_par0_go_out;
wire _guard1500 = early_reset_static_par0_go_out;
wire _guard1501 = ~_guard0;
wire _guard1502 = early_reset_static_par0_go_out;
wire _guard1503 = _guard1501 & _guard1502;
wire _guard1504 = early_reset_static_par0_go_out;
wire _guard1505 = early_reset_static_par0_go_out;
wire _guard1506 = early_reset_static_par0_go_out;
wire _guard1507 = ~_guard0;
wire _guard1508 = early_reset_static_par0_go_out;
wire _guard1509 = _guard1507 & _guard1508;
wire _guard1510 = early_reset_static_par0_go_out;
wire _guard1511 = early_reset_static_par0_go_out;
wire _guard1512 = ~_guard0;
wire _guard1513 = early_reset_static_par0_go_out;
wire _guard1514 = _guard1512 & _guard1513;
wire _guard1515 = early_reset_static_par0_go_out;
wire _guard1516 = ~_guard0;
wire _guard1517 = early_reset_static_par0_go_out;
wire _guard1518 = _guard1516 & _guard1517;
wire _guard1519 = early_reset_static_par0_go_out;
wire _guard1520 = early_reset_static_par0_go_out;
wire _guard1521 = early_reset_static_par0_go_out;
wire _guard1522 = early_reset_static_par0_go_out;
wire _guard1523 = ~_guard0;
wire _guard1524 = early_reset_static_par0_go_out;
wire _guard1525 = _guard1523 & _guard1524;
wire _guard1526 = early_reset_static_par0_go_out;
wire _guard1527 = early_reset_static_par0_go_out;
wire _guard1528 = early_reset_static_par0_go_out;
wire _guard1529 = early_reset_static_par0_go_out;
wire _guard1530 = early_reset_static_par0_go_out;
wire _guard1531 = early_reset_static_par0_go_out;
wire _guard1532 = early_reset_static_par0_go_out;
wire _guard1533 = ~_guard0;
wire _guard1534 = early_reset_static_par0_go_out;
wire _guard1535 = _guard1533 & _guard1534;
wire _guard1536 = early_reset_static_par0_go_out;
wire _guard1537 = early_reset_static_par0_go_out;
wire _guard1538 = early_reset_static_par0_go_out;
wire _guard1539 = ~_guard0;
wire _guard1540 = early_reset_static_par0_go_out;
wire _guard1541 = _guard1539 & _guard1540;
wire _guard1542 = early_reset_static_par0_go_out;
wire _guard1543 = early_reset_static_par0_go_out;
wire _guard1544 = early_reset_static_par0_go_out;
wire _guard1545 = ~_guard0;
wire _guard1546 = early_reset_static_par0_go_out;
wire _guard1547 = _guard1545 & _guard1546;
wire _guard1548 = early_reset_static_par0_go_out;
wire _guard1549 = early_reset_static_par0_go_out;
wire _guard1550 = early_reset_static_par0_go_out;
wire _guard1551 = early_reset_static_par0_go_out;
wire _guard1552 = early_reset_static_par0_go_out;
wire _guard1553 = early_reset_static_par0_go_out;
wire _guard1554 = ~_guard0;
wire _guard1555 = early_reset_static_par0_go_out;
wire _guard1556 = _guard1554 & _guard1555;
wire _guard1557 = early_reset_static_par_go_out;
wire _guard1558 = early_reset_static_par0_go_out;
wire _guard1559 = _guard1557 | _guard1558;
wire _guard1560 = fsm_out != 1'd0;
wire _guard1561 = early_reset_static_par_go_out;
wire _guard1562 = _guard1560 & _guard1561;
wire _guard1563 = fsm_out == 1'd0;
wire _guard1564 = early_reset_static_par_go_out;
wire _guard1565 = _guard1563 & _guard1564;
wire _guard1566 = fsm_out == 1'd0;
wire _guard1567 = early_reset_static_par0_go_out;
wire _guard1568 = _guard1566 & _guard1567;
wire _guard1569 = _guard1565 | _guard1568;
wire _guard1570 = fsm_out != 1'd0;
wire _guard1571 = early_reset_static_par0_go_out;
wire _guard1572 = _guard1570 & _guard1571;
wire _guard1573 = early_reset_static_par_go_out;
wire _guard1574 = early_reset_static_par_go_out;
wire _guard1575 = while_wrapper_early_reset_static_par0_go_out;
wire _guard1576 = early_reset_static_par0_go_out;
wire _guard1577 = early_reset_static_par0_go_out;
wire _guard1578 = early_reset_static_par0_go_out;
wire _guard1579 = early_reset_static_par0_go_out;
wire _guard1580 = cond_wire29_out;
wire _guard1581 = early_reset_static_par0_go_out;
wire _guard1582 = _guard1580 & _guard1581;
wire _guard1583 = cond_wire29_out;
wire _guard1584 = early_reset_static_par0_go_out;
wire _guard1585 = _guard1583 & _guard1584;
wire _guard1586 = cond_wire53_out;
wire _guard1587 = early_reset_static_par0_go_out;
wire _guard1588 = _guard1586 & _guard1587;
wire _guard1589 = cond_wire53_out;
wire _guard1590 = early_reset_static_par0_go_out;
wire _guard1591 = _guard1589 & _guard1590;
wire _guard1592 = cond_wire26_out;
wire _guard1593 = early_reset_static_par0_go_out;
wire _guard1594 = _guard1592 & _guard1593;
wire _guard1595 = cond_wire26_out;
wire _guard1596 = early_reset_static_par0_go_out;
wire _guard1597 = _guard1595 & _guard1596;
wire _guard1598 = cond_wire57_out;
wire _guard1599 = early_reset_static_par0_go_out;
wire _guard1600 = _guard1598 & _guard1599;
wire _guard1601 = cond_wire57_out;
wire _guard1602 = early_reset_static_par0_go_out;
wire _guard1603 = _guard1601 & _guard1602;
wire _guard1604 = cond_wire124_out;
wire _guard1605 = early_reset_static_par0_go_out;
wire _guard1606 = _guard1604 & _guard1605;
wire _guard1607 = cond_wire122_out;
wire _guard1608 = early_reset_static_par0_go_out;
wire _guard1609 = _guard1607 & _guard1608;
wire _guard1610 = fsm_out == 1'd0;
wire _guard1611 = cond_wire122_out;
wire _guard1612 = _guard1610 & _guard1611;
wire _guard1613 = fsm_out == 1'd0;
wire _guard1614 = _guard1612 & _guard1613;
wire _guard1615 = fsm_out == 1'd0;
wire _guard1616 = cond_wire124_out;
wire _guard1617 = _guard1615 & _guard1616;
wire _guard1618 = fsm_out == 1'd0;
wire _guard1619 = _guard1617 & _guard1618;
wire _guard1620 = _guard1614 | _guard1619;
wire _guard1621 = early_reset_static_par0_go_out;
wire _guard1622 = _guard1620 & _guard1621;
wire _guard1623 = fsm_out == 1'd0;
wire _guard1624 = cond_wire122_out;
wire _guard1625 = _guard1623 & _guard1624;
wire _guard1626 = fsm_out == 1'd0;
wire _guard1627 = _guard1625 & _guard1626;
wire _guard1628 = fsm_out == 1'd0;
wire _guard1629 = cond_wire124_out;
wire _guard1630 = _guard1628 & _guard1629;
wire _guard1631 = fsm_out == 1'd0;
wire _guard1632 = _guard1630 & _guard1631;
wire _guard1633 = _guard1627 | _guard1632;
wire _guard1634 = early_reset_static_par0_go_out;
wire _guard1635 = _guard1633 & _guard1634;
wire _guard1636 = fsm_out == 1'd0;
wire _guard1637 = cond_wire122_out;
wire _guard1638 = _guard1636 & _guard1637;
wire _guard1639 = fsm_out == 1'd0;
wire _guard1640 = _guard1638 & _guard1639;
wire _guard1641 = fsm_out == 1'd0;
wire _guard1642 = cond_wire124_out;
wire _guard1643 = _guard1641 & _guard1642;
wire _guard1644 = fsm_out == 1'd0;
wire _guard1645 = _guard1643 & _guard1644;
wire _guard1646 = _guard1640 | _guard1645;
wire _guard1647 = early_reset_static_par0_go_out;
wire _guard1648 = _guard1646 & _guard1647;
wire _guard1649 = cond_wire136_out;
wire _guard1650 = early_reset_static_par0_go_out;
wire _guard1651 = _guard1649 & _guard1650;
wire _guard1652 = cond_wire134_out;
wire _guard1653 = early_reset_static_par0_go_out;
wire _guard1654 = _guard1652 & _guard1653;
wire _guard1655 = fsm_out == 1'd0;
wire _guard1656 = cond_wire134_out;
wire _guard1657 = _guard1655 & _guard1656;
wire _guard1658 = fsm_out == 1'd0;
wire _guard1659 = _guard1657 & _guard1658;
wire _guard1660 = fsm_out == 1'd0;
wire _guard1661 = cond_wire136_out;
wire _guard1662 = _guard1660 & _guard1661;
wire _guard1663 = fsm_out == 1'd0;
wire _guard1664 = _guard1662 & _guard1663;
wire _guard1665 = _guard1659 | _guard1664;
wire _guard1666 = early_reset_static_par0_go_out;
wire _guard1667 = _guard1665 & _guard1666;
wire _guard1668 = fsm_out == 1'd0;
wire _guard1669 = cond_wire134_out;
wire _guard1670 = _guard1668 & _guard1669;
wire _guard1671 = fsm_out == 1'd0;
wire _guard1672 = _guard1670 & _guard1671;
wire _guard1673 = fsm_out == 1'd0;
wire _guard1674 = cond_wire136_out;
wire _guard1675 = _guard1673 & _guard1674;
wire _guard1676 = fsm_out == 1'd0;
wire _guard1677 = _guard1675 & _guard1676;
wire _guard1678 = _guard1672 | _guard1677;
wire _guard1679 = early_reset_static_par0_go_out;
wire _guard1680 = _guard1678 & _guard1679;
wire _guard1681 = fsm_out == 1'd0;
wire _guard1682 = cond_wire134_out;
wire _guard1683 = _guard1681 & _guard1682;
wire _guard1684 = fsm_out == 1'd0;
wire _guard1685 = _guard1683 & _guard1684;
wire _guard1686 = fsm_out == 1'd0;
wire _guard1687 = cond_wire136_out;
wire _guard1688 = _guard1686 & _guard1687;
wire _guard1689 = fsm_out == 1'd0;
wire _guard1690 = _guard1688 & _guard1689;
wire _guard1691 = _guard1685 | _guard1690;
wire _guard1692 = early_reset_static_par0_go_out;
wire _guard1693 = _guard1691 & _guard1692;
wire _guard1694 = cond_wire141_out;
wire _guard1695 = early_reset_static_par0_go_out;
wire _guard1696 = _guard1694 & _guard1695;
wire _guard1697 = cond_wire139_out;
wire _guard1698 = early_reset_static_par0_go_out;
wire _guard1699 = _guard1697 & _guard1698;
wire _guard1700 = fsm_out == 1'd0;
wire _guard1701 = cond_wire139_out;
wire _guard1702 = _guard1700 & _guard1701;
wire _guard1703 = fsm_out == 1'd0;
wire _guard1704 = _guard1702 & _guard1703;
wire _guard1705 = fsm_out == 1'd0;
wire _guard1706 = cond_wire141_out;
wire _guard1707 = _guard1705 & _guard1706;
wire _guard1708 = fsm_out == 1'd0;
wire _guard1709 = _guard1707 & _guard1708;
wire _guard1710 = _guard1704 | _guard1709;
wire _guard1711 = early_reset_static_par0_go_out;
wire _guard1712 = _guard1710 & _guard1711;
wire _guard1713 = fsm_out == 1'd0;
wire _guard1714 = cond_wire139_out;
wire _guard1715 = _guard1713 & _guard1714;
wire _guard1716 = fsm_out == 1'd0;
wire _guard1717 = _guard1715 & _guard1716;
wire _guard1718 = fsm_out == 1'd0;
wire _guard1719 = cond_wire141_out;
wire _guard1720 = _guard1718 & _guard1719;
wire _guard1721 = fsm_out == 1'd0;
wire _guard1722 = _guard1720 & _guard1721;
wire _guard1723 = _guard1717 | _guard1722;
wire _guard1724 = early_reset_static_par0_go_out;
wire _guard1725 = _guard1723 & _guard1724;
wire _guard1726 = fsm_out == 1'd0;
wire _guard1727 = cond_wire139_out;
wire _guard1728 = _guard1726 & _guard1727;
wire _guard1729 = fsm_out == 1'd0;
wire _guard1730 = _guard1728 & _guard1729;
wire _guard1731 = fsm_out == 1'd0;
wire _guard1732 = cond_wire141_out;
wire _guard1733 = _guard1731 & _guard1732;
wire _guard1734 = fsm_out == 1'd0;
wire _guard1735 = _guard1733 & _guard1734;
wire _guard1736 = _guard1730 | _guard1735;
wire _guard1737 = early_reset_static_par0_go_out;
wire _guard1738 = _guard1736 & _guard1737;
wire _guard1739 = cond_wire144_out;
wire _guard1740 = early_reset_static_par0_go_out;
wire _guard1741 = _guard1739 & _guard1740;
wire _guard1742 = cond_wire144_out;
wire _guard1743 = early_reset_static_par0_go_out;
wire _guard1744 = _guard1742 & _guard1743;
wire _guard1745 = cond_wire174_out;
wire _guard1746 = early_reset_static_par0_go_out;
wire _guard1747 = _guard1745 & _guard1746;
wire _guard1748 = cond_wire172_out;
wire _guard1749 = early_reset_static_par0_go_out;
wire _guard1750 = _guard1748 & _guard1749;
wire _guard1751 = fsm_out == 1'd0;
wire _guard1752 = cond_wire172_out;
wire _guard1753 = _guard1751 & _guard1752;
wire _guard1754 = fsm_out == 1'd0;
wire _guard1755 = _guard1753 & _guard1754;
wire _guard1756 = fsm_out == 1'd0;
wire _guard1757 = cond_wire174_out;
wire _guard1758 = _guard1756 & _guard1757;
wire _guard1759 = fsm_out == 1'd0;
wire _guard1760 = _guard1758 & _guard1759;
wire _guard1761 = _guard1755 | _guard1760;
wire _guard1762 = early_reset_static_par0_go_out;
wire _guard1763 = _guard1761 & _guard1762;
wire _guard1764 = fsm_out == 1'd0;
wire _guard1765 = cond_wire172_out;
wire _guard1766 = _guard1764 & _guard1765;
wire _guard1767 = fsm_out == 1'd0;
wire _guard1768 = _guard1766 & _guard1767;
wire _guard1769 = fsm_out == 1'd0;
wire _guard1770 = cond_wire174_out;
wire _guard1771 = _guard1769 & _guard1770;
wire _guard1772 = fsm_out == 1'd0;
wire _guard1773 = _guard1771 & _guard1772;
wire _guard1774 = _guard1768 | _guard1773;
wire _guard1775 = early_reset_static_par0_go_out;
wire _guard1776 = _guard1774 & _guard1775;
wire _guard1777 = fsm_out == 1'd0;
wire _guard1778 = cond_wire172_out;
wire _guard1779 = _guard1777 & _guard1778;
wire _guard1780 = fsm_out == 1'd0;
wire _guard1781 = _guard1779 & _guard1780;
wire _guard1782 = fsm_out == 1'd0;
wire _guard1783 = cond_wire174_out;
wire _guard1784 = _guard1782 & _guard1783;
wire _guard1785 = fsm_out == 1'd0;
wire _guard1786 = _guard1784 & _guard1785;
wire _guard1787 = _guard1781 | _guard1786;
wire _guard1788 = early_reset_static_par0_go_out;
wire _guard1789 = _guard1787 & _guard1788;
wire _guard1790 = cond_wire193_out;
wire _guard1791 = early_reset_static_par0_go_out;
wire _guard1792 = _guard1790 & _guard1791;
wire _guard1793 = cond_wire193_out;
wire _guard1794 = early_reset_static_par0_go_out;
wire _guard1795 = _guard1793 & _guard1794;
wire _guard1796 = cond_wire222_out;
wire _guard1797 = early_reset_static_par0_go_out;
wire _guard1798 = _guard1796 & _guard1797;
wire _guard1799 = cond_wire222_out;
wire _guard1800 = early_reset_static_par0_go_out;
wire _guard1801 = _guard1799 & _guard1800;
wire _guard1802 = cond_wire197_out;
wire _guard1803 = early_reset_static_par0_go_out;
wire _guard1804 = _guard1802 & _guard1803;
wire _guard1805 = cond_wire197_out;
wire _guard1806 = early_reset_static_par0_go_out;
wire _guard1807 = _guard1805 & _guard1806;
wire _guard1808 = early_reset_static_par_go_out;
wire _guard1809 = cond_wire_out;
wire _guard1810 = early_reset_static_par0_go_out;
wire _guard1811 = _guard1809 & _guard1810;
wire _guard1812 = _guard1808 | _guard1811;
wire _guard1813 = early_reset_static_par_go_out;
wire _guard1814 = cond_wire_out;
wire _guard1815 = early_reset_static_par0_go_out;
wire _guard1816 = _guard1814 & _guard1815;
wire _guard1817 = early_reset_static_par0_go_out;
wire _guard1818 = early_reset_static_par0_go_out;
wire _guard1819 = early_reset_static_par0_go_out;
wire _guard1820 = early_reset_static_par0_go_out;
wire _guard1821 = early_reset_static_par0_go_out;
wire _guard1822 = early_reset_static_par0_go_out;
wire _guard1823 = early_reset_static_par_go_out;
wire _guard1824 = early_reset_static_par0_go_out;
wire _guard1825 = _guard1823 | _guard1824;
wire _guard1826 = early_reset_static_par_go_out;
wire _guard1827 = early_reset_static_par0_go_out;
wire _guard1828 = early_reset_static_par0_go_out;
wire _guard1829 = early_reset_static_par0_go_out;
wire _guard1830 = early_reset_static_par0_go_out;
wire _guard1831 = early_reset_static_par0_go_out;
wire _guard1832 = early_reset_static_par0_go_out;
wire _guard1833 = early_reset_static_par0_go_out;
wire _guard1834 = early_reset_static_par0_go_out;
wire _guard1835 = early_reset_static_par0_go_out;
wire _guard1836 = early_reset_static_par0_go_out;
wire _guard1837 = early_reset_static_par0_go_out;
wire _guard1838 = early_reset_static_par0_go_out;
wire _guard1839 = early_reset_static_par0_go_out;
wire _guard1840 = early_reset_static_par_go_out;
wire _guard1841 = early_reset_static_par0_go_out;
wire _guard1842 = _guard1840 | _guard1841;
wire _guard1843 = early_reset_static_par_go_out;
wire _guard1844 = early_reset_static_par0_go_out;
wire _guard1845 = early_reset_static_par_go_out;
wire _guard1846 = early_reset_static_par0_go_out;
wire _guard1847 = _guard1845 | _guard1846;
wire _guard1848 = early_reset_static_par0_go_out;
wire _guard1849 = early_reset_static_par_go_out;
wire _guard1850 = early_reset_static_par_go_out;
wire _guard1851 = early_reset_static_par0_go_out;
wire _guard1852 = _guard1850 | _guard1851;
wire _guard1853 = early_reset_static_par_go_out;
wire _guard1854 = early_reset_static_par0_go_out;
wire _guard1855 = early_reset_static_par_go_out;
wire _guard1856 = early_reset_static_par0_go_out;
wire _guard1857 = _guard1855 | _guard1856;
wire _guard1858 = early_reset_static_par_go_out;
wire _guard1859 = early_reset_static_par0_go_out;
wire _guard1860 = early_reset_static_par_go_out;
wire _guard1861 = early_reset_static_par0_go_out;
wire _guard1862 = _guard1860 | _guard1861;
wire _guard1863 = early_reset_static_par0_go_out;
wire _guard1864 = early_reset_static_par_go_out;
wire _guard1865 = early_reset_static_par0_go_out;
wire _guard1866 = early_reset_static_par0_go_out;
wire _guard1867 = early_reset_static_par0_go_out;
wire _guard1868 = early_reset_static_par0_go_out;
wire _guard1869 = early_reset_static_par0_go_out;
wire _guard1870 = early_reset_static_par0_go_out;
wire _guard1871 = ~_guard0;
wire _guard1872 = early_reset_static_par0_go_out;
wire _guard1873 = _guard1871 & _guard1872;
wire _guard1874 = early_reset_static_par0_go_out;
wire _guard1875 = early_reset_static_par0_go_out;
wire _guard1876 = early_reset_static_par0_go_out;
wire _guard1877 = early_reset_static_par0_go_out;
wire _guard1878 = ~_guard0;
wire _guard1879 = early_reset_static_par0_go_out;
wire _guard1880 = _guard1878 & _guard1879;
wire _guard1881 = ~_guard0;
wire _guard1882 = early_reset_static_par0_go_out;
wire _guard1883 = _guard1881 & _guard1882;
wire _guard1884 = early_reset_static_par0_go_out;
wire _guard1885 = early_reset_static_par0_go_out;
wire _guard1886 = early_reset_static_par0_go_out;
wire _guard1887 = ~_guard0;
wire _guard1888 = early_reset_static_par0_go_out;
wire _guard1889 = _guard1887 & _guard1888;
wire _guard1890 = early_reset_static_par0_go_out;
wire _guard1891 = ~_guard0;
wire _guard1892 = early_reset_static_par0_go_out;
wire _guard1893 = _guard1891 & _guard1892;
wire _guard1894 = early_reset_static_par0_go_out;
wire _guard1895 = early_reset_static_par0_go_out;
wire _guard1896 = early_reset_static_par0_go_out;
wire _guard1897 = ~_guard0;
wire _guard1898 = early_reset_static_par0_go_out;
wire _guard1899 = _guard1897 & _guard1898;
wire _guard1900 = early_reset_static_par0_go_out;
wire _guard1901 = early_reset_static_par0_go_out;
wire _guard1902 = early_reset_static_par0_go_out;
wire _guard1903 = early_reset_static_par0_go_out;
wire _guard1904 = early_reset_static_par0_go_out;
wire _guard1905 = early_reset_static_par0_go_out;
wire _guard1906 = early_reset_static_par0_go_out;
wire _guard1907 = early_reset_static_par0_go_out;
wire _guard1908 = early_reset_static_par0_go_out;
wire _guard1909 = early_reset_static_par0_go_out;
wire _guard1910 = early_reset_static_par0_go_out;
wire _guard1911 = early_reset_static_par0_go_out;
wire _guard1912 = ~_guard0;
wire _guard1913 = early_reset_static_par0_go_out;
wire _guard1914 = _guard1912 & _guard1913;
wire _guard1915 = ~_guard0;
wire _guard1916 = early_reset_static_par0_go_out;
wire _guard1917 = _guard1915 & _guard1916;
wire _guard1918 = early_reset_static_par0_go_out;
wire _guard1919 = ~_guard0;
wire _guard1920 = early_reset_static_par0_go_out;
wire _guard1921 = _guard1919 & _guard1920;
wire _guard1922 = early_reset_static_par0_go_out;
wire _guard1923 = early_reset_static_par0_go_out;
wire _guard1924 = early_reset_static_par0_go_out;
wire _guard1925 = early_reset_static_par0_go_out;
wire _guard1926 = early_reset_static_par0_go_out;
wire _guard1927 = early_reset_static_par0_go_out;
wire _guard1928 = ~_guard0;
wire _guard1929 = early_reset_static_par0_go_out;
wire _guard1930 = _guard1928 & _guard1929;
wire _guard1931 = early_reset_static_par0_go_out;
wire _guard1932 = ~_guard0;
wire _guard1933 = early_reset_static_par0_go_out;
wire _guard1934 = _guard1932 & _guard1933;
wire _guard1935 = early_reset_static_par0_go_out;
wire _guard1936 = early_reset_static_par0_go_out;
wire _guard1937 = early_reset_static_par0_go_out;
wire _guard1938 = early_reset_static_par0_go_out;
wire _guard1939 = early_reset_static_par0_go_out;
wire _guard1940 = early_reset_static_par0_go_out;
wire _guard1941 = ~_guard0;
wire _guard1942 = early_reset_static_par0_go_out;
wire _guard1943 = _guard1941 & _guard1942;
wire _guard1944 = early_reset_static_par0_go_out;
wire _guard1945 = cond_wire7_out;
wire _guard1946 = early_reset_static_par0_go_out;
wire _guard1947 = _guard1945 & _guard1946;
wire _guard1948 = cond_wire5_out;
wire _guard1949 = early_reset_static_par0_go_out;
wire _guard1950 = _guard1948 & _guard1949;
wire _guard1951 = fsm_out == 1'd0;
wire _guard1952 = cond_wire5_out;
wire _guard1953 = _guard1951 & _guard1952;
wire _guard1954 = fsm_out == 1'd0;
wire _guard1955 = _guard1953 & _guard1954;
wire _guard1956 = fsm_out == 1'd0;
wire _guard1957 = cond_wire7_out;
wire _guard1958 = _guard1956 & _guard1957;
wire _guard1959 = fsm_out == 1'd0;
wire _guard1960 = _guard1958 & _guard1959;
wire _guard1961 = _guard1955 | _guard1960;
wire _guard1962 = early_reset_static_par0_go_out;
wire _guard1963 = _guard1961 & _guard1962;
wire _guard1964 = fsm_out == 1'd0;
wire _guard1965 = cond_wire5_out;
wire _guard1966 = _guard1964 & _guard1965;
wire _guard1967 = fsm_out == 1'd0;
wire _guard1968 = _guard1966 & _guard1967;
wire _guard1969 = fsm_out == 1'd0;
wire _guard1970 = cond_wire7_out;
wire _guard1971 = _guard1969 & _guard1970;
wire _guard1972 = fsm_out == 1'd0;
wire _guard1973 = _guard1971 & _guard1972;
wire _guard1974 = _guard1968 | _guard1973;
wire _guard1975 = early_reset_static_par0_go_out;
wire _guard1976 = _guard1974 & _guard1975;
wire _guard1977 = fsm_out == 1'd0;
wire _guard1978 = cond_wire5_out;
wire _guard1979 = _guard1977 & _guard1978;
wire _guard1980 = fsm_out == 1'd0;
wire _guard1981 = _guard1979 & _guard1980;
wire _guard1982 = fsm_out == 1'd0;
wire _guard1983 = cond_wire7_out;
wire _guard1984 = _guard1982 & _guard1983;
wire _guard1985 = fsm_out == 1'd0;
wire _guard1986 = _guard1984 & _guard1985;
wire _guard1987 = _guard1981 | _guard1986;
wire _guard1988 = early_reset_static_par0_go_out;
wire _guard1989 = _guard1987 & _guard1988;
wire _guard1990 = cond_wire26_out;
wire _guard1991 = early_reset_static_par0_go_out;
wire _guard1992 = _guard1990 & _guard1991;
wire _guard1993 = cond_wire26_out;
wire _guard1994 = early_reset_static_par0_go_out;
wire _guard1995 = _guard1993 & _guard1994;
wire _guard1996 = cond_wire37_out;
wire _guard1997 = early_reset_static_par0_go_out;
wire _guard1998 = _guard1996 & _guard1997;
wire _guard1999 = cond_wire35_out;
wire _guard2000 = early_reset_static_par0_go_out;
wire _guard2001 = _guard1999 & _guard2000;
wire _guard2002 = fsm_out == 1'd0;
wire _guard2003 = cond_wire35_out;
wire _guard2004 = _guard2002 & _guard2003;
wire _guard2005 = fsm_out == 1'd0;
wire _guard2006 = _guard2004 & _guard2005;
wire _guard2007 = fsm_out == 1'd0;
wire _guard2008 = cond_wire37_out;
wire _guard2009 = _guard2007 & _guard2008;
wire _guard2010 = fsm_out == 1'd0;
wire _guard2011 = _guard2009 & _guard2010;
wire _guard2012 = _guard2006 | _guard2011;
wire _guard2013 = early_reset_static_par0_go_out;
wire _guard2014 = _guard2012 & _guard2013;
wire _guard2015 = fsm_out == 1'd0;
wire _guard2016 = cond_wire35_out;
wire _guard2017 = _guard2015 & _guard2016;
wire _guard2018 = fsm_out == 1'd0;
wire _guard2019 = _guard2017 & _guard2018;
wire _guard2020 = fsm_out == 1'd0;
wire _guard2021 = cond_wire37_out;
wire _guard2022 = _guard2020 & _guard2021;
wire _guard2023 = fsm_out == 1'd0;
wire _guard2024 = _guard2022 & _guard2023;
wire _guard2025 = _guard2019 | _guard2024;
wire _guard2026 = early_reset_static_par0_go_out;
wire _guard2027 = _guard2025 & _guard2026;
wire _guard2028 = fsm_out == 1'd0;
wire _guard2029 = cond_wire35_out;
wire _guard2030 = _guard2028 & _guard2029;
wire _guard2031 = fsm_out == 1'd0;
wire _guard2032 = _guard2030 & _guard2031;
wire _guard2033 = fsm_out == 1'd0;
wire _guard2034 = cond_wire37_out;
wire _guard2035 = _guard2033 & _guard2034;
wire _guard2036 = fsm_out == 1'd0;
wire _guard2037 = _guard2035 & _guard2036;
wire _guard2038 = _guard2032 | _guard2037;
wire _guard2039 = early_reset_static_par0_go_out;
wire _guard2040 = _guard2038 & _guard2039;
wire _guard2041 = cond_wire45_out;
wire _guard2042 = early_reset_static_par0_go_out;
wire _guard2043 = _guard2041 & _guard2042;
wire _guard2044 = cond_wire45_out;
wire _guard2045 = early_reset_static_par0_go_out;
wire _guard2046 = _guard2044 & _guard2045;
wire _guard2047 = cond_wire78_out;
wire _guard2048 = early_reset_static_par0_go_out;
wire _guard2049 = _guard2047 & _guard2048;
wire _guard2050 = cond_wire78_out;
wire _guard2051 = early_reset_static_par0_go_out;
wire _guard2052 = _guard2050 & _guard2051;
wire _guard2053 = cond_wire61_out;
wire _guard2054 = early_reset_static_par0_go_out;
wire _guard2055 = _guard2053 & _guard2054;
wire _guard2056 = cond_wire61_out;
wire _guard2057 = early_reset_static_par0_go_out;
wire _guard2058 = _guard2056 & _guard2057;
wire _guard2059 = cond_wire103_out;
wire _guard2060 = early_reset_static_par0_go_out;
wire _guard2061 = _guard2059 & _guard2060;
wire _guard2062 = cond_wire101_out;
wire _guard2063 = early_reset_static_par0_go_out;
wire _guard2064 = _guard2062 & _guard2063;
wire _guard2065 = fsm_out == 1'd0;
wire _guard2066 = cond_wire101_out;
wire _guard2067 = _guard2065 & _guard2066;
wire _guard2068 = fsm_out == 1'd0;
wire _guard2069 = _guard2067 & _guard2068;
wire _guard2070 = fsm_out == 1'd0;
wire _guard2071 = cond_wire103_out;
wire _guard2072 = _guard2070 & _guard2071;
wire _guard2073 = fsm_out == 1'd0;
wire _guard2074 = _guard2072 & _guard2073;
wire _guard2075 = _guard2069 | _guard2074;
wire _guard2076 = early_reset_static_par0_go_out;
wire _guard2077 = _guard2075 & _guard2076;
wire _guard2078 = fsm_out == 1'd0;
wire _guard2079 = cond_wire101_out;
wire _guard2080 = _guard2078 & _guard2079;
wire _guard2081 = fsm_out == 1'd0;
wire _guard2082 = _guard2080 & _guard2081;
wire _guard2083 = fsm_out == 1'd0;
wire _guard2084 = cond_wire103_out;
wire _guard2085 = _guard2083 & _guard2084;
wire _guard2086 = fsm_out == 1'd0;
wire _guard2087 = _guard2085 & _guard2086;
wire _guard2088 = _guard2082 | _guard2087;
wire _guard2089 = early_reset_static_par0_go_out;
wire _guard2090 = _guard2088 & _guard2089;
wire _guard2091 = fsm_out == 1'd0;
wire _guard2092 = cond_wire101_out;
wire _guard2093 = _guard2091 & _guard2092;
wire _guard2094 = fsm_out == 1'd0;
wire _guard2095 = _guard2093 & _guard2094;
wire _guard2096 = fsm_out == 1'd0;
wire _guard2097 = cond_wire103_out;
wire _guard2098 = _guard2096 & _guard2097;
wire _guard2099 = fsm_out == 1'd0;
wire _guard2100 = _guard2098 & _guard2099;
wire _guard2101 = _guard2095 | _guard2100;
wire _guard2102 = early_reset_static_par0_go_out;
wire _guard2103 = _guard2101 & _guard2102;
wire _guard2104 = cond_wire98_out;
wire _guard2105 = early_reset_static_par0_go_out;
wire _guard2106 = _guard2104 & _guard2105;
wire _guard2107 = cond_wire98_out;
wire _guard2108 = early_reset_static_par0_go_out;
wire _guard2109 = _guard2107 & _guard2108;
wire _guard2110 = cond_wire161_out;
wire _guard2111 = early_reset_static_par0_go_out;
wire _guard2112 = _guard2110 & _guard2111;
wire _guard2113 = cond_wire159_out;
wire _guard2114 = early_reset_static_par0_go_out;
wire _guard2115 = _guard2113 & _guard2114;
wire _guard2116 = fsm_out == 1'd0;
wire _guard2117 = cond_wire159_out;
wire _guard2118 = _guard2116 & _guard2117;
wire _guard2119 = fsm_out == 1'd0;
wire _guard2120 = _guard2118 & _guard2119;
wire _guard2121 = fsm_out == 1'd0;
wire _guard2122 = cond_wire161_out;
wire _guard2123 = _guard2121 & _guard2122;
wire _guard2124 = fsm_out == 1'd0;
wire _guard2125 = _guard2123 & _guard2124;
wire _guard2126 = _guard2120 | _guard2125;
wire _guard2127 = early_reset_static_par0_go_out;
wire _guard2128 = _guard2126 & _guard2127;
wire _guard2129 = fsm_out == 1'd0;
wire _guard2130 = cond_wire159_out;
wire _guard2131 = _guard2129 & _guard2130;
wire _guard2132 = fsm_out == 1'd0;
wire _guard2133 = _guard2131 & _guard2132;
wire _guard2134 = fsm_out == 1'd0;
wire _guard2135 = cond_wire161_out;
wire _guard2136 = _guard2134 & _guard2135;
wire _guard2137 = fsm_out == 1'd0;
wire _guard2138 = _guard2136 & _guard2137;
wire _guard2139 = _guard2133 | _guard2138;
wire _guard2140 = early_reset_static_par0_go_out;
wire _guard2141 = _guard2139 & _guard2140;
wire _guard2142 = fsm_out == 1'd0;
wire _guard2143 = cond_wire159_out;
wire _guard2144 = _guard2142 & _guard2143;
wire _guard2145 = fsm_out == 1'd0;
wire _guard2146 = _guard2144 & _guard2145;
wire _guard2147 = fsm_out == 1'd0;
wire _guard2148 = cond_wire161_out;
wire _guard2149 = _guard2147 & _guard2148;
wire _guard2150 = fsm_out == 1'd0;
wire _guard2151 = _guard2149 & _guard2150;
wire _guard2152 = _guard2146 | _guard2151;
wire _guard2153 = early_reset_static_par0_go_out;
wire _guard2154 = _guard2152 & _guard2153;
wire _guard2155 = cond_wire156_out;
wire _guard2156 = early_reset_static_par0_go_out;
wire _guard2157 = _guard2155 & _guard2156;
wire _guard2158 = cond_wire156_out;
wire _guard2159 = early_reset_static_par0_go_out;
wire _guard2160 = _guard2158 & _guard2159;
wire _guard2161 = cond_wire140_out;
wire _guard2162 = early_reset_static_par0_go_out;
wire _guard2163 = _guard2161 & _guard2162;
wire _guard2164 = cond_wire140_out;
wire _guard2165 = early_reset_static_par0_go_out;
wire _guard2166 = _guard2164 & _guard2165;
wire _guard2167 = cond_wire152_out;
wire _guard2168 = early_reset_static_par0_go_out;
wire _guard2169 = _guard2167 & _guard2168;
wire _guard2170 = cond_wire152_out;
wire _guard2171 = early_reset_static_par0_go_out;
wire _guard2172 = _guard2170 & _guard2171;
wire _guard2173 = cond_wire105_out;
wire _guard2174 = early_reset_static_par0_go_out;
wire _guard2175 = _guard2173 & _guard2174;
wire _guard2176 = cond_wire105_out;
wire _guard2177 = early_reset_static_par0_go_out;
wire _guard2178 = _guard2176 & _guard2177;
wire _guard2179 = early_reset_static_par0_go_out;
wire _guard2180 = early_reset_static_par0_go_out;
wire _guard2181 = early_reset_static_par0_go_out;
wire _guard2182 = early_reset_static_par0_go_out;
wire _guard2183 = early_reset_static_par0_go_out;
wire _guard2184 = early_reset_static_par0_go_out;
wire _guard2185 = early_reset_static_par_go_out;
wire _guard2186 = early_reset_static_par0_go_out;
wire _guard2187 = _guard2185 | _guard2186;
wire _guard2188 = early_reset_static_par0_go_out;
wire _guard2189 = early_reset_static_par_go_out;
wire _guard2190 = early_reset_static_par0_go_out;
wire _guard2191 = early_reset_static_par0_go_out;
wire _guard2192 = early_reset_static_par0_go_out;
wire _guard2193 = early_reset_static_par0_go_out;
wire _guard2194 = early_reset_static_par0_go_out;
wire _guard2195 = early_reset_static_par0_go_out;
wire _guard2196 = early_reset_static_par0_go_out;
wire _guard2197 = early_reset_static_par0_go_out;
wire _guard2198 = early_reset_static_par_go_out;
wire _guard2199 = early_reset_static_par0_go_out;
wire _guard2200 = _guard2198 | _guard2199;
wire _guard2201 = early_reset_static_par_go_out;
wire _guard2202 = early_reset_static_par0_go_out;
wire _guard2203 = early_reset_static_par0_go_out;
wire _guard2204 = early_reset_static_par0_go_out;
wire _guard2205 = early_reset_static_par0_go_out;
wire _guard2206 = ~_guard0;
wire _guard2207 = early_reset_static_par0_go_out;
wire _guard2208 = _guard2206 & _guard2207;
wire _guard2209 = early_reset_static_par0_go_out;
wire _guard2210 = early_reset_static_par0_go_out;
wire _guard2211 = early_reset_static_par0_go_out;
wire _guard2212 = ~_guard0;
wire _guard2213 = early_reset_static_par0_go_out;
wire _guard2214 = _guard2212 & _guard2213;
wire _guard2215 = ~_guard0;
wire _guard2216 = early_reset_static_par0_go_out;
wire _guard2217 = _guard2215 & _guard2216;
wire _guard2218 = early_reset_static_par0_go_out;
wire _guard2219 = early_reset_static_par0_go_out;
wire _guard2220 = ~_guard0;
wire _guard2221 = early_reset_static_par0_go_out;
wire _guard2222 = _guard2220 & _guard2221;
wire _guard2223 = early_reset_static_par0_go_out;
wire _guard2224 = early_reset_static_par0_go_out;
wire _guard2225 = early_reset_static_par0_go_out;
wire _guard2226 = early_reset_static_par0_go_out;
wire _guard2227 = early_reset_static_par0_go_out;
wire _guard2228 = early_reset_static_par0_go_out;
wire _guard2229 = early_reset_static_par0_go_out;
wire _guard2230 = early_reset_static_par0_go_out;
wire _guard2231 = early_reset_static_par0_go_out;
wire _guard2232 = ~_guard0;
wire _guard2233 = early_reset_static_par0_go_out;
wire _guard2234 = _guard2232 & _guard2233;
wire _guard2235 = early_reset_static_par0_go_out;
wire _guard2236 = early_reset_static_par0_go_out;
wire _guard2237 = ~_guard0;
wire _guard2238 = early_reset_static_par0_go_out;
wire _guard2239 = _guard2237 & _guard2238;
wire _guard2240 = early_reset_static_par0_go_out;
wire _guard2241 = early_reset_static_par0_go_out;
wire _guard2242 = ~_guard0;
wire _guard2243 = early_reset_static_par0_go_out;
wire _guard2244 = _guard2242 & _guard2243;
wire _guard2245 = early_reset_static_par0_go_out;
wire _guard2246 = ~_guard0;
wire _guard2247 = early_reset_static_par0_go_out;
wire _guard2248 = _guard2246 & _guard2247;
wire _guard2249 = early_reset_static_par0_go_out;
wire _guard2250 = ~_guard0;
wire _guard2251 = early_reset_static_par0_go_out;
wire _guard2252 = _guard2250 & _guard2251;
wire _guard2253 = early_reset_static_par0_go_out;
wire _guard2254 = early_reset_static_par0_go_out;
wire _guard2255 = early_reset_static_par0_go_out;
wire _guard2256 = ~_guard0;
wire _guard2257 = early_reset_static_par0_go_out;
wire _guard2258 = _guard2256 & _guard2257;
wire _guard2259 = early_reset_static_par0_go_out;
wire _guard2260 = ~_guard0;
wire _guard2261 = early_reset_static_par0_go_out;
wire _guard2262 = _guard2260 & _guard2261;
wire _guard2263 = early_reset_static_par0_go_out;
wire _guard2264 = ~_guard0;
wire _guard2265 = early_reset_static_par0_go_out;
wire _guard2266 = _guard2264 & _guard2265;
wire _guard2267 = early_reset_static_par0_go_out;
wire _guard2268 = early_reset_static_par0_go_out;
wire _guard2269 = early_reset_static_par0_go_out;
wire _guard2270 = early_reset_static_par0_go_out;
wire _guard2271 = early_reset_static_par0_go_out;
wire _guard2272 = early_reset_static_par0_go_out;
wire _guard2273 = early_reset_static_par0_go_out;
wire _guard2274 = ~_guard0;
wire _guard2275 = early_reset_static_par0_go_out;
wire _guard2276 = _guard2274 & _guard2275;
wire _guard2277 = ~_guard0;
wire _guard2278 = early_reset_static_par0_go_out;
wire _guard2279 = _guard2277 & _guard2278;
wire _guard2280 = early_reset_static_par0_go_out;
wire _guard2281 = early_reset_static_par0_go_out;
wire _guard2282 = early_reset_static_par0_go_out;
wire _guard2283 = early_reset_static_par0_go_out;
wire _guard2284 = early_reset_static_par0_go_out;
wire _guard2285 = ~_guard0;
wire _guard2286 = early_reset_static_par0_go_out;
wire _guard2287 = _guard2285 & _guard2286;
wire _guard2288 = early_reset_static_par0_go_out;
wire _guard2289 = early_reset_static_par0_go_out;
wire _guard2290 = early_reset_static_par0_go_out;
wire _guard2291 = early_reset_static_par0_go_out;
wire _guard2292 = early_reset_static_par0_go_out;
wire _guard2293 = early_reset_static_par0_go_out;
wire _guard2294 = early_reset_static_par0_go_out;
wire _guard2295 = cond_wire42_out;
wire _guard2296 = early_reset_static_par0_go_out;
wire _guard2297 = _guard2295 & _guard2296;
wire _guard2298 = cond_wire40_out;
wire _guard2299 = early_reset_static_par0_go_out;
wire _guard2300 = _guard2298 & _guard2299;
wire _guard2301 = fsm_out == 1'd0;
wire _guard2302 = cond_wire40_out;
wire _guard2303 = _guard2301 & _guard2302;
wire _guard2304 = fsm_out == 1'd0;
wire _guard2305 = _guard2303 & _guard2304;
wire _guard2306 = fsm_out == 1'd0;
wire _guard2307 = cond_wire42_out;
wire _guard2308 = _guard2306 & _guard2307;
wire _guard2309 = fsm_out == 1'd0;
wire _guard2310 = _guard2308 & _guard2309;
wire _guard2311 = _guard2305 | _guard2310;
wire _guard2312 = early_reset_static_par0_go_out;
wire _guard2313 = _guard2311 & _guard2312;
wire _guard2314 = fsm_out == 1'd0;
wire _guard2315 = cond_wire40_out;
wire _guard2316 = _guard2314 & _guard2315;
wire _guard2317 = fsm_out == 1'd0;
wire _guard2318 = _guard2316 & _guard2317;
wire _guard2319 = fsm_out == 1'd0;
wire _guard2320 = cond_wire42_out;
wire _guard2321 = _guard2319 & _guard2320;
wire _guard2322 = fsm_out == 1'd0;
wire _guard2323 = _guard2321 & _guard2322;
wire _guard2324 = _guard2318 | _guard2323;
wire _guard2325 = early_reset_static_par0_go_out;
wire _guard2326 = _guard2324 & _guard2325;
wire _guard2327 = fsm_out == 1'd0;
wire _guard2328 = cond_wire40_out;
wire _guard2329 = _guard2327 & _guard2328;
wire _guard2330 = fsm_out == 1'd0;
wire _guard2331 = _guard2329 & _guard2330;
wire _guard2332 = fsm_out == 1'd0;
wire _guard2333 = cond_wire42_out;
wire _guard2334 = _guard2332 & _guard2333;
wire _guard2335 = fsm_out == 1'd0;
wire _guard2336 = _guard2334 & _guard2335;
wire _guard2337 = _guard2331 | _guard2336;
wire _guard2338 = early_reset_static_par0_go_out;
wire _guard2339 = _guard2337 & _guard2338;
wire _guard2340 = cond_wire39_out;
wire _guard2341 = early_reset_static_par0_go_out;
wire _guard2342 = _guard2340 & _guard2341;
wire _guard2343 = cond_wire39_out;
wire _guard2344 = early_reset_static_par0_go_out;
wire _guard2345 = _guard2343 & _guard2344;
wire _guard2346 = cond_wire41_out;
wire _guard2347 = early_reset_static_par0_go_out;
wire _guard2348 = _guard2346 & _guard2347;
wire _guard2349 = cond_wire41_out;
wire _guard2350 = early_reset_static_par0_go_out;
wire _guard2351 = _guard2349 & _guard2350;
wire _guard2352 = cond_wire11_out;
wire _guard2353 = early_reset_static_par0_go_out;
wire _guard2354 = _guard2352 & _guard2353;
wire _guard2355 = cond_wire11_out;
wire _guard2356 = early_reset_static_par0_go_out;
wire _guard2357 = _guard2355 & _guard2356;
wire _guard2358 = cond_wire72_out;
wire _guard2359 = early_reset_static_par0_go_out;
wire _guard2360 = _guard2358 & _guard2359;
wire _guard2361 = cond_wire72_out;
wire _guard2362 = early_reset_static_par0_go_out;
wire _guard2363 = _guard2361 & _guard2362;
wire _guard2364 = cond_wire107_out;
wire _guard2365 = early_reset_static_par0_go_out;
wire _guard2366 = _guard2364 & _guard2365;
wire _guard2367 = cond_wire107_out;
wire _guard2368 = early_reset_static_par0_go_out;
wire _guard2369 = _guard2367 & _guard2368;
wire _guard2370 = cond_wire116_out;
wire _guard2371 = early_reset_static_par0_go_out;
wire _guard2372 = _guard2370 & _guard2371;
wire _guard2373 = cond_wire114_out;
wire _guard2374 = early_reset_static_par0_go_out;
wire _guard2375 = _guard2373 & _guard2374;
wire _guard2376 = fsm_out == 1'd0;
wire _guard2377 = cond_wire114_out;
wire _guard2378 = _guard2376 & _guard2377;
wire _guard2379 = fsm_out == 1'd0;
wire _guard2380 = _guard2378 & _guard2379;
wire _guard2381 = fsm_out == 1'd0;
wire _guard2382 = cond_wire116_out;
wire _guard2383 = _guard2381 & _guard2382;
wire _guard2384 = fsm_out == 1'd0;
wire _guard2385 = _guard2383 & _guard2384;
wire _guard2386 = _guard2380 | _guard2385;
wire _guard2387 = early_reset_static_par0_go_out;
wire _guard2388 = _guard2386 & _guard2387;
wire _guard2389 = fsm_out == 1'd0;
wire _guard2390 = cond_wire114_out;
wire _guard2391 = _guard2389 & _guard2390;
wire _guard2392 = fsm_out == 1'd0;
wire _guard2393 = _guard2391 & _guard2392;
wire _guard2394 = fsm_out == 1'd0;
wire _guard2395 = cond_wire116_out;
wire _guard2396 = _guard2394 & _guard2395;
wire _guard2397 = fsm_out == 1'd0;
wire _guard2398 = _guard2396 & _guard2397;
wire _guard2399 = _guard2393 | _guard2398;
wire _guard2400 = early_reset_static_par0_go_out;
wire _guard2401 = _guard2399 & _guard2400;
wire _guard2402 = fsm_out == 1'd0;
wire _guard2403 = cond_wire114_out;
wire _guard2404 = _guard2402 & _guard2403;
wire _guard2405 = fsm_out == 1'd0;
wire _guard2406 = _guard2404 & _guard2405;
wire _guard2407 = fsm_out == 1'd0;
wire _guard2408 = cond_wire116_out;
wire _guard2409 = _guard2407 & _guard2408;
wire _guard2410 = fsm_out == 1'd0;
wire _guard2411 = _guard2409 & _guard2410;
wire _guard2412 = _guard2406 | _guard2411;
wire _guard2413 = early_reset_static_par0_go_out;
wire _guard2414 = _guard2412 & _guard2413;
wire _guard2415 = cond_wire128_out;
wire _guard2416 = early_reset_static_par0_go_out;
wire _guard2417 = _guard2415 & _guard2416;
wire _guard2418 = cond_wire126_out;
wire _guard2419 = early_reset_static_par0_go_out;
wire _guard2420 = _guard2418 & _guard2419;
wire _guard2421 = fsm_out == 1'd0;
wire _guard2422 = cond_wire126_out;
wire _guard2423 = _guard2421 & _guard2422;
wire _guard2424 = fsm_out == 1'd0;
wire _guard2425 = _guard2423 & _guard2424;
wire _guard2426 = fsm_out == 1'd0;
wire _guard2427 = cond_wire128_out;
wire _guard2428 = _guard2426 & _guard2427;
wire _guard2429 = fsm_out == 1'd0;
wire _guard2430 = _guard2428 & _guard2429;
wire _guard2431 = _guard2425 | _guard2430;
wire _guard2432 = early_reset_static_par0_go_out;
wire _guard2433 = _guard2431 & _guard2432;
wire _guard2434 = fsm_out == 1'd0;
wire _guard2435 = cond_wire126_out;
wire _guard2436 = _guard2434 & _guard2435;
wire _guard2437 = fsm_out == 1'd0;
wire _guard2438 = _guard2436 & _guard2437;
wire _guard2439 = fsm_out == 1'd0;
wire _guard2440 = cond_wire128_out;
wire _guard2441 = _guard2439 & _guard2440;
wire _guard2442 = fsm_out == 1'd0;
wire _guard2443 = _guard2441 & _guard2442;
wire _guard2444 = _guard2438 | _guard2443;
wire _guard2445 = early_reset_static_par0_go_out;
wire _guard2446 = _guard2444 & _guard2445;
wire _guard2447 = fsm_out == 1'd0;
wire _guard2448 = cond_wire126_out;
wire _guard2449 = _guard2447 & _guard2448;
wire _guard2450 = fsm_out == 1'd0;
wire _guard2451 = _guard2449 & _guard2450;
wire _guard2452 = fsm_out == 1'd0;
wire _guard2453 = cond_wire128_out;
wire _guard2454 = _guard2452 & _guard2453;
wire _guard2455 = fsm_out == 1'd0;
wire _guard2456 = _guard2454 & _guard2455;
wire _guard2457 = _guard2451 | _guard2456;
wire _guard2458 = early_reset_static_par0_go_out;
wire _guard2459 = _guard2457 & _guard2458;
wire _guard2460 = cond_wire132_out;
wire _guard2461 = early_reset_static_par0_go_out;
wire _guard2462 = _guard2460 & _guard2461;
wire _guard2463 = cond_wire130_out;
wire _guard2464 = early_reset_static_par0_go_out;
wire _guard2465 = _guard2463 & _guard2464;
wire _guard2466 = fsm_out == 1'd0;
wire _guard2467 = cond_wire130_out;
wire _guard2468 = _guard2466 & _guard2467;
wire _guard2469 = fsm_out == 1'd0;
wire _guard2470 = _guard2468 & _guard2469;
wire _guard2471 = fsm_out == 1'd0;
wire _guard2472 = cond_wire132_out;
wire _guard2473 = _guard2471 & _guard2472;
wire _guard2474 = fsm_out == 1'd0;
wire _guard2475 = _guard2473 & _guard2474;
wire _guard2476 = _guard2470 | _guard2475;
wire _guard2477 = early_reset_static_par0_go_out;
wire _guard2478 = _guard2476 & _guard2477;
wire _guard2479 = fsm_out == 1'd0;
wire _guard2480 = cond_wire130_out;
wire _guard2481 = _guard2479 & _guard2480;
wire _guard2482 = fsm_out == 1'd0;
wire _guard2483 = _guard2481 & _guard2482;
wire _guard2484 = fsm_out == 1'd0;
wire _guard2485 = cond_wire132_out;
wire _guard2486 = _guard2484 & _guard2485;
wire _guard2487 = fsm_out == 1'd0;
wire _guard2488 = _guard2486 & _guard2487;
wire _guard2489 = _guard2483 | _guard2488;
wire _guard2490 = early_reset_static_par0_go_out;
wire _guard2491 = _guard2489 & _guard2490;
wire _guard2492 = fsm_out == 1'd0;
wire _guard2493 = cond_wire130_out;
wire _guard2494 = _guard2492 & _guard2493;
wire _guard2495 = fsm_out == 1'd0;
wire _guard2496 = _guard2494 & _guard2495;
wire _guard2497 = fsm_out == 1'd0;
wire _guard2498 = cond_wire132_out;
wire _guard2499 = _guard2497 & _guard2498;
wire _guard2500 = fsm_out == 1'd0;
wire _guard2501 = _guard2499 & _guard2500;
wire _guard2502 = _guard2496 | _guard2501;
wire _guard2503 = early_reset_static_par0_go_out;
wire _guard2504 = _guard2502 & _guard2503;
wire _guard2505 = cond_wire131_out;
wire _guard2506 = early_reset_static_par0_go_out;
wire _guard2507 = _guard2505 & _guard2506;
wire _guard2508 = cond_wire131_out;
wire _guard2509 = early_reset_static_par0_go_out;
wire _guard2510 = _guard2508 & _guard2509;
wire _guard2511 = cond_wire127_out;
wire _guard2512 = early_reset_static_par0_go_out;
wire _guard2513 = _guard2511 & _guard2512;
wire _guard2514 = cond_wire127_out;
wire _guard2515 = early_reset_static_par0_go_out;
wire _guard2516 = _guard2514 & _guard2515;
wire _guard2517 = cond_wire190_out;
wire _guard2518 = early_reset_static_par0_go_out;
wire _guard2519 = _guard2517 & _guard2518;
wire _guard2520 = cond_wire188_out;
wire _guard2521 = early_reset_static_par0_go_out;
wire _guard2522 = _guard2520 & _guard2521;
wire _guard2523 = fsm_out == 1'd0;
wire _guard2524 = cond_wire188_out;
wire _guard2525 = _guard2523 & _guard2524;
wire _guard2526 = fsm_out == 1'd0;
wire _guard2527 = _guard2525 & _guard2526;
wire _guard2528 = fsm_out == 1'd0;
wire _guard2529 = cond_wire190_out;
wire _guard2530 = _guard2528 & _guard2529;
wire _guard2531 = fsm_out == 1'd0;
wire _guard2532 = _guard2530 & _guard2531;
wire _guard2533 = _guard2527 | _guard2532;
wire _guard2534 = early_reset_static_par0_go_out;
wire _guard2535 = _guard2533 & _guard2534;
wire _guard2536 = fsm_out == 1'd0;
wire _guard2537 = cond_wire188_out;
wire _guard2538 = _guard2536 & _guard2537;
wire _guard2539 = fsm_out == 1'd0;
wire _guard2540 = _guard2538 & _guard2539;
wire _guard2541 = fsm_out == 1'd0;
wire _guard2542 = cond_wire190_out;
wire _guard2543 = _guard2541 & _guard2542;
wire _guard2544 = fsm_out == 1'd0;
wire _guard2545 = _guard2543 & _guard2544;
wire _guard2546 = _guard2540 | _guard2545;
wire _guard2547 = early_reset_static_par0_go_out;
wire _guard2548 = _guard2546 & _guard2547;
wire _guard2549 = fsm_out == 1'd0;
wire _guard2550 = cond_wire188_out;
wire _guard2551 = _guard2549 & _guard2550;
wire _guard2552 = fsm_out == 1'd0;
wire _guard2553 = _guard2551 & _guard2552;
wire _guard2554 = fsm_out == 1'd0;
wire _guard2555 = cond_wire190_out;
wire _guard2556 = _guard2554 & _guard2555;
wire _guard2557 = fsm_out == 1'd0;
wire _guard2558 = _guard2556 & _guard2557;
wire _guard2559 = _guard2553 | _guard2558;
wire _guard2560 = early_reset_static_par0_go_out;
wire _guard2561 = _guard2559 & _guard2560;
wire _guard2562 = cond_wire214_out;
wire _guard2563 = early_reset_static_par0_go_out;
wire _guard2564 = _guard2562 & _guard2563;
wire _guard2565 = cond_wire214_out;
wire _guard2566 = early_reset_static_par0_go_out;
wire _guard2567 = _guard2565 & _guard2566;
wire _guard2568 = cond_wire256_out;
wire _guard2569 = early_reset_static_par0_go_out;
wire _guard2570 = _guard2568 & _guard2569;
wire _guard2571 = cond_wire254_out;
wire _guard2572 = early_reset_static_par0_go_out;
wire _guard2573 = _guard2571 & _guard2572;
wire _guard2574 = fsm_out == 1'd0;
wire _guard2575 = cond_wire254_out;
wire _guard2576 = _guard2574 & _guard2575;
wire _guard2577 = fsm_out == 1'd0;
wire _guard2578 = _guard2576 & _guard2577;
wire _guard2579 = fsm_out == 1'd0;
wire _guard2580 = cond_wire256_out;
wire _guard2581 = _guard2579 & _guard2580;
wire _guard2582 = fsm_out == 1'd0;
wire _guard2583 = _guard2581 & _guard2582;
wire _guard2584 = _guard2578 | _guard2583;
wire _guard2585 = early_reset_static_par0_go_out;
wire _guard2586 = _guard2584 & _guard2585;
wire _guard2587 = fsm_out == 1'd0;
wire _guard2588 = cond_wire254_out;
wire _guard2589 = _guard2587 & _guard2588;
wire _guard2590 = fsm_out == 1'd0;
wire _guard2591 = _guard2589 & _guard2590;
wire _guard2592 = fsm_out == 1'd0;
wire _guard2593 = cond_wire256_out;
wire _guard2594 = _guard2592 & _guard2593;
wire _guard2595 = fsm_out == 1'd0;
wire _guard2596 = _guard2594 & _guard2595;
wire _guard2597 = _guard2591 | _guard2596;
wire _guard2598 = early_reset_static_par0_go_out;
wire _guard2599 = _guard2597 & _guard2598;
wire _guard2600 = fsm_out == 1'd0;
wire _guard2601 = cond_wire254_out;
wire _guard2602 = _guard2600 & _guard2601;
wire _guard2603 = fsm_out == 1'd0;
wire _guard2604 = _guard2602 & _guard2603;
wire _guard2605 = fsm_out == 1'd0;
wire _guard2606 = cond_wire256_out;
wire _guard2607 = _guard2605 & _guard2606;
wire _guard2608 = fsm_out == 1'd0;
wire _guard2609 = _guard2607 & _guard2608;
wire _guard2610 = _guard2604 | _guard2609;
wire _guard2611 = early_reset_static_par0_go_out;
wire _guard2612 = _guard2610 & _guard2611;
wire _guard2613 = early_reset_static_par_go_out;
wire _guard2614 = cond_wire4_out;
wire _guard2615 = early_reset_static_par0_go_out;
wire _guard2616 = _guard2614 & _guard2615;
wire _guard2617 = _guard2613 | _guard2616;
wire _guard2618 = early_reset_static_par_go_out;
wire _guard2619 = cond_wire4_out;
wire _guard2620 = early_reset_static_par0_go_out;
wire _guard2621 = _guard2619 & _guard2620;
wire _guard2622 = early_reset_static_par_go_out;
wire _guard2623 = cond_wire34_out;
wire _guard2624 = early_reset_static_par0_go_out;
wire _guard2625 = _guard2623 & _guard2624;
wire _guard2626 = _guard2622 | _guard2625;
wire _guard2627 = early_reset_static_par_go_out;
wire _guard2628 = cond_wire34_out;
wire _guard2629 = early_reset_static_par0_go_out;
wire _guard2630 = _guard2628 & _guard2629;
wire _guard2631 = early_reset_static_par0_go_out;
wire _guard2632 = early_reset_static_par0_go_out;
wire _guard2633 = early_reset_static_par0_go_out;
wire _guard2634 = early_reset_static_par0_go_out;
wire _guard2635 = early_reset_static_par0_go_out;
wire _guard2636 = early_reset_static_par0_go_out;
wire _guard2637 = early_reset_static_par0_go_out;
wire _guard2638 = early_reset_static_par0_go_out;
wire _guard2639 = early_reset_static_par_go_out;
wire _guard2640 = early_reset_static_par0_go_out;
wire _guard2641 = _guard2639 | _guard2640;
wire _guard2642 = early_reset_static_par_go_out;
wire _guard2643 = early_reset_static_par0_go_out;
wire _guard2644 = early_reset_static_par0_go_out;
wire _guard2645 = early_reset_static_par0_go_out;
wire _guard2646 = early_reset_static_par0_go_out;
wire _guard2647 = early_reset_static_par0_go_out;
wire _guard2648 = early_reset_static_par0_go_out;
wire _guard2649 = early_reset_static_par0_go_out;
wire _guard2650 = early_reset_static_par0_go_out;
wire _guard2651 = early_reset_static_par0_go_out;
wire _guard2652 = early_reset_static_par0_go_out;
wire _guard2653 = early_reset_static_par0_go_out;
wire _guard2654 = ~_guard0;
wire _guard2655 = early_reset_static_par0_go_out;
wire _guard2656 = _guard2654 & _guard2655;
wire _guard2657 = early_reset_static_par0_go_out;
wire _guard2658 = early_reset_static_par0_go_out;
wire _guard2659 = ~_guard0;
wire _guard2660 = early_reset_static_par0_go_out;
wire _guard2661 = _guard2659 & _guard2660;
wire _guard2662 = early_reset_static_par0_go_out;
wire _guard2663 = ~_guard0;
wire _guard2664 = early_reset_static_par0_go_out;
wire _guard2665 = _guard2663 & _guard2664;
wire _guard2666 = ~_guard0;
wire _guard2667 = early_reset_static_par0_go_out;
wire _guard2668 = _guard2666 & _guard2667;
wire _guard2669 = early_reset_static_par0_go_out;
wire _guard2670 = ~_guard0;
wire _guard2671 = early_reset_static_par0_go_out;
wire _guard2672 = _guard2670 & _guard2671;
wire _guard2673 = early_reset_static_par0_go_out;
wire _guard2674 = ~_guard0;
wire _guard2675 = early_reset_static_par0_go_out;
wire _guard2676 = _guard2674 & _guard2675;
wire _guard2677 = early_reset_static_par0_go_out;
wire _guard2678 = ~_guard0;
wire _guard2679 = early_reset_static_par0_go_out;
wire _guard2680 = _guard2678 & _guard2679;
wire _guard2681 = early_reset_static_par0_go_out;
wire _guard2682 = early_reset_static_par0_go_out;
wire _guard2683 = early_reset_static_par0_go_out;
wire _guard2684 = early_reset_static_par0_go_out;
wire _guard2685 = ~_guard0;
wire _guard2686 = early_reset_static_par0_go_out;
wire _guard2687 = _guard2685 & _guard2686;
wire _guard2688 = early_reset_static_par0_go_out;
wire _guard2689 = early_reset_static_par0_go_out;
wire _guard2690 = ~_guard0;
wire _guard2691 = early_reset_static_par0_go_out;
wire _guard2692 = _guard2690 & _guard2691;
wire _guard2693 = early_reset_static_par0_go_out;
wire _guard2694 = early_reset_static_par0_go_out;
wire _guard2695 = early_reset_static_par0_go_out;
wire _guard2696 = early_reset_static_par0_go_out;
wire _guard2697 = ~_guard0;
wire _guard2698 = early_reset_static_par0_go_out;
wire _guard2699 = _guard2697 & _guard2698;
wire _guard2700 = ~_guard0;
wire _guard2701 = early_reset_static_par0_go_out;
wire _guard2702 = _guard2700 & _guard2701;
wire _guard2703 = early_reset_static_par0_go_out;
wire _guard2704 = ~_guard0;
wire _guard2705 = early_reset_static_par0_go_out;
wire _guard2706 = _guard2704 & _guard2705;
wire _guard2707 = early_reset_static_par0_go_out;
wire _guard2708 = early_reset_static_par0_go_out;
wire _guard2709 = early_reset_static_par0_go_out;
wire _guard2710 = early_reset_static_par0_go_out;
wire _guard2711 = early_reset_static_par0_go_out;
wire _guard2712 = ~_guard0;
wire _guard2713 = early_reset_static_par0_go_out;
wire _guard2714 = _guard2712 & _guard2713;
wire _guard2715 = early_reset_static_par0_go_out;
wire _guard2716 = early_reset_static_par0_go_out;
wire _guard2717 = ~_guard0;
wire _guard2718 = early_reset_static_par0_go_out;
wire _guard2719 = _guard2717 & _guard2718;
wire _guard2720 = early_reset_static_par0_go_out;
wire _guard2721 = early_reset_static_par0_go_out;
wire _guard2722 = early_reset_static_par0_go_out;
wire _guard2723 = early_reset_static_par0_go_out;
wire _guard2724 = ~_guard0;
wire _guard2725 = early_reset_static_par0_go_out;
wire _guard2726 = _guard2724 & _guard2725;
wire _guard2727 = early_reset_static_par0_go_out;
wire _guard2728 = ~_guard0;
wire _guard2729 = early_reset_static_par0_go_out;
wire _guard2730 = _guard2728 & _guard2729;
wire _guard2731 = early_reset_static_par0_go_out;
wire _guard2732 = early_reset_static_par0_go_out;
wire _guard2733 = early_reset_static_par0_go_out;
wire _guard2734 = ~_guard0;
wire _guard2735 = early_reset_static_par0_go_out;
wire _guard2736 = _guard2734 & _guard2735;
wire _guard2737 = early_reset_static_par0_go_out;
wire _guard2738 = early_reset_static_par0_go_out;
wire _guard2739 = early_reset_static_par0_go_out;
wire _guard2740 = early_reset_static_par0_go_out;
wire _guard2741 = early_reset_static_par0_go_out;
wire _guard2742 = early_reset_static_par0_go_out;
wire _guard2743 = early_reset_static_par0_go_out;
wire _guard2744 = early_reset_static_par0_go_out;
wire _guard2745 = early_reset_static_par0_go_out;
wire _guard2746 = early_reset_static_par0_go_out;
wire _guard2747 = early_reset_static_par0_go_out;
wire _guard2748 = early_reset_static_par0_go_out;
wire _guard2749 = early_reset_static_par0_go_out;
wire _guard2750 = cond_wire_out;
wire _guard2751 = early_reset_static_par0_go_out;
wire _guard2752 = _guard2750 & _guard2751;
wire _guard2753 = cond_wire_out;
wire _guard2754 = early_reset_static_par0_go_out;
wire _guard2755 = _guard2753 & _guard2754;
wire _guard2756 = cond_wire17_out;
wire _guard2757 = early_reset_static_par0_go_out;
wire _guard2758 = _guard2756 & _guard2757;
wire _guard2759 = cond_wire15_out;
wire _guard2760 = early_reset_static_par0_go_out;
wire _guard2761 = _guard2759 & _guard2760;
wire _guard2762 = fsm_out == 1'd0;
wire _guard2763 = cond_wire15_out;
wire _guard2764 = _guard2762 & _guard2763;
wire _guard2765 = fsm_out == 1'd0;
wire _guard2766 = _guard2764 & _guard2765;
wire _guard2767 = fsm_out == 1'd0;
wire _guard2768 = cond_wire17_out;
wire _guard2769 = _guard2767 & _guard2768;
wire _guard2770 = fsm_out == 1'd0;
wire _guard2771 = _guard2769 & _guard2770;
wire _guard2772 = _guard2766 | _guard2771;
wire _guard2773 = early_reset_static_par0_go_out;
wire _guard2774 = _guard2772 & _guard2773;
wire _guard2775 = fsm_out == 1'd0;
wire _guard2776 = cond_wire15_out;
wire _guard2777 = _guard2775 & _guard2776;
wire _guard2778 = fsm_out == 1'd0;
wire _guard2779 = _guard2777 & _guard2778;
wire _guard2780 = fsm_out == 1'd0;
wire _guard2781 = cond_wire17_out;
wire _guard2782 = _guard2780 & _guard2781;
wire _guard2783 = fsm_out == 1'd0;
wire _guard2784 = _guard2782 & _guard2783;
wire _guard2785 = _guard2779 | _guard2784;
wire _guard2786 = early_reset_static_par0_go_out;
wire _guard2787 = _guard2785 & _guard2786;
wire _guard2788 = fsm_out == 1'd0;
wire _guard2789 = cond_wire15_out;
wire _guard2790 = _guard2788 & _guard2789;
wire _guard2791 = fsm_out == 1'd0;
wire _guard2792 = _guard2790 & _guard2791;
wire _guard2793 = fsm_out == 1'd0;
wire _guard2794 = cond_wire17_out;
wire _guard2795 = _guard2793 & _guard2794;
wire _guard2796 = fsm_out == 1'd0;
wire _guard2797 = _guard2795 & _guard2796;
wire _guard2798 = _guard2792 | _guard2797;
wire _guard2799 = early_reset_static_par0_go_out;
wire _guard2800 = _guard2798 & _guard2799;
wire _guard2801 = cond_wire27_out;
wire _guard2802 = early_reset_static_par0_go_out;
wire _guard2803 = _guard2801 & _guard2802;
wire _guard2804 = cond_wire25_out;
wire _guard2805 = early_reset_static_par0_go_out;
wire _guard2806 = _guard2804 & _guard2805;
wire _guard2807 = fsm_out == 1'd0;
wire _guard2808 = cond_wire25_out;
wire _guard2809 = _guard2807 & _guard2808;
wire _guard2810 = fsm_out == 1'd0;
wire _guard2811 = _guard2809 & _guard2810;
wire _guard2812 = fsm_out == 1'd0;
wire _guard2813 = cond_wire27_out;
wire _guard2814 = _guard2812 & _guard2813;
wire _guard2815 = fsm_out == 1'd0;
wire _guard2816 = _guard2814 & _guard2815;
wire _guard2817 = _guard2811 | _guard2816;
wire _guard2818 = early_reset_static_par0_go_out;
wire _guard2819 = _guard2817 & _guard2818;
wire _guard2820 = fsm_out == 1'd0;
wire _guard2821 = cond_wire25_out;
wire _guard2822 = _guard2820 & _guard2821;
wire _guard2823 = fsm_out == 1'd0;
wire _guard2824 = _guard2822 & _guard2823;
wire _guard2825 = fsm_out == 1'd0;
wire _guard2826 = cond_wire27_out;
wire _guard2827 = _guard2825 & _guard2826;
wire _guard2828 = fsm_out == 1'd0;
wire _guard2829 = _guard2827 & _guard2828;
wire _guard2830 = _guard2824 | _guard2829;
wire _guard2831 = early_reset_static_par0_go_out;
wire _guard2832 = _guard2830 & _guard2831;
wire _guard2833 = fsm_out == 1'd0;
wire _guard2834 = cond_wire25_out;
wire _guard2835 = _guard2833 & _guard2834;
wire _guard2836 = fsm_out == 1'd0;
wire _guard2837 = _guard2835 & _guard2836;
wire _guard2838 = fsm_out == 1'd0;
wire _guard2839 = cond_wire27_out;
wire _guard2840 = _guard2838 & _guard2839;
wire _guard2841 = fsm_out == 1'd0;
wire _guard2842 = _guard2840 & _guard2841;
wire _guard2843 = _guard2837 | _guard2842;
wire _guard2844 = early_reset_static_par0_go_out;
wire _guard2845 = _guard2843 & _guard2844;
wire _guard2846 = cond_wire16_out;
wire _guard2847 = early_reset_static_par0_go_out;
wire _guard2848 = _guard2846 & _guard2847;
wire _guard2849 = cond_wire16_out;
wire _guard2850 = early_reset_static_par0_go_out;
wire _guard2851 = _guard2849 & _guard2850;
wire _guard2852 = cond_wire21_out;
wire _guard2853 = early_reset_static_par0_go_out;
wire _guard2854 = _guard2852 & _guard2853;
wire _guard2855 = cond_wire21_out;
wire _guard2856 = early_reset_static_par0_go_out;
wire _guard2857 = _guard2855 & _guard2856;
wire _guard2858 = cond_wire82_out;
wire _guard2859 = early_reset_static_par0_go_out;
wire _guard2860 = _guard2858 & _guard2859;
wire _guard2861 = cond_wire82_out;
wire _guard2862 = early_reset_static_par0_go_out;
wire _guard2863 = _guard2861 & _guard2862;
wire _guard2864 = cond_wire91_out;
wire _guard2865 = early_reset_static_par0_go_out;
wire _guard2866 = _guard2864 & _guard2865;
wire _guard2867 = cond_wire89_out;
wire _guard2868 = early_reset_static_par0_go_out;
wire _guard2869 = _guard2867 & _guard2868;
wire _guard2870 = fsm_out == 1'd0;
wire _guard2871 = cond_wire89_out;
wire _guard2872 = _guard2870 & _guard2871;
wire _guard2873 = fsm_out == 1'd0;
wire _guard2874 = _guard2872 & _guard2873;
wire _guard2875 = fsm_out == 1'd0;
wire _guard2876 = cond_wire91_out;
wire _guard2877 = _guard2875 & _guard2876;
wire _guard2878 = fsm_out == 1'd0;
wire _guard2879 = _guard2877 & _guard2878;
wire _guard2880 = _guard2874 | _guard2879;
wire _guard2881 = early_reset_static_par0_go_out;
wire _guard2882 = _guard2880 & _guard2881;
wire _guard2883 = fsm_out == 1'd0;
wire _guard2884 = cond_wire89_out;
wire _guard2885 = _guard2883 & _guard2884;
wire _guard2886 = fsm_out == 1'd0;
wire _guard2887 = _guard2885 & _guard2886;
wire _guard2888 = fsm_out == 1'd0;
wire _guard2889 = cond_wire91_out;
wire _guard2890 = _guard2888 & _guard2889;
wire _guard2891 = fsm_out == 1'd0;
wire _guard2892 = _guard2890 & _guard2891;
wire _guard2893 = _guard2887 | _guard2892;
wire _guard2894 = early_reset_static_par0_go_out;
wire _guard2895 = _guard2893 & _guard2894;
wire _guard2896 = fsm_out == 1'd0;
wire _guard2897 = cond_wire89_out;
wire _guard2898 = _guard2896 & _guard2897;
wire _guard2899 = fsm_out == 1'd0;
wire _guard2900 = _guard2898 & _guard2899;
wire _guard2901 = fsm_out == 1'd0;
wire _guard2902 = cond_wire91_out;
wire _guard2903 = _guard2901 & _guard2902;
wire _guard2904 = fsm_out == 1'd0;
wire _guard2905 = _guard2903 & _guard2904;
wire _guard2906 = _guard2900 | _guard2905;
wire _guard2907 = early_reset_static_par0_go_out;
wire _guard2908 = _guard2906 & _guard2907;
wire _guard2909 = cond_wire65_out;
wire _guard2910 = early_reset_static_par0_go_out;
wire _guard2911 = _guard2909 & _guard2910;
wire _guard2912 = cond_wire65_out;
wire _guard2913 = early_reset_static_par0_go_out;
wire _guard2914 = _guard2912 & _guard2913;
wire _guard2915 = cond_wire108_out;
wire _guard2916 = early_reset_static_par0_go_out;
wire _guard2917 = _guard2915 & _guard2916;
wire _guard2918 = cond_wire106_out;
wire _guard2919 = early_reset_static_par0_go_out;
wire _guard2920 = _guard2918 & _guard2919;
wire _guard2921 = fsm_out == 1'd0;
wire _guard2922 = cond_wire106_out;
wire _guard2923 = _guard2921 & _guard2922;
wire _guard2924 = fsm_out == 1'd0;
wire _guard2925 = _guard2923 & _guard2924;
wire _guard2926 = fsm_out == 1'd0;
wire _guard2927 = cond_wire108_out;
wire _guard2928 = _guard2926 & _guard2927;
wire _guard2929 = fsm_out == 1'd0;
wire _guard2930 = _guard2928 & _guard2929;
wire _guard2931 = _guard2925 | _guard2930;
wire _guard2932 = early_reset_static_par0_go_out;
wire _guard2933 = _guard2931 & _guard2932;
wire _guard2934 = fsm_out == 1'd0;
wire _guard2935 = cond_wire106_out;
wire _guard2936 = _guard2934 & _guard2935;
wire _guard2937 = fsm_out == 1'd0;
wire _guard2938 = _guard2936 & _guard2937;
wire _guard2939 = fsm_out == 1'd0;
wire _guard2940 = cond_wire108_out;
wire _guard2941 = _guard2939 & _guard2940;
wire _guard2942 = fsm_out == 1'd0;
wire _guard2943 = _guard2941 & _guard2942;
wire _guard2944 = _guard2938 | _guard2943;
wire _guard2945 = early_reset_static_par0_go_out;
wire _guard2946 = _guard2944 & _guard2945;
wire _guard2947 = fsm_out == 1'd0;
wire _guard2948 = cond_wire106_out;
wire _guard2949 = _guard2947 & _guard2948;
wire _guard2950 = fsm_out == 1'd0;
wire _guard2951 = _guard2949 & _guard2950;
wire _guard2952 = fsm_out == 1'd0;
wire _guard2953 = cond_wire108_out;
wire _guard2954 = _guard2952 & _guard2953;
wire _guard2955 = fsm_out == 1'd0;
wire _guard2956 = _guard2954 & _guard2955;
wire _guard2957 = _guard2951 | _guard2956;
wire _guard2958 = early_reset_static_par0_go_out;
wire _guard2959 = _guard2957 & _guard2958;
wire _guard2960 = cond_wire82_out;
wire _guard2961 = early_reset_static_par0_go_out;
wire _guard2962 = _guard2960 & _guard2961;
wire _guard2963 = cond_wire82_out;
wire _guard2964 = early_reset_static_par0_go_out;
wire _guard2965 = _guard2963 & _guard2964;
wire _guard2966 = cond_wire107_out;
wire _guard2967 = early_reset_static_par0_go_out;
wire _guard2968 = _guard2966 & _guard2967;
wire _guard2969 = cond_wire107_out;
wire _guard2970 = early_reset_static_par0_go_out;
wire _guard2971 = _guard2969 & _guard2970;
wire _guard2972 = cond_wire160_out;
wire _guard2973 = early_reset_static_par0_go_out;
wire _guard2974 = _guard2972 & _guard2973;
wire _guard2975 = cond_wire160_out;
wire _guard2976 = early_reset_static_par0_go_out;
wire _guard2977 = _guard2975 & _guard2976;
wire _guard2978 = cond_wire164_out;
wire _guard2979 = early_reset_static_par0_go_out;
wire _guard2980 = _guard2978 & _guard2979;
wire _guard2981 = cond_wire164_out;
wire _guard2982 = early_reset_static_par0_go_out;
wire _guard2983 = _guard2981 & _guard2982;
wire _guard2984 = cond_wire178_out;
wire _guard2985 = early_reset_static_par0_go_out;
wire _guard2986 = _guard2984 & _guard2985;
wire _guard2987 = cond_wire176_out;
wire _guard2988 = early_reset_static_par0_go_out;
wire _guard2989 = _guard2987 & _guard2988;
wire _guard2990 = fsm_out == 1'd0;
wire _guard2991 = cond_wire176_out;
wire _guard2992 = _guard2990 & _guard2991;
wire _guard2993 = fsm_out == 1'd0;
wire _guard2994 = _guard2992 & _guard2993;
wire _guard2995 = fsm_out == 1'd0;
wire _guard2996 = cond_wire178_out;
wire _guard2997 = _guard2995 & _guard2996;
wire _guard2998 = fsm_out == 1'd0;
wire _guard2999 = _guard2997 & _guard2998;
wire _guard3000 = _guard2994 | _guard2999;
wire _guard3001 = early_reset_static_par0_go_out;
wire _guard3002 = _guard3000 & _guard3001;
wire _guard3003 = fsm_out == 1'd0;
wire _guard3004 = cond_wire176_out;
wire _guard3005 = _guard3003 & _guard3004;
wire _guard3006 = fsm_out == 1'd0;
wire _guard3007 = _guard3005 & _guard3006;
wire _guard3008 = fsm_out == 1'd0;
wire _guard3009 = cond_wire178_out;
wire _guard3010 = _guard3008 & _guard3009;
wire _guard3011 = fsm_out == 1'd0;
wire _guard3012 = _guard3010 & _guard3011;
wire _guard3013 = _guard3007 | _guard3012;
wire _guard3014 = early_reset_static_par0_go_out;
wire _guard3015 = _guard3013 & _guard3014;
wire _guard3016 = fsm_out == 1'd0;
wire _guard3017 = cond_wire176_out;
wire _guard3018 = _guard3016 & _guard3017;
wire _guard3019 = fsm_out == 1'd0;
wire _guard3020 = _guard3018 & _guard3019;
wire _guard3021 = fsm_out == 1'd0;
wire _guard3022 = cond_wire178_out;
wire _guard3023 = _guard3021 & _guard3022;
wire _guard3024 = fsm_out == 1'd0;
wire _guard3025 = _guard3023 & _guard3024;
wire _guard3026 = _guard3020 | _guard3025;
wire _guard3027 = early_reset_static_par0_go_out;
wire _guard3028 = _guard3026 & _guard3027;
wire _guard3029 = cond_wire202_out;
wire _guard3030 = early_reset_static_par0_go_out;
wire _guard3031 = _guard3029 & _guard3030;
wire _guard3032 = cond_wire200_out;
wire _guard3033 = early_reset_static_par0_go_out;
wire _guard3034 = _guard3032 & _guard3033;
wire _guard3035 = fsm_out == 1'd0;
wire _guard3036 = cond_wire200_out;
wire _guard3037 = _guard3035 & _guard3036;
wire _guard3038 = fsm_out == 1'd0;
wire _guard3039 = _guard3037 & _guard3038;
wire _guard3040 = fsm_out == 1'd0;
wire _guard3041 = cond_wire202_out;
wire _guard3042 = _guard3040 & _guard3041;
wire _guard3043 = fsm_out == 1'd0;
wire _guard3044 = _guard3042 & _guard3043;
wire _guard3045 = _guard3039 | _guard3044;
wire _guard3046 = early_reset_static_par0_go_out;
wire _guard3047 = _guard3045 & _guard3046;
wire _guard3048 = fsm_out == 1'd0;
wire _guard3049 = cond_wire200_out;
wire _guard3050 = _guard3048 & _guard3049;
wire _guard3051 = fsm_out == 1'd0;
wire _guard3052 = _guard3050 & _guard3051;
wire _guard3053 = fsm_out == 1'd0;
wire _guard3054 = cond_wire202_out;
wire _guard3055 = _guard3053 & _guard3054;
wire _guard3056 = fsm_out == 1'd0;
wire _guard3057 = _guard3055 & _guard3056;
wire _guard3058 = _guard3052 | _guard3057;
wire _guard3059 = early_reset_static_par0_go_out;
wire _guard3060 = _guard3058 & _guard3059;
wire _guard3061 = fsm_out == 1'd0;
wire _guard3062 = cond_wire200_out;
wire _guard3063 = _guard3061 & _guard3062;
wire _guard3064 = fsm_out == 1'd0;
wire _guard3065 = _guard3063 & _guard3064;
wire _guard3066 = fsm_out == 1'd0;
wire _guard3067 = cond_wire202_out;
wire _guard3068 = _guard3066 & _guard3067;
wire _guard3069 = fsm_out == 1'd0;
wire _guard3070 = _guard3068 & _guard3069;
wire _guard3071 = _guard3065 | _guard3070;
wire _guard3072 = early_reset_static_par0_go_out;
wire _guard3073 = _guard3071 & _guard3072;
wire _guard3074 = cond_wire207_out;
wire _guard3075 = early_reset_static_par0_go_out;
wire _guard3076 = _guard3074 & _guard3075;
wire _guard3077 = cond_wire205_out;
wire _guard3078 = early_reset_static_par0_go_out;
wire _guard3079 = _guard3077 & _guard3078;
wire _guard3080 = fsm_out == 1'd0;
wire _guard3081 = cond_wire205_out;
wire _guard3082 = _guard3080 & _guard3081;
wire _guard3083 = fsm_out == 1'd0;
wire _guard3084 = _guard3082 & _guard3083;
wire _guard3085 = fsm_out == 1'd0;
wire _guard3086 = cond_wire207_out;
wire _guard3087 = _guard3085 & _guard3086;
wire _guard3088 = fsm_out == 1'd0;
wire _guard3089 = _guard3087 & _guard3088;
wire _guard3090 = _guard3084 | _guard3089;
wire _guard3091 = early_reset_static_par0_go_out;
wire _guard3092 = _guard3090 & _guard3091;
wire _guard3093 = fsm_out == 1'd0;
wire _guard3094 = cond_wire205_out;
wire _guard3095 = _guard3093 & _guard3094;
wire _guard3096 = fsm_out == 1'd0;
wire _guard3097 = _guard3095 & _guard3096;
wire _guard3098 = fsm_out == 1'd0;
wire _guard3099 = cond_wire207_out;
wire _guard3100 = _guard3098 & _guard3099;
wire _guard3101 = fsm_out == 1'd0;
wire _guard3102 = _guard3100 & _guard3101;
wire _guard3103 = _guard3097 | _guard3102;
wire _guard3104 = early_reset_static_par0_go_out;
wire _guard3105 = _guard3103 & _guard3104;
wire _guard3106 = fsm_out == 1'd0;
wire _guard3107 = cond_wire205_out;
wire _guard3108 = _guard3106 & _guard3107;
wire _guard3109 = fsm_out == 1'd0;
wire _guard3110 = _guard3108 & _guard3109;
wire _guard3111 = fsm_out == 1'd0;
wire _guard3112 = cond_wire207_out;
wire _guard3113 = _guard3111 & _guard3112;
wire _guard3114 = fsm_out == 1'd0;
wire _guard3115 = _guard3113 & _guard3114;
wire _guard3116 = _guard3110 | _guard3115;
wire _guard3117 = early_reset_static_par0_go_out;
wire _guard3118 = _guard3116 & _guard3117;
wire _guard3119 = cond_wire173_out;
wire _guard3120 = early_reset_static_par0_go_out;
wire _guard3121 = _guard3119 & _guard3120;
wire _guard3122 = cond_wire173_out;
wire _guard3123 = early_reset_static_par0_go_out;
wire _guard3124 = _guard3122 & _guard3123;
wire _guard3125 = cond_wire211_out;
wire _guard3126 = early_reset_static_par0_go_out;
wire _guard3127 = _guard3125 & _guard3126;
wire _guard3128 = cond_wire209_out;
wire _guard3129 = early_reset_static_par0_go_out;
wire _guard3130 = _guard3128 & _guard3129;
wire _guard3131 = fsm_out == 1'd0;
wire _guard3132 = cond_wire209_out;
wire _guard3133 = _guard3131 & _guard3132;
wire _guard3134 = fsm_out == 1'd0;
wire _guard3135 = _guard3133 & _guard3134;
wire _guard3136 = fsm_out == 1'd0;
wire _guard3137 = cond_wire211_out;
wire _guard3138 = _guard3136 & _guard3137;
wire _guard3139 = fsm_out == 1'd0;
wire _guard3140 = _guard3138 & _guard3139;
wire _guard3141 = _guard3135 | _guard3140;
wire _guard3142 = early_reset_static_par0_go_out;
wire _guard3143 = _guard3141 & _guard3142;
wire _guard3144 = fsm_out == 1'd0;
wire _guard3145 = cond_wire209_out;
wire _guard3146 = _guard3144 & _guard3145;
wire _guard3147 = fsm_out == 1'd0;
wire _guard3148 = _guard3146 & _guard3147;
wire _guard3149 = fsm_out == 1'd0;
wire _guard3150 = cond_wire211_out;
wire _guard3151 = _guard3149 & _guard3150;
wire _guard3152 = fsm_out == 1'd0;
wire _guard3153 = _guard3151 & _guard3152;
wire _guard3154 = _guard3148 | _guard3153;
wire _guard3155 = early_reset_static_par0_go_out;
wire _guard3156 = _guard3154 & _guard3155;
wire _guard3157 = fsm_out == 1'd0;
wire _guard3158 = cond_wire209_out;
wire _guard3159 = _guard3157 & _guard3158;
wire _guard3160 = fsm_out == 1'd0;
wire _guard3161 = _guard3159 & _guard3160;
wire _guard3162 = fsm_out == 1'd0;
wire _guard3163 = cond_wire211_out;
wire _guard3164 = _guard3162 & _guard3163;
wire _guard3165 = fsm_out == 1'd0;
wire _guard3166 = _guard3164 & _guard3165;
wire _guard3167 = _guard3161 | _guard3166;
wire _guard3168 = early_reset_static_par0_go_out;
wire _guard3169 = _guard3167 & _guard3168;
wire _guard3170 = cond_wire255_out;
wire _guard3171 = early_reset_static_par0_go_out;
wire _guard3172 = _guard3170 & _guard3171;
wire _guard3173 = cond_wire255_out;
wire _guard3174 = early_reset_static_par0_go_out;
wire _guard3175 = _guard3173 & _guard3174;
wire _guard3176 = early_reset_static_par_go_out;
wire _guard3177 = early_reset_static_par0_go_out;
wire _guard3178 = _guard3176 | _guard3177;
wire _guard3179 = early_reset_static_par0_go_out;
wire _guard3180 = early_reset_static_par_go_out;
wire _guard3181 = early_reset_static_par_go_out;
wire _guard3182 = early_reset_static_par0_go_out;
wire _guard3183 = _guard3181 | _guard3182;
wire _guard3184 = early_reset_static_par0_go_out;
wire _guard3185 = early_reset_static_par_go_out;
wire _guard3186 = early_reset_static_par_go_out;
wire _guard3187 = early_reset_static_par0_go_out;
wire _guard3188 = _guard3186 | _guard3187;
wire _guard3189 = early_reset_static_par_go_out;
wire _guard3190 = early_reset_static_par0_go_out;
wire _guard3191 = early_reset_static_par0_go_out;
wire _guard3192 = early_reset_static_par0_go_out;
wire _guard3193 = early_reset_static_par0_go_out;
wire _guard3194 = early_reset_static_par0_go_out;
wire _guard3195 = early_reset_static_par0_go_out;
wire _guard3196 = ~_guard0;
wire _guard3197 = early_reset_static_par0_go_out;
wire _guard3198 = _guard3196 & _guard3197;
wire _guard3199 = early_reset_static_par0_go_out;
wire _guard3200 = early_reset_static_par0_go_out;
wire _guard3201 = ~_guard0;
wire _guard3202 = early_reset_static_par0_go_out;
wire _guard3203 = _guard3201 & _guard3202;
wire _guard3204 = early_reset_static_par0_go_out;
wire _guard3205 = early_reset_static_par0_go_out;
wire _guard3206 = early_reset_static_par0_go_out;
wire _guard3207 = early_reset_static_par0_go_out;
wire _guard3208 = early_reset_static_par0_go_out;
wire _guard3209 = early_reset_static_par0_go_out;
wire _guard3210 = early_reset_static_par0_go_out;
wire _guard3211 = early_reset_static_par0_go_out;
wire _guard3212 = ~_guard0;
wire _guard3213 = early_reset_static_par0_go_out;
wire _guard3214 = _guard3212 & _guard3213;
wire _guard3215 = early_reset_static_par0_go_out;
wire _guard3216 = ~_guard0;
wire _guard3217 = early_reset_static_par0_go_out;
wire _guard3218 = _guard3216 & _guard3217;
wire _guard3219 = early_reset_static_par0_go_out;
wire _guard3220 = early_reset_static_par0_go_out;
wire _guard3221 = early_reset_static_par0_go_out;
wire _guard3222 = early_reset_static_par0_go_out;
wire _guard3223 = early_reset_static_par0_go_out;
wire _guard3224 = early_reset_static_par0_go_out;
wire _guard3225 = early_reset_static_par0_go_out;
wire _guard3226 = ~_guard0;
wire _guard3227 = early_reset_static_par0_go_out;
wire _guard3228 = _guard3226 & _guard3227;
wire _guard3229 = early_reset_static_par0_go_out;
wire _guard3230 = ~_guard0;
wire _guard3231 = early_reset_static_par0_go_out;
wire _guard3232 = _guard3230 & _guard3231;
wire _guard3233 = ~_guard0;
wire _guard3234 = early_reset_static_par0_go_out;
wire _guard3235 = _guard3233 & _guard3234;
wire _guard3236 = early_reset_static_par0_go_out;
wire _guard3237 = ~_guard0;
wire _guard3238 = early_reset_static_par0_go_out;
wire _guard3239 = _guard3237 & _guard3238;
wire _guard3240 = early_reset_static_par0_go_out;
wire _guard3241 = early_reset_static_par0_go_out;
wire _guard3242 = early_reset_static_par0_go_out;
wire _guard3243 = early_reset_static_par0_go_out;
wire _guard3244 = early_reset_static_par0_go_out;
wire _guard3245 = early_reset_static_par0_go_out;
wire _guard3246 = early_reset_static_par0_go_out;
wire _guard3247 = early_reset_static_par0_go_out;
wire _guard3248 = early_reset_static_par0_go_out;
wire _guard3249 = early_reset_static_par0_go_out;
wire _guard3250 = early_reset_static_par0_go_out;
wire _guard3251 = early_reset_static_par0_go_out;
wire _guard3252 = ~_guard0;
wire _guard3253 = early_reset_static_par0_go_out;
wire _guard3254 = _guard3252 & _guard3253;
wire _guard3255 = early_reset_static_par0_go_out;
wire _guard3256 = ~_guard0;
wire _guard3257 = early_reset_static_par0_go_out;
wire _guard3258 = _guard3256 & _guard3257;
wire _guard3259 = early_reset_static_par0_go_out;
wire _guard3260 = early_reset_static_par0_go_out;
wire _guard3261 = early_reset_static_par0_go_out;
wire _guard3262 = ~_guard0;
wire _guard3263 = early_reset_static_par0_go_out;
wire _guard3264 = _guard3262 & _guard3263;
wire _guard3265 = early_reset_static_par0_go_out;
wire _guard3266 = early_reset_static_par0_go_out;
wire _guard3267 = early_reset_static_par0_go_out;
wire _guard3268 = early_reset_static_par0_go_out;
wire _guard3269 = early_reset_static_par0_go_out;
wire _guard3270 = early_reset_static_par0_go_out;
wire _guard3271 = early_reset_static_par0_go_out;
wire _guard3272 = ~_guard0;
wire _guard3273 = early_reset_static_par0_go_out;
wire _guard3274 = _guard3272 & _guard3273;
wire _guard3275 = early_reset_static_par0_go_out;
wire _guard3276 = ~_guard0;
wire _guard3277 = early_reset_static_par0_go_out;
wire _guard3278 = _guard3276 & _guard3277;
wire _guard3279 = early_reset_static_par0_go_out;
wire _guard3280 = ~_guard0;
wire _guard3281 = early_reset_static_par0_go_out;
wire _guard3282 = _guard3280 & _guard3281;
wire _guard3283 = ~_guard0;
wire _guard3284 = early_reset_static_par0_go_out;
wire _guard3285 = _guard3283 & _guard3284;
wire _guard3286 = early_reset_static_par0_go_out;
wire _guard3287 = early_reset_static_par0_go_out;
wire _guard3288 = early_reset_static_par0_go_out;
wire _guard3289 = early_reset_static_par0_go_out;
wire _guard3290 = ~_guard0;
wire _guard3291 = early_reset_static_par0_go_out;
wire _guard3292 = _guard3290 & _guard3291;
wire _guard3293 = wrapper_early_reset_static_par_done_out;
wire _guard3294 = ~_guard3293;
wire _guard3295 = fsm0_out == 2'd0;
wire _guard3296 = _guard3294 & _guard3295;
wire _guard3297 = tdcc_go_out;
wire _guard3298 = _guard3296 & _guard3297;
wire _guard3299 = early_reset_static_par0_go_out;
wire _guard3300 = early_reset_static_par0_go_out;
wire _guard3301 = cond_wire12_out;
wire _guard3302 = early_reset_static_par0_go_out;
wire _guard3303 = _guard3301 & _guard3302;
wire _guard3304 = cond_wire10_out;
wire _guard3305 = early_reset_static_par0_go_out;
wire _guard3306 = _guard3304 & _guard3305;
wire _guard3307 = fsm_out == 1'd0;
wire _guard3308 = cond_wire10_out;
wire _guard3309 = _guard3307 & _guard3308;
wire _guard3310 = fsm_out == 1'd0;
wire _guard3311 = _guard3309 & _guard3310;
wire _guard3312 = fsm_out == 1'd0;
wire _guard3313 = cond_wire12_out;
wire _guard3314 = _guard3312 & _guard3313;
wire _guard3315 = fsm_out == 1'd0;
wire _guard3316 = _guard3314 & _guard3315;
wire _guard3317 = _guard3311 | _guard3316;
wire _guard3318 = early_reset_static_par0_go_out;
wire _guard3319 = _guard3317 & _guard3318;
wire _guard3320 = fsm_out == 1'd0;
wire _guard3321 = cond_wire10_out;
wire _guard3322 = _guard3320 & _guard3321;
wire _guard3323 = fsm_out == 1'd0;
wire _guard3324 = _guard3322 & _guard3323;
wire _guard3325 = fsm_out == 1'd0;
wire _guard3326 = cond_wire12_out;
wire _guard3327 = _guard3325 & _guard3326;
wire _guard3328 = fsm_out == 1'd0;
wire _guard3329 = _guard3327 & _guard3328;
wire _guard3330 = _guard3324 | _guard3329;
wire _guard3331 = early_reset_static_par0_go_out;
wire _guard3332 = _guard3330 & _guard3331;
wire _guard3333 = fsm_out == 1'd0;
wire _guard3334 = cond_wire10_out;
wire _guard3335 = _guard3333 & _guard3334;
wire _guard3336 = fsm_out == 1'd0;
wire _guard3337 = _guard3335 & _guard3336;
wire _guard3338 = fsm_out == 1'd0;
wire _guard3339 = cond_wire12_out;
wire _guard3340 = _guard3338 & _guard3339;
wire _guard3341 = fsm_out == 1'd0;
wire _guard3342 = _guard3340 & _guard3341;
wire _guard3343 = _guard3337 | _guard3342;
wire _guard3344 = early_reset_static_par0_go_out;
wire _guard3345 = _guard3343 & _guard3344;
wire _guard3346 = cond_wire66_out;
wire _guard3347 = early_reset_static_par0_go_out;
wire _guard3348 = _guard3346 & _guard3347;
wire _guard3349 = cond_wire64_out;
wire _guard3350 = early_reset_static_par0_go_out;
wire _guard3351 = _guard3349 & _guard3350;
wire _guard3352 = fsm_out == 1'd0;
wire _guard3353 = cond_wire64_out;
wire _guard3354 = _guard3352 & _guard3353;
wire _guard3355 = fsm_out == 1'd0;
wire _guard3356 = _guard3354 & _guard3355;
wire _guard3357 = fsm_out == 1'd0;
wire _guard3358 = cond_wire66_out;
wire _guard3359 = _guard3357 & _guard3358;
wire _guard3360 = fsm_out == 1'd0;
wire _guard3361 = _guard3359 & _guard3360;
wire _guard3362 = _guard3356 | _guard3361;
wire _guard3363 = early_reset_static_par0_go_out;
wire _guard3364 = _guard3362 & _guard3363;
wire _guard3365 = fsm_out == 1'd0;
wire _guard3366 = cond_wire64_out;
wire _guard3367 = _guard3365 & _guard3366;
wire _guard3368 = fsm_out == 1'd0;
wire _guard3369 = _guard3367 & _guard3368;
wire _guard3370 = fsm_out == 1'd0;
wire _guard3371 = cond_wire66_out;
wire _guard3372 = _guard3370 & _guard3371;
wire _guard3373 = fsm_out == 1'd0;
wire _guard3374 = _guard3372 & _guard3373;
wire _guard3375 = _guard3369 | _guard3374;
wire _guard3376 = early_reset_static_par0_go_out;
wire _guard3377 = _guard3375 & _guard3376;
wire _guard3378 = fsm_out == 1'd0;
wire _guard3379 = cond_wire64_out;
wire _guard3380 = _guard3378 & _guard3379;
wire _guard3381 = fsm_out == 1'd0;
wire _guard3382 = _guard3380 & _guard3381;
wire _guard3383 = fsm_out == 1'd0;
wire _guard3384 = cond_wire66_out;
wire _guard3385 = _guard3383 & _guard3384;
wire _guard3386 = fsm_out == 1'd0;
wire _guard3387 = _guard3385 & _guard3386;
wire _guard3388 = _guard3382 | _guard3387;
wire _guard3389 = early_reset_static_par0_go_out;
wire _guard3390 = _guard3388 & _guard3389;
wire _guard3391 = cond_wire123_out;
wire _guard3392 = early_reset_static_par0_go_out;
wire _guard3393 = _guard3391 & _guard3392;
wire _guard3394 = cond_wire123_out;
wire _guard3395 = early_reset_static_par0_go_out;
wire _guard3396 = _guard3394 & _guard3395;
wire _guard3397 = cond_wire160_out;
wire _guard3398 = early_reset_static_par0_go_out;
wire _guard3399 = _guard3397 & _guard3398;
wire _guard3400 = cond_wire160_out;
wire _guard3401 = early_reset_static_par0_go_out;
wire _guard3402 = _guard3400 & _guard3401;
wire _guard3403 = cond_wire206_out;
wire _guard3404 = early_reset_static_par0_go_out;
wire _guard3405 = _guard3403 & _guard3404;
wire _guard3406 = cond_wire206_out;
wire _guard3407 = early_reset_static_par0_go_out;
wire _guard3408 = _guard3406 & _guard3407;
wire _guard3409 = cond_wire227_out;
wire _guard3410 = early_reset_static_par0_go_out;
wire _guard3411 = _guard3409 & _guard3410;
wire _guard3412 = cond_wire225_out;
wire _guard3413 = early_reset_static_par0_go_out;
wire _guard3414 = _guard3412 & _guard3413;
wire _guard3415 = fsm_out == 1'd0;
wire _guard3416 = cond_wire225_out;
wire _guard3417 = _guard3415 & _guard3416;
wire _guard3418 = fsm_out == 1'd0;
wire _guard3419 = _guard3417 & _guard3418;
wire _guard3420 = fsm_out == 1'd0;
wire _guard3421 = cond_wire227_out;
wire _guard3422 = _guard3420 & _guard3421;
wire _guard3423 = fsm_out == 1'd0;
wire _guard3424 = _guard3422 & _guard3423;
wire _guard3425 = _guard3419 | _guard3424;
wire _guard3426 = early_reset_static_par0_go_out;
wire _guard3427 = _guard3425 & _guard3426;
wire _guard3428 = fsm_out == 1'd0;
wire _guard3429 = cond_wire225_out;
wire _guard3430 = _guard3428 & _guard3429;
wire _guard3431 = fsm_out == 1'd0;
wire _guard3432 = _guard3430 & _guard3431;
wire _guard3433 = fsm_out == 1'd0;
wire _guard3434 = cond_wire227_out;
wire _guard3435 = _guard3433 & _guard3434;
wire _guard3436 = fsm_out == 1'd0;
wire _guard3437 = _guard3435 & _guard3436;
wire _guard3438 = _guard3432 | _guard3437;
wire _guard3439 = early_reset_static_par0_go_out;
wire _guard3440 = _guard3438 & _guard3439;
wire _guard3441 = fsm_out == 1'd0;
wire _guard3442 = cond_wire225_out;
wire _guard3443 = _guard3441 & _guard3442;
wire _guard3444 = fsm_out == 1'd0;
wire _guard3445 = _guard3443 & _guard3444;
wire _guard3446 = fsm_out == 1'd0;
wire _guard3447 = cond_wire227_out;
wire _guard3448 = _guard3446 & _guard3447;
wire _guard3449 = fsm_out == 1'd0;
wire _guard3450 = _guard3448 & _guard3449;
wire _guard3451 = _guard3445 | _guard3450;
wire _guard3452 = early_reset_static_par0_go_out;
wire _guard3453 = _guard3451 & _guard3452;
wire _guard3454 = cond_wire230_out;
wire _guard3455 = early_reset_static_par0_go_out;
wire _guard3456 = _guard3454 & _guard3455;
wire _guard3457 = cond_wire230_out;
wire _guard3458 = early_reset_static_par0_go_out;
wire _guard3459 = _guard3457 & _guard3458;
wire _guard3460 = cond_wire240_out;
wire _guard3461 = early_reset_static_par0_go_out;
wire _guard3462 = _guard3460 & _guard3461;
wire _guard3463 = cond_wire238_out;
wire _guard3464 = early_reset_static_par0_go_out;
wire _guard3465 = _guard3463 & _guard3464;
wire _guard3466 = fsm_out == 1'd0;
wire _guard3467 = cond_wire238_out;
wire _guard3468 = _guard3466 & _guard3467;
wire _guard3469 = fsm_out == 1'd0;
wire _guard3470 = _guard3468 & _guard3469;
wire _guard3471 = fsm_out == 1'd0;
wire _guard3472 = cond_wire240_out;
wire _guard3473 = _guard3471 & _guard3472;
wire _guard3474 = fsm_out == 1'd0;
wire _guard3475 = _guard3473 & _guard3474;
wire _guard3476 = _guard3470 | _guard3475;
wire _guard3477 = early_reset_static_par0_go_out;
wire _guard3478 = _guard3476 & _guard3477;
wire _guard3479 = fsm_out == 1'd0;
wire _guard3480 = cond_wire238_out;
wire _guard3481 = _guard3479 & _guard3480;
wire _guard3482 = fsm_out == 1'd0;
wire _guard3483 = _guard3481 & _guard3482;
wire _guard3484 = fsm_out == 1'd0;
wire _guard3485 = cond_wire240_out;
wire _guard3486 = _guard3484 & _guard3485;
wire _guard3487 = fsm_out == 1'd0;
wire _guard3488 = _guard3486 & _guard3487;
wire _guard3489 = _guard3483 | _guard3488;
wire _guard3490 = early_reset_static_par0_go_out;
wire _guard3491 = _guard3489 & _guard3490;
wire _guard3492 = fsm_out == 1'd0;
wire _guard3493 = cond_wire238_out;
wire _guard3494 = _guard3492 & _guard3493;
wire _guard3495 = fsm_out == 1'd0;
wire _guard3496 = _guard3494 & _guard3495;
wire _guard3497 = fsm_out == 1'd0;
wire _guard3498 = cond_wire240_out;
wire _guard3499 = _guard3497 & _guard3498;
wire _guard3500 = fsm_out == 1'd0;
wire _guard3501 = _guard3499 & _guard3500;
wire _guard3502 = _guard3496 | _guard3501;
wire _guard3503 = early_reset_static_par0_go_out;
wire _guard3504 = _guard3502 & _guard3503;
wire _guard3505 = cond_wire222_out;
wire _guard3506 = early_reset_static_par0_go_out;
wire _guard3507 = _guard3505 & _guard3506;
wire _guard3508 = cond_wire222_out;
wire _guard3509 = early_reset_static_par0_go_out;
wire _guard3510 = _guard3508 & _guard3509;
wire _guard3511 = early_reset_static_par_go_out;
wire _guard3512 = cond_wire_out;
wire _guard3513 = early_reset_static_par0_go_out;
wire _guard3514 = _guard3512 & _guard3513;
wire _guard3515 = _guard3511 | _guard3514;
wire _guard3516 = early_reset_static_par_go_out;
wire _guard3517 = cond_wire_out;
wire _guard3518 = early_reset_static_par0_go_out;
wire _guard3519 = _guard3517 & _guard3518;
wire _guard3520 = early_reset_static_par_go_out;
wire _guard3521 = cond_wire19_out;
wire _guard3522 = early_reset_static_par0_go_out;
wire _guard3523 = _guard3521 & _guard3522;
wire _guard3524 = _guard3520 | _guard3523;
wire _guard3525 = early_reset_static_par_go_out;
wire _guard3526 = cond_wire19_out;
wire _guard3527 = early_reset_static_par0_go_out;
wire _guard3528 = _guard3526 & _guard3527;
wire _guard3529 = early_reset_static_par_go_out;
wire _guard3530 = cond_wire29_out;
wire _guard3531 = early_reset_static_par0_go_out;
wire _guard3532 = _guard3530 & _guard3531;
wire _guard3533 = _guard3529 | _guard3532;
wire _guard3534 = early_reset_static_par_go_out;
wire _guard3535 = cond_wire29_out;
wire _guard3536 = early_reset_static_par0_go_out;
wire _guard3537 = _guard3535 & _guard3536;
wire _guard3538 = early_reset_static_par_go_out;
wire _guard3539 = cond_wire39_out;
wire _guard3540 = early_reset_static_par0_go_out;
wire _guard3541 = _guard3539 & _guard3540;
wire _guard3542 = _guard3538 | _guard3541;
wire _guard3543 = cond_wire39_out;
wire _guard3544 = early_reset_static_par0_go_out;
wire _guard3545 = _guard3543 & _guard3544;
wire _guard3546 = early_reset_static_par_go_out;
wire _guard3547 = cond_wire171_out;
wire _guard3548 = early_reset_static_par0_go_out;
wire _guard3549 = _guard3547 & _guard3548;
wire _guard3550 = cond_wire171_out;
wire _guard3551 = early_reset_static_par0_go_out;
wire _guard3552 = _guard3550 & _guard3551;
wire _guard3553 = early_reset_static_par0_go_out;
wire _guard3554 = early_reset_static_par0_go_out;
wire _guard3555 = early_reset_static_par0_go_out;
wire _guard3556 = early_reset_static_par0_go_out;
wire _guard3557 = early_reset_static_par0_go_out;
wire _guard3558 = early_reset_static_par0_go_out;
wire _guard3559 = early_reset_static_par0_go_out;
wire _guard3560 = early_reset_static_par0_go_out;
wire _guard3561 = early_reset_static_par_go_out;
wire _guard3562 = early_reset_static_par0_go_out;
wire _guard3563 = _guard3561 | _guard3562;
wire _guard3564 = early_reset_static_par0_go_out;
wire _guard3565 = early_reset_static_par_go_out;
wire _guard3566 = early_reset_static_par0_go_out;
wire _guard3567 = early_reset_static_par0_go_out;
wire _guard3568 = early_reset_static_par0_go_out;
wire _guard3569 = early_reset_static_par0_go_out;
wire _guard3570 = early_reset_static_par_go_out;
wire _guard3571 = early_reset_static_par0_go_out;
wire _guard3572 = _guard3570 | _guard3571;
wire _guard3573 = early_reset_static_par0_go_out;
wire _guard3574 = early_reset_static_par_go_out;
wire _guard3575 = early_reset_static_par_go_out;
wire _guard3576 = early_reset_static_par0_go_out;
wire _guard3577 = _guard3575 | _guard3576;
wire _guard3578 = early_reset_static_par0_go_out;
wire _guard3579 = early_reset_static_par_go_out;
wire _guard3580 = early_reset_static_par_go_out;
wire _guard3581 = early_reset_static_par0_go_out;
wire _guard3582 = _guard3580 | _guard3581;
wire _guard3583 = early_reset_static_par0_go_out;
wire _guard3584 = early_reset_static_par_go_out;
wire _guard3585 = early_reset_static_par0_go_out;
wire _guard3586 = early_reset_static_par0_go_out;
wire _guard3587 = early_reset_static_par0_go_out;
wire _guard3588 = early_reset_static_par0_go_out;
wire _guard3589 = early_reset_static_par0_go_out;
wire _guard3590 = early_reset_static_par0_go_out;
wire _guard3591 = early_reset_static_par0_go_out;
wire _guard3592 = early_reset_static_par0_go_out;
wire _guard3593 = early_reset_static_par0_go_out;
wire _guard3594 = early_reset_static_par0_go_out;
wire _guard3595 = early_reset_static_par0_go_out;
wire _guard3596 = early_reset_static_par0_go_out;
wire _guard3597 = early_reset_static_par0_go_out;
wire _guard3598 = early_reset_static_par0_go_out;
wire _guard3599 = early_reset_static_par0_go_out;
wire _guard3600 = early_reset_static_par0_go_out;
wire _guard3601 = early_reset_static_par0_go_out;
wire _guard3602 = early_reset_static_par0_go_out;
wire _guard3603 = early_reset_static_par0_go_out;
wire _guard3604 = early_reset_static_par0_go_out;
wire _guard3605 = early_reset_static_par0_go_out;
wire _guard3606 = early_reset_static_par0_go_out;
wire _guard3607 = early_reset_static_par0_go_out;
wire _guard3608 = early_reset_static_par0_go_out;
wire _guard3609 = ~_guard0;
wire _guard3610 = early_reset_static_par0_go_out;
wire _guard3611 = _guard3609 & _guard3610;
wire _guard3612 = early_reset_static_par0_go_out;
wire _guard3613 = early_reset_static_par0_go_out;
wire _guard3614 = early_reset_static_par0_go_out;
wire _guard3615 = early_reset_static_par0_go_out;
wire _guard3616 = early_reset_static_par0_go_out;
wire _guard3617 = early_reset_static_par0_go_out;
wire _guard3618 = early_reset_static_par0_go_out;
wire _guard3619 = ~_guard0;
wire _guard3620 = early_reset_static_par0_go_out;
wire _guard3621 = _guard3619 & _guard3620;
wire _guard3622 = early_reset_static_par0_go_out;
wire _guard3623 = early_reset_static_par0_go_out;
wire _guard3624 = early_reset_static_par0_go_out;
wire _guard3625 = early_reset_static_par0_go_out;
wire _guard3626 = early_reset_static_par0_go_out;
wire _guard3627 = early_reset_static_par0_go_out;
wire _guard3628 = early_reset_static_par0_go_out;
wire _guard3629 = early_reset_static_par0_go_out;
wire _guard3630 = early_reset_static_par0_go_out;
wire _guard3631 = early_reset_static_par0_go_out;
wire _guard3632 = ~_guard0;
wire _guard3633 = early_reset_static_par0_go_out;
wire _guard3634 = _guard3632 & _guard3633;
wire _guard3635 = early_reset_static_par0_go_out;
wire _guard3636 = ~_guard0;
wire _guard3637 = early_reset_static_par0_go_out;
wire _guard3638 = _guard3636 & _guard3637;
wire _guard3639 = early_reset_static_par0_go_out;
wire _guard3640 = ~_guard0;
wire _guard3641 = early_reset_static_par0_go_out;
wire _guard3642 = _guard3640 & _guard3641;
wire _guard3643 = ~_guard0;
wire _guard3644 = early_reset_static_par0_go_out;
wire _guard3645 = _guard3643 & _guard3644;
wire _guard3646 = early_reset_static_par0_go_out;
wire _guard3647 = ~_guard0;
wire _guard3648 = early_reset_static_par0_go_out;
wire _guard3649 = _guard3647 & _guard3648;
wire _guard3650 = early_reset_static_par0_go_out;
wire _guard3651 = early_reset_static_par0_go_out;
wire _guard3652 = ~_guard0;
wire _guard3653 = early_reset_static_par0_go_out;
wire _guard3654 = _guard3652 & _guard3653;
wire _guard3655 = ~_guard0;
wire _guard3656 = early_reset_static_par0_go_out;
wire _guard3657 = _guard3655 & _guard3656;
wire _guard3658 = early_reset_static_par0_go_out;
wire _guard3659 = early_reset_static_par0_go_out;
wire _guard3660 = early_reset_static_par0_go_out;
wire _guard3661 = ~_guard0;
wire _guard3662 = early_reset_static_par0_go_out;
wire _guard3663 = _guard3661 & _guard3662;
wire _guard3664 = early_reset_static_par0_go_out;
wire _guard3665 = early_reset_static_par0_go_out;
wire _guard3666 = early_reset_static_par0_go_out;
wire _guard3667 = early_reset_static_par0_go_out;
wire _guard3668 = early_reset_static_par0_go_out;
wire _guard3669 = early_reset_static_par0_go_out;
wire _guard3670 = early_reset_static_par0_go_out;
wire _guard3671 = early_reset_static_par0_go_out;
wire _guard3672 = early_reset_static_par0_go_out;
wire _guard3673 = early_reset_static_par0_go_out;
wire _guard3674 = early_reset_static_par0_go_out;
wire _guard3675 = early_reset_static_par0_go_out;
wire _guard3676 = early_reset_static_par0_go_out;
wire _guard3677 = early_reset_static_par0_go_out;
wire _guard3678 = early_reset_static_par0_go_out;
wire _guard3679 = early_reset_static_par0_go_out;
wire _guard3680 = ~_guard0;
wire _guard3681 = early_reset_static_par0_go_out;
wire _guard3682 = _guard3680 & _guard3681;
wire _guard3683 = early_reset_static_par0_go_out;
wire _guard3684 = ~_guard0;
wire _guard3685 = early_reset_static_par0_go_out;
wire _guard3686 = _guard3684 & _guard3685;
wire _guard3687 = ~_guard0;
wire _guard3688 = early_reset_static_par0_go_out;
wire _guard3689 = _guard3687 & _guard3688;
wire _guard3690 = early_reset_static_par0_go_out;
wire _guard3691 = early_reset_static_par0_go_out;
wire _guard3692 = early_reset_static_par0_go_out;
wire _guard3693 = early_reset_static_par0_go_out;
wire _guard3694 = ~_guard0;
wire _guard3695 = early_reset_static_par0_go_out;
wire _guard3696 = _guard3694 & _guard3695;
wire _guard3697 = fsm_out == 1'd0;
wire _guard3698 = signal_reg_out;
wire _guard3699 = _guard3697 & _guard3698;
wire _guard3700 = cond_wire31_out;
wire _guard3701 = early_reset_static_par0_go_out;
wire _guard3702 = _guard3700 & _guard3701;
wire _guard3703 = cond_wire31_out;
wire _guard3704 = early_reset_static_par0_go_out;
wire _guard3705 = _guard3703 & _guard3704;
wire _guard3706 = cond_wire79_out;
wire _guard3707 = early_reset_static_par0_go_out;
wire _guard3708 = _guard3706 & _guard3707;
wire _guard3709 = cond_wire77_out;
wire _guard3710 = early_reset_static_par0_go_out;
wire _guard3711 = _guard3709 & _guard3710;
wire _guard3712 = fsm_out == 1'd0;
wire _guard3713 = cond_wire77_out;
wire _guard3714 = _guard3712 & _guard3713;
wire _guard3715 = fsm_out == 1'd0;
wire _guard3716 = _guard3714 & _guard3715;
wire _guard3717 = fsm_out == 1'd0;
wire _guard3718 = cond_wire79_out;
wire _guard3719 = _guard3717 & _guard3718;
wire _guard3720 = fsm_out == 1'd0;
wire _guard3721 = _guard3719 & _guard3720;
wire _guard3722 = _guard3716 | _guard3721;
wire _guard3723 = early_reset_static_par0_go_out;
wire _guard3724 = _guard3722 & _guard3723;
wire _guard3725 = fsm_out == 1'd0;
wire _guard3726 = cond_wire77_out;
wire _guard3727 = _guard3725 & _guard3726;
wire _guard3728 = fsm_out == 1'd0;
wire _guard3729 = _guard3727 & _guard3728;
wire _guard3730 = fsm_out == 1'd0;
wire _guard3731 = cond_wire79_out;
wire _guard3732 = _guard3730 & _guard3731;
wire _guard3733 = fsm_out == 1'd0;
wire _guard3734 = _guard3732 & _guard3733;
wire _guard3735 = _guard3729 | _guard3734;
wire _guard3736 = early_reset_static_par0_go_out;
wire _guard3737 = _guard3735 & _guard3736;
wire _guard3738 = fsm_out == 1'd0;
wire _guard3739 = cond_wire77_out;
wire _guard3740 = _guard3738 & _guard3739;
wire _guard3741 = fsm_out == 1'd0;
wire _guard3742 = _guard3740 & _guard3741;
wire _guard3743 = fsm_out == 1'd0;
wire _guard3744 = cond_wire79_out;
wire _guard3745 = _guard3743 & _guard3744;
wire _guard3746 = fsm_out == 1'd0;
wire _guard3747 = _guard3745 & _guard3746;
wire _guard3748 = _guard3742 | _guard3747;
wire _guard3749 = early_reset_static_par0_go_out;
wire _guard3750 = _guard3748 & _guard3749;
wire _guard3751 = cond_wire87_out;
wire _guard3752 = early_reset_static_par0_go_out;
wire _guard3753 = _guard3751 & _guard3752;
wire _guard3754 = cond_wire85_out;
wire _guard3755 = early_reset_static_par0_go_out;
wire _guard3756 = _guard3754 & _guard3755;
wire _guard3757 = fsm_out == 1'd0;
wire _guard3758 = cond_wire85_out;
wire _guard3759 = _guard3757 & _guard3758;
wire _guard3760 = fsm_out == 1'd0;
wire _guard3761 = _guard3759 & _guard3760;
wire _guard3762 = fsm_out == 1'd0;
wire _guard3763 = cond_wire87_out;
wire _guard3764 = _guard3762 & _guard3763;
wire _guard3765 = fsm_out == 1'd0;
wire _guard3766 = _guard3764 & _guard3765;
wire _guard3767 = _guard3761 | _guard3766;
wire _guard3768 = early_reset_static_par0_go_out;
wire _guard3769 = _guard3767 & _guard3768;
wire _guard3770 = fsm_out == 1'd0;
wire _guard3771 = cond_wire85_out;
wire _guard3772 = _guard3770 & _guard3771;
wire _guard3773 = fsm_out == 1'd0;
wire _guard3774 = _guard3772 & _guard3773;
wire _guard3775 = fsm_out == 1'd0;
wire _guard3776 = cond_wire87_out;
wire _guard3777 = _guard3775 & _guard3776;
wire _guard3778 = fsm_out == 1'd0;
wire _guard3779 = _guard3777 & _guard3778;
wire _guard3780 = _guard3774 | _guard3779;
wire _guard3781 = early_reset_static_par0_go_out;
wire _guard3782 = _guard3780 & _guard3781;
wire _guard3783 = fsm_out == 1'd0;
wire _guard3784 = cond_wire85_out;
wire _guard3785 = _guard3783 & _guard3784;
wire _guard3786 = fsm_out == 1'd0;
wire _guard3787 = _guard3785 & _guard3786;
wire _guard3788 = fsm_out == 1'd0;
wire _guard3789 = cond_wire87_out;
wire _guard3790 = _guard3788 & _guard3789;
wire _guard3791 = fsm_out == 1'd0;
wire _guard3792 = _guard3790 & _guard3791;
wire _guard3793 = _guard3787 | _guard3792;
wire _guard3794 = early_reset_static_par0_go_out;
wire _guard3795 = _guard3793 & _guard3794;
wire _guard3796 = cond_wire95_out;
wire _guard3797 = early_reset_static_par0_go_out;
wire _guard3798 = _guard3796 & _guard3797;
wire _guard3799 = cond_wire93_out;
wire _guard3800 = early_reset_static_par0_go_out;
wire _guard3801 = _guard3799 & _guard3800;
wire _guard3802 = fsm_out == 1'd0;
wire _guard3803 = cond_wire93_out;
wire _guard3804 = _guard3802 & _guard3803;
wire _guard3805 = fsm_out == 1'd0;
wire _guard3806 = _guard3804 & _guard3805;
wire _guard3807 = fsm_out == 1'd0;
wire _guard3808 = cond_wire95_out;
wire _guard3809 = _guard3807 & _guard3808;
wire _guard3810 = fsm_out == 1'd0;
wire _guard3811 = _guard3809 & _guard3810;
wire _guard3812 = _guard3806 | _guard3811;
wire _guard3813 = early_reset_static_par0_go_out;
wire _guard3814 = _guard3812 & _guard3813;
wire _guard3815 = fsm_out == 1'd0;
wire _guard3816 = cond_wire93_out;
wire _guard3817 = _guard3815 & _guard3816;
wire _guard3818 = fsm_out == 1'd0;
wire _guard3819 = _guard3817 & _guard3818;
wire _guard3820 = fsm_out == 1'd0;
wire _guard3821 = cond_wire95_out;
wire _guard3822 = _guard3820 & _guard3821;
wire _guard3823 = fsm_out == 1'd0;
wire _guard3824 = _guard3822 & _guard3823;
wire _guard3825 = _guard3819 | _guard3824;
wire _guard3826 = early_reset_static_par0_go_out;
wire _guard3827 = _guard3825 & _guard3826;
wire _guard3828 = fsm_out == 1'd0;
wire _guard3829 = cond_wire93_out;
wire _guard3830 = _guard3828 & _guard3829;
wire _guard3831 = fsm_out == 1'd0;
wire _guard3832 = _guard3830 & _guard3831;
wire _guard3833 = fsm_out == 1'd0;
wire _guard3834 = cond_wire95_out;
wire _guard3835 = _guard3833 & _guard3834;
wire _guard3836 = fsm_out == 1'd0;
wire _guard3837 = _guard3835 & _guard3836;
wire _guard3838 = _guard3832 | _guard3837;
wire _guard3839 = early_reset_static_par0_go_out;
wire _guard3840 = _guard3838 & _guard3839;
wire _guard3841 = cond_wire112_out;
wire _guard3842 = early_reset_static_par0_go_out;
wire _guard3843 = _guard3841 & _guard3842;
wire _guard3844 = cond_wire110_out;
wire _guard3845 = early_reset_static_par0_go_out;
wire _guard3846 = _guard3844 & _guard3845;
wire _guard3847 = fsm_out == 1'd0;
wire _guard3848 = cond_wire110_out;
wire _guard3849 = _guard3847 & _guard3848;
wire _guard3850 = fsm_out == 1'd0;
wire _guard3851 = _guard3849 & _guard3850;
wire _guard3852 = fsm_out == 1'd0;
wire _guard3853 = cond_wire112_out;
wire _guard3854 = _guard3852 & _guard3853;
wire _guard3855 = fsm_out == 1'd0;
wire _guard3856 = _guard3854 & _guard3855;
wire _guard3857 = _guard3851 | _guard3856;
wire _guard3858 = early_reset_static_par0_go_out;
wire _guard3859 = _guard3857 & _guard3858;
wire _guard3860 = fsm_out == 1'd0;
wire _guard3861 = cond_wire110_out;
wire _guard3862 = _guard3860 & _guard3861;
wire _guard3863 = fsm_out == 1'd0;
wire _guard3864 = _guard3862 & _guard3863;
wire _guard3865 = fsm_out == 1'd0;
wire _guard3866 = cond_wire112_out;
wire _guard3867 = _guard3865 & _guard3866;
wire _guard3868 = fsm_out == 1'd0;
wire _guard3869 = _guard3867 & _guard3868;
wire _guard3870 = _guard3864 | _guard3869;
wire _guard3871 = early_reset_static_par0_go_out;
wire _guard3872 = _guard3870 & _guard3871;
wire _guard3873 = fsm_out == 1'd0;
wire _guard3874 = cond_wire110_out;
wire _guard3875 = _guard3873 & _guard3874;
wire _guard3876 = fsm_out == 1'd0;
wire _guard3877 = _guard3875 & _guard3876;
wire _guard3878 = fsm_out == 1'd0;
wire _guard3879 = cond_wire112_out;
wire _guard3880 = _guard3878 & _guard3879;
wire _guard3881 = fsm_out == 1'd0;
wire _guard3882 = _guard3880 & _guard3881;
wire _guard3883 = _guard3877 | _guard3882;
wire _guard3884 = early_reset_static_par0_go_out;
wire _guard3885 = _guard3883 & _guard3884;
wire _guard3886 = cond_wire90_out;
wire _guard3887 = early_reset_static_par0_go_out;
wire _guard3888 = _guard3886 & _guard3887;
wire _guard3889 = cond_wire90_out;
wire _guard3890 = early_reset_static_par0_go_out;
wire _guard3891 = _guard3889 & _guard3890;
wire _guard3892 = cond_wire186_out;
wire _guard3893 = early_reset_static_par0_go_out;
wire _guard3894 = _guard3892 & _guard3893;
wire _guard3895 = cond_wire184_out;
wire _guard3896 = early_reset_static_par0_go_out;
wire _guard3897 = _guard3895 & _guard3896;
wire _guard3898 = fsm_out == 1'd0;
wire _guard3899 = cond_wire184_out;
wire _guard3900 = _guard3898 & _guard3899;
wire _guard3901 = fsm_out == 1'd0;
wire _guard3902 = _guard3900 & _guard3901;
wire _guard3903 = fsm_out == 1'd0;
wire _guard3904 = cond_wire186_out;
wire _guard3905 = _guard3903 & _guard3904;
wire _guard3906 = fsm_out == 1'd0;
wire _guard3907 = _guard3905 & _guard3906;
wire _guard3908 = _guard3902 | _guard3907;
wire _guard3909 = early_reset_static_par0_go_out;
wire _guard3910 = _guard3908 & _guard3909;
wire _guard3911 = fsm_out == 1'd0;
wire _guard3912 = cond_wire184_out;
wire _guard3913 = _guard3911 & _guard3912;
wire _guard3914 = fsm_out == 1'd0;
wire _guard3915 = _guard3913 & _guard3914;
wire _guard3916 = fsm_out == 1'd0;
wire _guard3917 = cond_wire186_out;
wire _guard3918 = _guard3916 & _guard3917;
wire _guard3919 = fsm_out == 1'd0;
wire _guard3920 = _guard3918 & _guard3919;
wire _guard3921 = _guard3915 | _guard3920;
wire _guard3922 = early_reset_static_par0_go_out;
wire _guard3923 = _guard3921 & _guard3922;
wire _guard3924 = fsm_out == 1'd0;
wire _guard3925 = cond_wire184_out;
wire _guard3926 = _guard3924 & _guard3925;
wire _guard3927 = fsm_out == 1'd0;
wire _guard3928 = _guard3926 & _guard3927;
wire _guard3929 = fsm_out == 1'd0;
wire _guard3930 = cond_wire186_out;
wire _guard3931 = _guard3929 & _guard3930;
wire _guard3932 = fsm_out == 1'd0;
wire _guard3933 = _guard3931 & _guard3932;
wire _guard3934 = _guard3928 | _guard3933;
wire _guard3935 = early_reset_static_par0_go_out;
wire _guard3936 = _guard3934 & _guard3935;
wire _guard3937 = cond_wire194_out;
wire _guard3938 = early_reset_static_par0_go_out;
wire _guard3939 = _guard3937 & _guard3938;
wire _guard3940 = cond_wire192_out;
wire _guard3941 = early_reset_static_par0_go_out;
wire _guard3942 = _guard3940 & _guard3941;
wire _guard3943 = fsm_out == 1'd0;
wire _guard3944 = cond_wire192_out;
wire _guard3945 = _guard3943 & _guard3944;
wire _guard3946 = fsm_out == 1'd0;
wire _guard3947 = _guard3945 & _guard3946;
wire _guard3948 = fsm_out == 1'd0;
wire _guard3949 = cond_wire194_out;
wire _guard3950 = _guard3948 & _guard3949;
wire _guard3951 = fsm_out == 1'd0;
wire _guard3952 = _guard3950 & _guard3951;
wire _guard3953 = _guard3947 | _guard3952;
wire _guard3954 = early_reset_static_par0_go_out;
wire _guard3955 = _guard3953 & _guard3954;
wire _guard3956 = fsm_out == 1'd0;
wire _guard3957 = cond_wire192_out;
wire _guard3958 = _guard3956 & _guard3957;
wire _guard3959 = fsm_out == 1'd0;
wire _guard3960 = _guard3958 & _guard3959;
wire _guard3961 = fsm_out == 1'd0;
wire _guard3962 = cond_wire194_out;
wire _guard3963 = _guard3961 & _guard3962;
wire _guard3964 = fsm_out == 1'd0;
wire _guard3965 = _guard3963 & _guard3964;
wire _guard3966 = _guard3960 | _guard3965;
wire _guard3967 = early_reset_static_par0_go_out;
wire _guard3968 = _guard3966 & _guard3967;
wire _guard3969 = fsm_out == 1'd0;
wire _guard3970 = cond_wire192_out;
wire _guard3971 = _guard3969 & _guard3970;
wire _guard3972 = fsm_out == 1'd0;
wire _guard3973 = _guard3971 & _guard3972;
wire _guard3974 = fsm_out == 1'd0;
wire _guard3975 = cond_wire194_out;
wire _guard3976 = _guard3974 & _guard3975;
wire _guard3977 = fsm_out == 1'd0;
wire _guard3978 = _guard3976 & _guard3977;
wire _guard3979 = _guard3973 | _guard3978;
wire _guard3980 = early_reset_static_par0_go_out;
wire _guard3981 = _guard3979 & _guard3980;
wire _guard3982 = cond_wire215_out;
wire _guard3983 = early_reset_static_par0_go_out;
wire _guard3984 = _guard3982 & _guard3983;
wire _guard3985 = cond_wire213_out;
wire _guard3986 = early_reset_static_par0_go_out;
wire _guard3987 = _guard3985 & _guard3986;
wire _guard3988 = fsm_out == 1'd0;
wire _guard3989 = cond_wire213_out;
wire _guard3990 = _guard3988 & _guard3989;
wire _guard3991 = fsm_out == 1'd0;
wire _guard3992 = _guard3990 & _guard3991;
wire _guard3993 = fsm_out == 1'd0;
wire _guard3994 = cond_wire215_out;
wire _guard3995 = _guard3993 & _guard3994;
wire _guard3996 = fsm_out == 1'd0;
wire _guard3997 = _guard3995 & _guard3996;
wire _guard3998 = _guard3992 | _guard3997;
wire _guard3999 = early_reset_static_par0_go_out;
wire _guard4000 = _guard3998 & _guard3999;
wire _guard4001 = fsm_out == 1'd0;
wire _guard4002 = cond_wire213_out;
wire _guard4003 = _guard4001 & _guard4002;
wire _guard4004 = fsm_out == 1'd0;
wire _guard4005 = _guard4003 & _guard4004;
wire _guard4006 = fsm_out == 1'd0;
wire _guard4007 = cond_wire215_out;
wire _guard4008 = _guard4006 & _guard4007;
wire _guard4009 = fsm_out == 1'd0;
wire _guard4010 = _guard4008 & _guard4009;
wire _guard4011 = _guard4005 | _guard4010;
wire _guard4012 = early_reset_static_par0_go_out;
wire _guard4013 = _guard4011 & _guard4012;
wire _guard4014 = fsm_out == 1'd0;
wire _guard4015 = cond_wire213_out;
wire _guard4016 = _guard4014 & _guard4015;
wire _guard4017 = fsm_out == 1'd0;
wire _guard4018 = _guard4016 & _guard4017;
wire _guard4019 = fsm_out == 1'd0;
wire _guard4020 = cond_wire215_out;
wire _guard4021 = _guard4019 & _guard4020;
wire _guard4022 = fsm_out == 1'd0;
wire _guard4023 = _guard4021 & _guard4022;
wire _guard4024 = _guard4018 | _guard4023;
wire _guard4025 = early_reset_static_par0_go_out;
wire _guard4026 = _guard4024 & _guard4025;
wire _guard4027 = cond_wire219_out;
wire _guard4028 = early_reset_static_par0_go_out;
wire _guard4029 = _guard4027 & _guard4028;
wire _guard4030 = cond_wire217_out;
wire _guard4031 = early_reset_static_par0_go_out;
wire _guard4032 = _guard4030 & _guard4031;
wire _guard4033 = fsm_out == 1'd0;
wire _guard4034 = cond_wire217_out;
wire _guard4035 = _guard4033 & _guard4034;
wire _guard4036 = fsm_out == 1'd0;
wire _guard4037 = _guard4035 & _guard4036;
wire _guard4038 = fsm_out == 1'd0;
wire _guard4039 = cond_wire219_out;
wire _guard4040 = _guard4038 & _guard4039;
wire _guard4041 = fsm_out == 1'd0;
wire _guard4042 = _guard4040 & _guard4041;
wire _guard4043 = _guard4037 | _guard4042;
wire _guard4044 = early_reset_static_par0_go_out;
wire _guard4045 = _guard4043 & _guard4044;
wire _guard4046 = fsm_out == 1'd0;
wire _guard4047 = cond_wire217_out;
wire _guard4048 = _guard4046 & _guard4047;
wire _guard4049 = fsm_out == 1'd0;
wire _guard4050 = _guard4048 & _guard4049;
wire _guard4051 = fsm_out == 1'd0;
wire _guard4052 = cond_wire219_out;
wire _guard4053 = _guard4051 & _guard4052;
wire _guard4054 = fsm_out == 1'd0;
wire _guard4055 = _guard4053 & _guard4054;
wire _guard4056 = _guard4050 | _guard4055;
wire _guard4057 = early_reset_static_par0_go_out;
wire _guard4058 = _guard4056 & _guard4057;
wire _guard4059 = fsm_out == 1'd0;
wire _guard4060 = cond_wire217_out;
wire _guard4061 = _guard4059 & _guard4060;
wire _guard4062 = fsm_out == 1'd0;
wire _guard4063 = _guard4061 & _guard4062;
wire _guard4064 = fsm_out == 1'd0;
wire _guard4065 = cond_wire219_out;
wire _guard4066 = _guard4064 & _guard4065;
wire _guard4067 = fsm_out == 1'd0;
wire _guard4068 = _guard4066 & _guard4067;
wire _guard4069 = _guard4063 | _guard4068;
wire _guard4070 = early_reset_static_par0_go_out;
wire _guard4071 = _guard4069 & _guard4070;
wire _guard4072 = cond_wire239_out;
wire _guard4073 = early_reset_static_par0_go_out;
wire _guard4074 = _guard4072 & _guard4073;
wire _guard4075 = cond_wire239_out;
wire _guard4076 = early_reset_static_par0_go_out;
wire _guard4077 = _guard4075 & _guard4076;
wire _guard4078 = cond_wire247_out;
wire _guard4079 = early_reset_static_par0_go_out;
wire _guard4080 = _guard4078 & _guard4079;
wire _guard4081 = cond_wire247_out;
wire _guard4082 = early_reset_static_par0_go_out;
wire _guard4083 = _guard4081 & _guard4082;
wire _guard4084 = cond_wire226_out;
wire _guard4085 = early_reset_static_par0_go_out;
wire _guard4086 = _guard4084 & _guard4085;
wire _guard4087 = cond_wire226_out;
wire _guard4088 = early_reset_static_par0_go_out;
wire _guard4089 = _guard4087 & _guard4088;
wire _guard4090 = cond_wire19_out;
wire _guard4091 = early_reset_static_par0_go_out;
wire _guard4092 = _guard4090 & _guard4091;
wire _guard4093 = cond_wire19_out;
wire _guard4094 = early_reset_static_par0_go_out;
wire _guard4095 = _guard4093 & _guard4094;
wire _guard4096 = early_reset_static_par_go_out;
wire _guard4097 = cond_wire24_out;
wire _guard4098 = early_reset_static_par0_go_out;
wire _guard4099 = _guard4097 & _guard4098;
wire _guard4100 = _guard4096 | _guard4099;
wire _guard4101 = early_reset_static_par_go_out;
wire _guard4102 = cond_wire24_out;
wire _guard4103 = early_reset_static_par0_go_out;
wire _guard4104 = _guard4102 & _guard4103;
wire _guard4105 = cond_wire29_out;
wire _guard4106 = early_reset_static_par0_go_out;
wire _guard4107 = _guard4105 & _guard4106;
wire _guard4108 = cond_wire29_out;
wire _guard4109 = early_reset_static_par0_go_out;
wire _guard4110 = _guard4108 & _guard4109;
wire _guard4111 = early_reset_static_par_go_out;
wire _guard4112 = early_reset_static_par0_go_out;
wire _guard4113 = early_reset_static_par_go_out;
wire _guard4114 = early_reset_static_par0_go_out;
wire _guard4115 = early_reset_static_par0_go_out;
wire _guard4116 = early_reset_static_par0_go_out;
wire _guard4117 = early_reset_static_par0_go_out;
wire _guard4118 = early_reset_static_par0_go_out;
wire _guard4119 = early_reset_static_par_go_out;
wire _guard4120 = early_reset_static_par0_go_out;
wire _guard4121 = _guard4119 | _guard4120;
wire _guard4122 = early_reset_static_par_go_out;
wire _guard4123 = early_reset_static_par0_go_out;
wire _guard4124 = early_reset_static_par0_go_out;
wire _guard4125 = early_reset_static_par0_go_out;
wire _guard4126 = early_reset_static_par_go_out;
wire _guard4127 = early_reset_static_par0_go_out;
wire _guard4128 = _guard4126 | _guard4127;
wire _guard4129 = early_reset_static_par0_go_out;
wire _guard4130 = early_reset_static_par_go_out;
wire _guard4131 = early_reset_static_par0_go_out;
wire _guard4132 = early_reset_static_par0_go_out;
wire _guard4133 = early_reset_static_par_go_out;
wire _guard4134 = early_reset_static_par0_go_out;
wire _guard4135 = _guard4133 | _guard4134;
wire _guard4136 = early_reset_static_par0_go_out;
wire _guard4137 = early_reset_static_par_go_out;
wire _guard4138 = early_reset_static_par0_go_out;
wire _guard4139 = early_reset_static_par0_go_out;
wire _guard4140 = early_reset_static_par0_go_out;
wire _guard4141 = early_reset_static_par0_go_out;
wire _guard4142 = early_reset_static_par0_go_out;
wire _guard4143 = early_reset_static_par0_go_out;
wire _guard4144 = early_reset_static_par0_go_out;
wire _guard4145 = early_reset_static_par0_go_out;
wire _guard4146 = early_reset_static_par0_go_out;
wire _guard4147 = ~_guard0;
wire _guard4148 = early_reset_static_par0_go_out;
wire _guard4149 = _guard4147 & _guard4148;
wire _guard4150 = early_reset_static_par0_go_out;
wire _guard4151 = early_reset_static_par0_go_out;
wire _guard4152 = early_reset_static_par0_go_out;
wire _guard4153 = early_reset_static_par0_go_out;
wire _guard4154 = ~_guard0;
wire _guard4155 = early_reset_static_par0_go_out;
wire _guard4156 = _guard4154 & _guard4155;
wire _guard4157 = early_reset_static_par0_go_out;
wire _guard4158 = early_reset_static_par0_go_out;
wire _guard4159 = early_reset_static_par0_go_out;
wire _guard4160 = early_reset_static_par0_go_out;
wire _guard4161 = early_reset_static_par0_go_out;
wire _guard4162 = early_reset_static_par0_go_out;
wire _guard4163 = early_reset_static_par0_go_out;
wire _guard4164 = early_reset_static_par0_go_out;
wire _guard4165 = early_reset_static_par0_go_out;
wire _guard4166 = early_reset_static_par0_go_out;
wire _guard4167 = early_reset_static_par0_go_out;
wire _guard4168 = early_reset_static_par0_go_out;
wire _guard4169 = early_reset_static_par0_go_out;
wire _guard4170 = ~_guard0;
wire _guard4171 = early_reset_static_par0_go_out;
wire _guard4172 = _guard4170 & _guard4171;
wire _guard4173 = early_reset_static_par0_go_out;
wire _guard4174 = ~_guard0;
wire _guard4175 = early_reset_static_par0_go_out;
wire _guard4176 = _guard4174 & _guard4175;
wire _guard4177 = early_reset_static_par0_go_out;
wire _guard4178 = early_reset_static_par0_go_out;
wire _guard4179 = ~_guard0;
wire _guard4180 = early_reset_static_par0_go_out;
wire _guard4181 = _guard4179 & _guard4180;
wire _guard4182 = early_reset_static_par0_go_out;
wire _guard4183 = early_reset_static_par0_go_out;
wire _guard4184 = early_reset_static_par0_go_out;
wire _guard4185 = early_reset_static_par0_go_out;
wire _guard4186 = early_reset_static_par0_go_out;
wire _guard4187 = early_reset_static_par0_go_out;
wire _guard4188 = early_reset_static_par0_go_out;
wire _guard4189 = ~_guard0;
wire _guard4190 = early_reset_static_par0_go_out;
wire _guard4191 = _guard4189 & _guard4190;
wire _guard4192 = early_reset_static_par0_go_out;
wire _guard4193 = early_reset_static_par0_go_out;
wire _guard4194 = early_reset_static_par0_go_out;
wire _guard4195 = early_reset_static_par0_go_out;
wire _guard4196 = early_reset_static_par0_go_out;
wire _guard4197 = ~_guard0;
wire _guard4198 = early_reset_static_par0_go_out;
wire _guard4199 = _guard4197 & _guard4198;
wire _guard4200 = early_reset_static_par0_go_out;
wire _guard4201 = early_reset_static_par0_go_out;
wire _guard4202 = early_reset_static_par0_go_out;
wire _guard4203 = ~_guard0;
wire _guard4204 = early_reset_static_par0_go_out;
wire _guard4205 = _guard4203 & _guard4204;
wire _guard4206 = early_reset_static_par0_go_out;
wire _guard4207 = early_reset_static_par0_go_out;
wire _guard4208 = early_reset_static_par0_go_out;
wire _guard4209 = early_reset_static_par0_go_out;
wire _guard4210 = ~_guard0;
wire _guard4211 = early_reset_static_par0_go_out;
wire _guard4212 = _guard4210 & _guard4211;
wire _guard4213 = early_reset_static_par0_go_out;
wire _guard4214 = early_reset_static_par0_go_out;
wire _guard4215 = early_reset_static_par0_go_out;
wire _guard4216 = early_reset_static_par0_go_out;
wire _guard4217 = early_reset_static_par0_go_out;
wire _guard4218 = fsm0_out == 2'd2;
wire _guard4219 = fsm0_out == 2'd0;
wire _guard4220 = wrapper_early_reset_static_par_done_out;
wire _guard4221 = _guard4219 & _guard4220;
wire _guard4222 = tdcc_go_out;
wire _guard4223 = _guard4221 & _guard4222;
wire _guard4224 = _guard4218 | _guard4223;
wire _guard4225 = fsm0_out == 2'd1;
wire _guard4226 = while_wrapper_early_reset_static_par0_done_out;
wire _guard4227 = _guard4225 & _guard4226;
wire _guard4228 = tdcc_go_out;
wire _guard4229 = _guard4227 & _guard4228;
wire _guard4230 = _guard4224 | _guard4229;
wire _guard4231 = fsm0_out == 2'd0;
wire _guard4232 = wrapper_early_reset_static_par_done_out;
wire _guard4233 = _guard4231 & _guard4232;
wire _guard4234 = tdcc_go_out;
wire _guard4235 = _guard4233 & _guard4234;
wire _guard4236 = fsm0_out == 2'd2;
wire _guard4237 = fsm0_out == 2'd1;
wire _guard4238 = while_wrapper_early_reset_static_par0_done_out;
wire _guard4239 = _guard4237 & _guard4238;
wire _guard4240 = tdcc_go_out;
wire _guard4241 = _guard4239 & _guard4240;
wire _guard4242 = early_reset_static_par0_go_out;
wire _guard4243 = early_reset_static_par0_go_out;
wire _guard4244 = early_reset_static_par0_go_out;
wire _guard4245 = early_reset_static_par0_go_out;
wire _guard4246 = early_reset_static_par0_go_out;
wire _guard4247 = early_reset_static_par0_go_out;
wire _guard4248 = early_reset_static_par0_go_out;
wire _guard4249 = early_reset_static_par0_go_out;
wire _guard4250 = cond_wire62_out;
wire _guard4251 = early_reset_static_par0_go_out;
wire _guard4252 = _guard4250 & _guard4251;
wire _guard4253 = cond_wire60_out;
wire _guard4254 = early_reset_static_par0_go_out;
wire _guard4255 = _guard4253 & _guard4254;
wire _guard4256 = fsm_out == 1'd0;
wire _guard4257 = cond_wire60_out;
wire _guard4258 = _guard4256 & _guard4257;
wire _guard4259 = fsm_out == 1'd0;
wire _guard4260 = _guard4258 & _guard4259;
wire _guard4261 = fsm_out == 1'd0;
wire _guard4262 = cond_wire62_out;
wire _guard4263 = _guard4261 & _guard4262;
wire _guard4264 = fsm_out == 1'd0;
wire _guard4265 = _guard4263 & _guard4264;
wire _guard4266 = _guard4260 | _guard4265;
wire _guard4267 = early_reset_static_par0_go_out;
wire _guard4268 = _guard4266 & _guard4267;
wire _guard4269 = fsm_out == 1'd0;
wire _guard4270 = cond_wire60_out;
wire _guard4271 = _guard4269 & _guard4270;
wire _guard4272 = fsm_out == 1'd0;
wire _guard4273 = _guard4271 & _guard4272;
wire _guard4274 = fsm_out == 1'd0;
wire _guard4275 = cond_wire62_out;
wire _guard4276 = _guard4274 & _guard4275;
wire _guard4277 = fsm_out == 1'd0;
wire _guard4278 = _guard4276 & _guard4277;
wire _guard4279 = _guard4273 | _guard4278;
wire _guard4280 = early_reset_static_par0_go_out;
wire _guard4281 = _guard4279 & _guard4280;
wire _guard4282 = fsm_out == 1'd0;
wire _guard4283 = cond_wire60_out;
wire _guard4284 = _guard4282 & _guard4283;
wire _guard4285 = fsm_out == 1'd0;
wire _guard4286 = _guard4284 & _guard4285;
wire _guard4287 = fsm_out == 1'd0;
wire _guard4288 = cond_wire62_out;
wire _guard4289 = _guard4287 & _guard4288;
wire _guard4290 = fsm_out == 1'd0;
wire _guard4291 = _guard4289 & _guard4290;
wire _guard4292 = _guard4286 | _guard4291;
wire _guard4293 = early_reset_static_par0_go_out;
wire _guard4294 = _guard4292 & _guard4293;
wire _guard4295 = cond_wire31_out;
wire _guard4296 = early_reset_static_par0_go_out;
wire _guard4297 = _guard4295 & _guard4296;
wire _guard4298 = cond_wire31_out;
wire _guard4299 = early_reset_static_par0_go_out;
wire _guard4300 = _guard4298 & _guard4299;
wire _guard4301 = cond_wire41_out;
wire _guard4302 = early_reset_static_par0_go_out;
wire _guard4303 = _guard4301 & _guard4302;
wire _guard4304 = cond_wire41_out;
wire _guard4305 = early_reset_static_par0_go_out;
wire _guard4306 = _guard4304 & _guard4305;
wire _guard4307 = cond_wire74_out;
wire _guard4308 = early_reset_static_par0_go_out;
wire _guard4309 = _guard4307 & _guard4308;
wire _guard4310 = cond_wire74_out;
wire _guard4311 = early_reset_static_par0_go_out;
wire _guard4312 = _guard4310 & _guard4311;
wire _guard4313 = cond_wire78_out;
wire _guard4314 = early_reset_static_par0_go_out;
wire _guard4315 = _guard4313 & _guard4314;
wire _guard4316 = cond_wire78_out;
wire _guard4317 = early_reset_static_par0_go_out;
wire _guard4318 = _guard4316 & _guard4317;
wire _guard4319 = cond_wire165_out;
wire _guard4320 = early_reset_static_par0_go_out;
wire _guard4321 = _guard4319 & _guard4320;
wire _guard4322 = cond_wire163_out;
wire _guard4323 = early_reset_static_par0_go_out;
wire _guard4324 = _guard4322 & _guard4323;
wire _guard4325 = fsm_out == 1'd0;
wire _guard4326 = cond_wire163_out;
wire _guard4327 = _guard4325 & _guard4326;
wire _guard4328 = fsm_out == 1'd0;
wire _guard4329 = _guard4327 & _guard4328;
wire _guard4330 = fsm_out == 1'd0;
wire _guard4331 = cond_wire165_out;
wire _guard4332 = _guard4330 & _guard4331;
wire _guard4333 = fsm_out == 1'd0;
wire _guard4334 = _guard4332 & _guard4333;
wire _guard4335 = _guard4329 | _guard4334;
wire _guard4336 = early_reset_static_par0_go_out;
wire _guard4337 = _guard4335 & _guard4336;
wire _guard4338 = fsm_out == 1'd0;
wire _guard4339 = cond_wire163_out;
wire _guard4340 = _guard4338 & _guard4339;
wire _guard4341 = fsm_out == 1'd0;
wire _guard4342 = _guard4340 & _guard4341;
wire _guard4343 = fsm_out == 1'd0;
wire _guard4344 = cond_wire165_out;
wire _guard4345 = _guard4343 & _guard4344;
wire _guard4346 = fsm_out == 1'd0;
wire _guard4347 = _guard4345 & _guard4346;
wire _guard4348 = _guard4342 | _guard4347;
wire _guard4349 = early_reset_static_par0_go_out;
wire _guard4350 = _guard4348 & _guard4349;
wire _guard4351 = fsm_out == 1'd0;
wire _guard4352 = cond_wire163_out;
wire _guard4353 = _guard4351 & _guard4352;
wire _guard4354 = fsm_out == 1'd0;
wire _guard4355 = _guard4353 & _guard4354;
wire _guard4356 = fsm_out == 1'd0;
wire _guard4357 = cond_wire165_out;
wire _guard4358 = _guard4356 & _guard4357;
wire _guard4359 = fsm_out == 1'd0;
wire _guard4360 = _guard4358 & _guard4359;
wire _guard4361 = _guard4355 | _guard4360;
wire _guard4362 = early_reset_static_par0_go_out;
wire _guard4363 = _guard4361 & _guard4362;
wire _guard4364 = cond_wire148_out;
wire _guard4365 = early_reset_static_par0_go_out;
wire _guard4366 = _guard4364 & _guard4365;
wire _guard4367 = cond_wire148_out;
wire _guard4368 = early_reset_static_par0_go_out;
wire _guard4369 = _guard4367 & _guard4368;
wire _guard4370 = cond_wire156_out;
wire _guard4371 = early_reset_static_par0_go_out;
wire _guard4372 = _guard4370 & _guard4371;
wire _guard4373 = cond_wire156_out;
wire _guard4374 = early_reset_static_par0_go_out;
wire _guard4375 = _guard4373 & _guard4374;
wire _guard4376 = cond_wire263_out;
wire _guard4377 = early_reset_static_par0_go_out;
wire _guard4378 = _guard4376 & _guard4377;
wire _guard4379 = cond_wire263_out;
wire _guard4380 = early_reset_static_par0_go_out;
wire _guard4381 = _guard4379 & _guard4380;
wire _guard4382 = cond_wire34_out;
wire _guard4383 = early_reset_static_par0_go_out;
wire _guard4384 = _guard4382 & _guard4383;
wire _guard4385 = cond_wire34_out;
wire _guard4386 = early_reset_static_par0_go_out;
wire _guard4387 = _guard4385 & _guard4386;
wire _guard4388 = early_reset_static_par_go_out;
wire _guard4389 = cond_wire138_out;
wire _guard4390 = early_reset_static_par0_go_out;
wire _guard4391 = _guard4389 & _guard4390;
wire _guard4392 = _guard4388 | _guard4391;
wire _guard4393 = early_reset_static_par_go_out;
wire _guard4394 = cond_wire138_out;
wire _guard4395 = early_reset_static_par0_go_out;
wire _guard4396 = _guard4394 & _guard4395;
wire _guard4397 = early_reset_static_par_go_out;
wire _guard4398 = early_reset_static_par0_go_out;
wire _guard4399 = _guard4397 | _guard4398;
wire _guard4400 = early_reset_static_par_go_out;
wire _guard4401 = early_reset_static_par0_go_out;
wire _guard4402 = early_reset_static_par_go_out;
wire _guard4403 = early_reset_static_par0_go_out;
wire _guard4404 = _guard4402 | _guard4403;
wire _guard4405 = early_reset_static_par0_go_out;
wire _guard4406 = early_reset_static_par_go_out;
wire _guard4407 = early_reset_static_par_go_out;
wire _guard4408 = early_reset_static_par0_go_out;
wire _guard4409 = _guard4407 | _guard4408;
wire _guard4410 = early_reset_static_par0_go_out;
wire _guard4411 = early_reset_static_par_go_out;
wire _guard4412 = early_reset_static_par0_go_out;
wire _guard4413 = early_reset_static_par0_go_out;
wire _guard4414 = early_reset_static_par_go_out;
wire _guard4415 = early_reset_static_par0_go_out;
wire _guard4416 = _guard4414 | _guard4415;
wire _guard4417 = early_reset_static_par_go_out;
wire _guard4418 = early_reset_static_par0_go_out;
wire _guard4419 = early_reset_static_par0_go_out;
wire _guard4420 = early_reset_static_par0_go_out;
wire _guard4421 = early_reset_static_par0_go_out;
wire _guard4422 = early_reset_static_par0_go_out;
wire _guard4423 = early_reset_static_par0_go_out;
wire _guard4424 = early_reset_static_par0_go_out;
wire _guard4425 = early_reset_static_par0_go_out;
wire _guard4426 = early_reset_static_par0_go_out;
wire _guard4427 = early_reset_static_par0_go_out;
wire _guard4428 = early_reset_static_par0_go_out;
wire _guard4429 = early_reset_static_par_go_out;
wire _guard4430 = early_reset_static_par0_go_out;
wire _guard4431 = _guard4429 | _guard4430;
wire _guard4432 = early_reset_static_par_go_out;
wire _guard4433 = early_reset_static_par0_go_out;
wire _guard4434 = early_reset_static_par0_go_out;
wire _guard4435 = early_reset_static_par0_go_out;
wire _guard4436 = early_reset_static_par0_go_out;
wire _guard4437 = early_reset_static_par0_go_out;
wire _guard4438 = early_reset_static_par0_go_out;
wire _guard4439 = early_reset_static_par0_go_out;
wire _guard4440 = early_reset_static_par0_go_out;
wire _guard4441 = early_reset_static_par0_go_out;
wire _guard4442 = early_reset_static_par0_go_out;
wire _guard4443 = early_reset_static_par0_go_out;
wire _guard4444 = early_reset_static_par0_go_out;
wire _guard4445 = ~_guard0;
wire _guard4446 = early_reset_static_par0_go_out;
wire _guard4447 = _guard4445 & _guard4446;
wire _guard4448 = early_reset_static_par0_go_out;
wire _guard4449 = early_reset_static_par0_go_out;
wire _guard4450 = early_reset_static_par0_go_out;
wire _guard4451 = early_reset_static_par0_go_out;
wire _guard4452 = early_reset_static_par0_go_out;
wire _guard4453 = ~_guard0;
wire _guard4454 = early_reset_static_par0_go_out;
wire _guard4455 = _guard4453 & _guard4454;
wire _guard4456 = early_reset_static_par0_go_out;
wire _guard4457 = early_reset_static_par0_go_out;
wire _guard4458 = early_reset_static_par0_go_out;
wire _guard4459 = early_reset_static_par0_go_out;
wire _guard4460 = early_reset_static_par0_go_out;
wire _guard4461 = ~_guard0;
wire _guard4462 = early_reset_static_par0_go_out;
wire _guard4463 = _guard4461 & _guard4462;
wire _guard4464 = early_reset_static_par0_go_out;
wire _guard4465 = early_reset_static_par0_go_out;
wire _guard4466 = ~_guard0;
wire _guard4467 = early_reset_static_par0_go_out;
wire _guard4468 = _guard4466 & _guard4467;
wire _guard4469 = early_reset_static_par0_go_out;
wire _guard4470 = early_reset_static_par0_go_out;
wire _guard4471 = ~_guard0;
wire _guard4472 = early_reset_static_par0_go_out;
wire _guard4473 = _guard4471 & _guard4472;
wire _guard4474 = ~_guard0;
wire _guard4475 = early_reset_static_par0_go_out;
wire _guard4476 = _guard4474 & _guard4475;
wire _guard4477 = early_reset_static_par0_go_out;
wire _guard4478 = ~_guard0;
wire _guard4479 = early_reset_static_par0_go_out;
wire _guard4480 = _guard4478 & _guard4479;
wire _guard4481 = early_reset_static_par0_go_out;
wire _guard4482 = early_reset_static_par0_go_out;
wire _guard4483 = early_reset_static_par0_go_out;
wire _guard4484 = ~_guard0;
wire _guard4485 = early_reset_static_par0_go_out;
wire _guard4486 = _guard4484 & _guard4485;
wire _guard4487 = early_reset_static_par0_go_out;
wire _guard4488 = early_reset_static_par0_go_out;
wire _guard4489 = ~_guard0;
wire _guard4490 = early_reset_static_par0_go_out;
wire _guard4491 = _guard4489 & _guard4490;
wire _guard4492 = early_reset_static_par0_go_out;
wire _guard4493 = early_reset_static_par0_go_out;
wire _guard4494 = ~_guard0;
wire _guard4495 = early_reset_static_par0_go_out;
wire _guard4496 = _guard4494 & _guard4495;
wire _guard4497 = early_reset_static_par0_go_out;
wire _guard4498 = early_reset_static_par0_go_out;
wire _guard4499 = early_reset_static_par0_go_out;
wire _guard4500 = early_reset_static_par0_go_out;
wire _guard4501 = ~_guard0;
wire _guard4502 = early_reset_static_par0_go_out;
wire _guard4503 = _guard4501 & _guard4502;
wire _guard4504 = early_reset_static_par0_go_out;
wire _guard4505 = ~_guard0;
wire _guard4506 = early_reset_static_par0_go_out;
wire _guard4507 = _guard4505 & _guard4506;
wire _guard4508 = ~_guard0;
wire _guard4509 = early_reset_static_par0_go_out;
wire _guard4510 = _guard4508 & _guard4509;
wire _guard4511 = early_reset_static_par0_go_out;
wire _guard4512 = early_reset_static_par0_go_out;
wire _guard4513 = ~_guard0;
wire _guard4514 = early_reset_static_par0_go_out;
wire _guard4515 = _guard4513 & _guard4514;
wire _guard4516 = early_reset_static_par0_go_out;
wire _guard4517 = early_reset_static_par0_go_out;
wire _guard4518 = early_reset_static_par0_go_out;
wire _guard4519 = early_reset_static_par0_go_out;
wire _guard4520 = early_reset_static_par0_go_out;
wire _guard4521 = early_reset_static_par0_go_out;
wire _guard4522 = ~_guard0;
wire _guard4523 = early_reset_static_par0_go_out;
wire _guard4524 = _guard4522 & _guard4523;
wire _guard4525 = early_reset_static_par0_go_out;
wire _guard4526 = ~_guard0;
wire _guard4527 = early_reset_static_par0_go_out;
wire _guard4528 = _guard4526 & _guard4527;
wire _guard4529 = early_reset_static_par0_go_out;
wire _guard4530 = early_reset_static_par0_go_out;
wire _guard4531 = early_reset_static_par0_go_out;
wire _guard4532 = early_reset_static_par0_go_out;
wire _guard4533 = early_reset_static_par0_go_out;
wire _guard4534 = early_reset_static_par0_go_out;
wire _guard4535 = early_reset_static_par0_go_out;
wire _guard4536 = early_reset_static_par0_go_out;
wire _guard4537 = ~_guard0;
wire _guard4538 = early_reset_static_par0_go_out;
wire _guard4539 = _guard4537 & _guard4538;
wire _guard4540 = early_reset_static_par0_go_out;
wire _guard4541 = ~_guard0;
wire _guard4542 = early_reset_static_par0_go_out;
wire _guard4543 = _guard4541 & _guard4542;
wire _guard4544 = early_reset_static_par0_go_out;
wire _guard4545 = early_reset_static_par0_go_out;
wire _guard4546 = early_reset_static_par0_go_out;
wire _guard4547 = early_reset_static_par0_go_out;
wire _guard4548 = early_reset_static_par0_go_out;
wire _guard4549 = early_reset_static_par0_go_out;
wire _guard4550 = early_reset_static_par0_go_out;
wire _guard4551 = early_reset_static_par0_go_out;
wire _guard4552 = early_reset_static_par_go_out;
wire _guard4553 = lt_iter_limit_out;
wire _guard4554 = early_reset_static_par_go_out;
wire _guard4555 = _guard4553 & _guard4554;
wire _guard4556 = lt_iter_limit_out;
wire _guard4557 = ~_guard4556;
wire _guard4558 = early_reset_static_par_go_out;
wire _guard4559 = _guard4557 & _guard4558;
wire _guard4560 = early_reset_static_par0_go_out;
wire _guard4561 = early_reset_static_par0_go_out;
wire _guard4562 = early_reset_static_par0_go_out;
wire _guard4563 = early_reset_static_par0_go_out;
wire _guard4564 = early_reset_static_par0_go_out;
wire _guard4565 = early_reset_static_par0_go_out;
wire _guard4566 = cond_wire4_out;
wire _guard4567 = early_reset_static_par0_go_out;
wire _guard4568 = _guard4566 & _guard4567;
wire _guard4569 = cond_wire4_out;
wire _guard4570 = early_reset_static_par0_go_out;
wire _guard4571 = _guard4569 & _guard4570;
wire _guard4572 = cond_wire6_out;
wire _guard4573 = early_reset_static_par0_go_out;
wire _guard4574 = _guard4572 & _guard4573;
wire _guard4575 = cond_wire6_out;
wire _guard4576 = early_reset_static_par0_go_out;
wire _guard4577 = _guard4575 & _guard4576;
wire _guard4578 = cond_wire22_out;
wire _guard4579 = early_reset_static_par0_go_out;
wire _guard4580 = _guard4578 & _guard4579;
wire _guard4581 = cond_wire20_out;
wire _guard4582 = early_reset_static_par0_go_out;
wire _guard4583 = _guard4581 & _guard4582;
wire _guard4584 = fsm_out == 1'd0;
wire _guard4585 = cond_wire20_out;
wire _guard4586 = _guard4584 & _guard4585;
wire _guard4587 = fsm_out == 1'd0;
wire _guard4588 = _guard4586 & _guard4587;
wire _guard4589 = fsm_out == 1'd0;
wire _guard4590 = cond_wire22_out;
wire _guard4591 = _guard4589 & _guard4590;
wire _guard4592 = fsm_out == 1'd0;
wire _guard4593 = _guard4591 & _guard4592;
wire _guard4594 = _guard4588 | _guard4593;
wire _guard4595 = early_reset_static_par0_go_out;
wire _guard4596 = _guard4594 & _guard4595;
wire _guard4597 = fsm_out == 1'd0;
wire _guard4598 = cond_wire20_out;
wire _guard4599 = _guard4597 & _guard4598;
wire _guard4600 = fsm_out == 1'd0;
wire _guard4601 = _guard4599 & _guard4600;
wire _guard4602 = fsm_out == 1'd0;
wire _guard4603 = cond_wire22_out;
wire _guard4604 = _guard4602 & _guard4603;
wire _guard4605 = fsm_out == 1'd0;
wire _guard4606 = _guard4604 & _guard4605;
wire _guard4607 = _guard4601 | _guard4606;
wire _guard4608 = early_reset_static_par0_go_out;
wire _guard4609 = _guard4607 & _guard4608;
wire _guard4610 = fsm_out == 1'd0;
wire _guard4611 = cond_wire20_out;
wire _guard4612 = _guard4610 & _guard4611;
wire _guard4613 = fsm_out == 1'd0;
wire _guard4614 = _guard4612 & _guard4613;
wire _guard4615 = fsm_out == 1'd0;
wire _guard4616 = cond_wire22_out;
wire _guard4617 = _guard4615 & _guard4616;
wire _guard4618 = fsm_out == 1'd0;
wire _guard4619 = _guard4617 & _guard4618;
wire _guard4620 = _guard4614 | _guard4619;
wire _guard4621 = early_reset_static_par0_go_out;
wire _guard4622 = _guard4620 & _guard4621;
wire _guard4623 = cond_wire53_out;
wire _guard4624 = early_reset_static_par0_go_out;
wire _guard4625 = _guard4623 & _guard4624;
wire _guard4626 = cond_wire53_out;
wire _guard4627 = early_reset_static_par0_go_out;
wire _guard4628 = _guard4626 & _guard4627;
wire _guard4629 = cond_wire99_out;
wire _guard4630 = early_reset_static_par0_go_out;
wire _guard4631 = _guard4629 & _guard4630;
wire _guard4632 = cond_wire97_out;
wire _guard4633 = early_reset_static_par0_go_out;
wire _guard4634 = _guard4632 & _guard4633;
wire _guard4635 = fsm_out == 1'd0;
wire _guard4636 = cond_wire97_out;
wire _guard4637 = _guard4635 & _guard4636;
wire _guard4638 = fsm_out == 1'd0;
wire _guard4639 = _guard4637 & _guard4638;
wire _guard4640 = fsm_out == 1'd0;
wire _guard4641 = cond_wire99_out;
wire _guard4642 = _guard4640 & _guard4641;
wire _guard4643 = fsm_out == 1'd0;
wire _guard4644 = _guard4642 & _guard4643;
wire _guard4645 = _guard4639 | _guard4644;
wire _guard4646 = early_reset_static_par0_go_out;
wire _guard4647 = _guard4645 & _guard4646;
wire _guard4648 = fsm_out == 1'd0;
wire _guard4649 = cond_wire97_out;
wire _guard4650 = _guard4648 & _guard4649;
wire _guard4651 = fsm_out == 1'd0;
wire _guard4652 = _guard4650 & _guard4651;
wire _guard4653 = fsm_out == 1'd0;
wire _guard4654 = cond_wire99_out;
wire _guard4655 = _guard4653 & _guard4654;
wire _guard4656 = fsm_out == 1'd0;
wire _guard4657 = _guard4655 & _guard4656;
wire _guard4658 = _guard4652 | _guard4657;
wire _guard4659 = early_reset_static_par0_go_out;
wire _guard4660 = _guard4658 & _guard4659;
wire _guard4661 = fsm_out == 1'd0;
wire _guard4662 = cond_wire97_out;
wire _guard4663 = _guard4661 & _guard4662;
wire _guard4664 = fsm_out == 1'd0;
wire _guard4665 = _guard4663 & _guard4664;
wire _guard4666 = fsm_out == 1'd0;
wire _guard4667 = cond_wire99_out;
wire _guard4668 = _guard4666 & _guard4667;
wire _guard4669 = fsm_out == 1'd0;
wire _guard4670 = _guard4668 & _guard4669;
wire _guard4671 = _guard4665 | _guard4670;
wire _guard4672 = early_reset_static_par0_go_out;
wire _guard4673 = _guard4671 & _guard4672;
wire _guard4674 = cond_wire105_out;
wire _guard4675 = early_reset_static_par0_go_out;
wire _guard4676 = _guard4674 & _guard4675;
wire _guard4677 = cond_wire105_out;
wire _guard4678 = early_reset_static_par0_go_out;
wire _guard4679 = _guard4677 & _guard4678;
wire _guard4680 = cond_wire149_out;
wire _guard4681 = early_reset_static_par0_go_out;
wire _guard4682 = _guard4680 & _guard4681;
wire _guard4683 = cond_wire147_out;
wire _guard4684 = early_reset_static_par0_go_out;
wire _guard4685 = _guard4683 & _guard4684;
wire _guard4686 = fsm_out == 1'd0;
wire _guard4687 = cond_wire147_out;
wire _guard4688 = _guard4686 & _guard4687;
wire _guard4689 = fsm_out == 1'd0;
wire _guard4690 = _guard4688 & _guard4689;
wire _guard4691 = fsm_out == 1'd0;
wire _guard4692 = cond_wire149_out;
wire _guard4693 = _guard4691 & _guard4692;
wire _guard4694 = fsm_out == 1'd0;
wire _guard4695 = _guard4693 & _guard4694;
wire _guard4696 = _guard4690 | _guard4695;
wire _guard4697 = early_reset_static_par0_go_out;
wire _guard4698 = _guard4696 & _guard4697;
wire _guard4699 = fsm_out == 1'd0;
wire _guard4700 = cond_wire147_out;
wire _guard4701 = _guard4699 & _guard4700;
wire _guard4702 = fsm_out == 1'd0;
wire _guard4703 = _guard4701 & _guard4702;
wire _guard4704 = fsm_out == 1'd0;
wire _guard4705 = cond_wire149_out;
wire _guard4706 = _guard4704 & _guard4705;
wire _guard4707 = fsm_out == 1'd0;
wire _guard4708 = _guard4706 & _guard4707;
wire _guard4709 = _guard4703 | _guard4708;
wire _guard4710 = early_reset_static_par0_go_out;
wire _guard4711 = _guard4709 & _guard4710;
wire _guard4712 = fsm_out == 1'd0;
wire _guard4713 = cond_wire147_out;
wire _guard4714 = _guard4712 & _guard4713;
wire _guard4715 = fsm_out == 1'd0;
wire _guard4716 = _guard4714 & _guard4715;
wire _guard4717 = fsm_out == 1'd0;
wire _guard4718 = cond_wire149_out;
wire _guard4719 = _guard4717 & _guard4718;
wire _guard4720 = fsm_out == 1'd0;
wire _guard4721 = _guard4719 & _guard4720;
wire _guard4722 = _guard4716 | _guard4721;
wire _guard4723 = early_reset_static_par0_go_out;
wire _guard4724 = _guard4722 & _guard4723;
wire _guard4725 = cond_wire144_out;
wire _guard4726 = early_reset_static_par0_go_out;
wire _guard4727 = _guard4725 & _guard4726;
wire _guard4728 = cond_wire144_out;
wire _guard4729 = early_reset_static_par0_go_out;
wire _guard4730 = _guard4728 & _guard4729;
wire _guard4731 = cond_wire185_out;
wire _guard4732 = early_reset_static_par0_go_out;
wire _guard4733 = _guard4731 & _guard4732;
wire _guard4734 = cond_wire185_out;
wire _guard4735 = early_reset_static_par0_go_out;
wire _guard4736 = _guard4734 & _guard4735;
wire _guard4737 = cond_wire235_out;
wire _guard4738 = early_reset_static_par0_go_out;
wire _guard4739 = _guard4737 & _guard4738;
wire _guard4740 = cond_wire233_out;
wire _guard4741 = early_reset_static_par0_go_out;
wire _guard4742 = _guard4740 & _guard4741;
wire _guard4743 = fsm_out == 1'd0;
wire _guard4744 = cond_wire233_out;
wire _guard4745 = _guard4743 & _guard4744;
wire _guard4746 = fsm_out == 1'd0;
wire _guard4747 = _guard4745 & _guard4746;
wire _guard4748 = fsm_out == 1'd0;
wire _guard4749 = cond_wire235_out;
wire _guard4750 = _guard4748 & _guard4749;
wire _guard4751 = fsm_out == 1'd0;
wire _guard4752 = _guard4750 & _guard4751;
wire _guard4753 = _guard4747 | _guard4752;
wire _guard4754 = early_reset_static_par0_go_out;
wire _guard4755 = _guard4753 & _guard4754;
wire _guard4756 = fsm_out == 1'd0;
wire _guard4757 = cond_wire233_out;
wire _guard4758 = _guard4756 & _guard4757;
wire _guard4759 = fsm_out == 1'd0;
wire _guard4760 = _guard4758 & _guard4759;
wire _guard4761 = fsm_out == 1'd0;
wire _guard4762 = cond_wire235_out;
wire _guard4763 = _guard4761 & _guard4762;
wire _guard4764 = fsm_out == 1'd0;
wire _guard4765 = _guard4763 & _guard4764;
wire _guard4766 = _guard4760 | _guard4765;
wire _guard4767 = early_reset_static_par0_go_out;
wire _guard4768 = _guard4766 & _guard4767;
wire _guard4769 = fsm_out == 1'd0;
wire _guard4770 = cond_wire233_out;
wire _guard4771 = _guard4769 & _guard4770;
wire _guard4772 = fsm_out == 1'd0;
wire _guard4773 = _guard4771 & _guard4772;
wire _guard4774 = fsm_out == 1'd0;
wire _guard4775 = cond_wire235_out;
wire _guard4776 = _guard4774 & _guard4775;
wire _guard4777 = fsm_out == 1'd0;
wire _guard4778 = _guard4776 & _guard4777;
wire _guard4779 = _guard4773 | _guard4778;
wire _guard4780 = early_reset_static_par0_go_out;
wire _guard4781 = _guard4779 & _guard4780;
wire _guard4782 = cond_wire237_out;
wire _guard4783 = early_reset_static_par0_go_out;
wire _guard4784 = _guard4782 & _guard4783;
wire _guard4785 = cond_wire237_out;
wire _guard4786 = early_reset_static_par0_go_out;
wire _guard4787 = _guard4785 & _guard4786;
wire _guard4788 = early_reset_static_par0_go_out;
wire _guard4789 = early_reset_static_par0_go_out;
wire _guard4790 = early_reset_static_par0_go_out;
wire _guard4791 = early_reset_static_par0_go_out;
wire _guard4792 = early_reset_static_par0_go_out;
wire _guard4793 = early_reset_static_par0_go_out;
wire _guard4794 = early_reset_static_par_go_out;
wire _guard4795 = early_reset_static_par0_go_out;
wire _guard4796 = _guard4794 | _guard4795;
wire _guard4797 = early_reset_static_par0_go_out;
wire _guard4798 = early_reset_static_par_go_out;
wire _guard4799 = early_reset_static_par0_go_out;
wire _guard4800 = early_reset_static_par0_go_out;
wire _guard4801 = early_reset_static_par0_go_out;
wire _guard4802 = early_reset_static_par0_go_out;
wire _guard4803 = early_reset_static_par_go_out;
wire _guard4804 = early_reset_static_par0_go_out;
wire _guard4805 = _guard4803 | _guard4804;
wire _guard4806 = early_reset_static_par_go_out;
wire _guard4807 = early_reset_static_par0_go_out;
wire _guard4808 = early_reset_static_par0_go_out;
wire _guard4809 = early_reset_static_par0_go_out;
wire _guard4810 = early_reset_static_par_go_out;
wire _guard4811 = early_reset_static_par0_go_out;
wire _guard4812 = _guard4810 | _guard4811;
wire _guard4813 = early_reset_static_par_go_out;
wire _guard4814 = early_reset_static_par0_go_out;
wire _guard4815 = early_reset_static_par0_go_out;
wire _guard4816 = early_reset_static_par0_go_out;
wire _guard4817 = early_reset_static_par0_go_out;
wire _guard4818 = early_reset_static_par0_go_out;
wire _guard4819 = ~_guard0;
wire _guard4820 = early_reset_static_par0_go_out;
wire _guard4821 = _guard4819 & _guard4820;
wire _guard4822 = early_reset_static_par0_go_out;
wire _guard4823 = early_reset_static_par0_go_out;
wire _guard4824 = early_reset_static_par0_go_out;
wire _guard4825 = ~_guard0;
wire _guard4826 = early_reset_static_par0_go_out;
wire _guard4827 = _guard4825 & _guard4826;
wire _guard4828 = early_reset_static_par0_go_out;
wire _guard4829 = early_reset_static_par0_go_out;
wire _guard4830 = early_reset_static_par0_go_out;
wire _guard4831 = early_reset_static_par0_go_out;
wire _guard4832 = ~_guard0;
wire _guard4833 = early_reset_static_par0_go_out;
wire _guard4834 = _guard4832 & _guard4833;
wire _guard4835 = early_reset_static_par0_go_out;
wire _guard4836 = early_reset_static_par0_go_out;
wire _guard4837 = early_reset_static_par0_go_out;
wire _guard4838 = ~_guard0;
wire _guard4839 = early_reset_static_par0_go_out;
wire _guard4840 = _guard4838 & _guard4839;
wire _guard4841 = ~_guard0;
wire _guard4842 = early_reset_static_par0_go_out;
wire _guard4843 = _guard4841 & _guard4842;
wire _guard4844 = early_reset_static_par0_go_out;
wire _guard4845 = ~_guard0;
wire _guard4846 = early_reset_static_par0_go_out;
wire _guard4847 = _guard4845 & _guard4846;
wire _guard4848 = early_reset_static_par0_go_out;
wire _guard4849 = early_reset_static_par0_go_out;
wire _guard4850 = early_reset_static_par0_go_out;
wire _guard4851 = early_reset_static_par0_go_out;
wire _guard4852 = early_reset_static_par0_go_out;
wire _guard4853 = ~_guard0;
wire _guard4854 = early_reset_static_par0_go_out;
wire _guard4855 = _guard4853 & _guard4854;
wire _guard4856 = early_reset_static_par0_go_out;
wire _guard4857 = early_reset_static_par0_go_out;
wire _guard4858 = early_reset_static_par0_go_out;
wire _guard4859 = early_reset_static_par0_go_out;
wire _guard4860 = early_reset_static_par0_go_out;
wire _guard4861 = early_reset_static_par0_go_out;
wire _guard4862 = ~_guard0;
wire _guard4863 = early_reset_static_par0_go_out;
wire _guard4864 = _guard4862 & _guard4863;
wire _guard4865 = early_reset_static_par0_go_out;
wire _guard4866 = early_reset_static_par0_go_out;
wire _guard4867 = early_reset_static_par0_go_out;
wire _guard4868 = early_reset_static_par0_go_out;
wire _guard4869 = early_reset_static_par0_go_out;
wire _guard4870 = ~_guard0;
wire _guard4871 = early_reset_static_par0_go_out;
wire _guard4872 = _guard4870 & _guard4871;
wire _guard4873 = early_reset_static_par0_go_out;
wire _guard4874 = ~_guard0;
wire _guard4875 = early_reset_static_par0_go_out;
wire _guard4876 = _guard4874 & _guard4875;
wire _guard4877 = ~_guard0;
wire _guard4878 = early_reset_static_par0_go_out;
wire _guard4879 = _guard4877 & _guard4878;
wire _guard4880 = early_reset_static_par0_go_out;
wire _guard4881 = early_reset_static_par0_go_out;
wire _guard4882 = early_reset_static_par0_go_out;
wire _guard4883 = early_reset_static_par0_go_out;
wire _guard4884 = ~_guard0;
wire _guard4885 = early_reset_static_par0_go_out;
wire _guard4886 = _guard4884 & _guard4885;
wire _guard4887 = early_reset_static_par0_go_out;
wire _guard4888 = early_reset_static_par0_go_out;
wire _guard4889 = early_reset_static_par0_go_out;
wire _guard4890 = early_reset_static_par0_go_out;
wire _guard4891 = early_reset_static_par0_go_out;
wire _guard4892 = ~_guard0;
wire _guard4893 = early_reset_static_par0_go_out;
wire _guard4894 = _guard4892 & _guard4893;
wire _guard4895 = early_reset_static_par0_go_out;
wire _guard4896 = ~_guard0;
wire _guard4897 = early_reset_static_par0_go_out;
wire _guard4898 = _guard4896 & _guard4897;
wire _guard4899 = ~_guard0;
wire _guard4900 = early_reset_static_par0_go_out;
wire _guard4901 = _guard4899 & _guard4900;
wire _guard4902 = early_reset_static_par0_go_out;
wire _guard4903 = ~_guard0;
wire _guard4904 = early_reset_static_par0_go_out;
wire _guard4905 = _guard4903 & _guard4904;
wire _guard4906 = early_reset_static_par0_go_out;
wire _guard4907 = early_reset_static_par0_go_out;
wire _guard4908 = early_reset_static_par0_go_out;
wire _guard4909 = early_reset_static_par0_go_out;
wire _guard4910 = early_reset_static_par0_go_out;
wire _guard4911 = early_reset_static_par0_go_out;
wire _guard4912 = early_reset_static_par0_go_out;
wire _guard4913 = ~_guard0;
wire _guard4914 = early_reset_static_par0_go_out;
wire _guard4915 = _guard4913 & _guard4914;
wire _guard4916 = early_reset_static_par0_go_out;
wire _guard4917 = early_reset_static_par0_go_out;
wire _guard4918 = early_reset_static_par0_go_out;
wire _guard4919 = early_reset_static_par0_go_out;
wire _guard4920 = ~_guard0;
wire _guard4921 = early_reset_static_par0_go_out;
wire _guard4922 = _guard4920 & _guard4921;
wire _guard4923 = ~_guard0;
wire _guard4924 = early_reset_static_par0_go_out;
wire _guard4925 = _guard4923 & _guard4924;
wire _guard4926 = early_reset_static_par0_go_out;
wire _guard4927 = early_reset_static_par0_go_out;
wire _guard4928 = ~_guard0;
wire _guard4929 = early_reset_static_par0_go_out;
wire _guard4930 = _guard4928 & _guard4929;
wire _guard4931 = early_reset_static_par0_go_out;
wire _guard4932 = early_reset_static_par0_go_out;
wire _guard4933 = ~_guard0;
wire _guard4934 = early_reset_static_par0_go_out;
wire _guard4935 = _guard4933 & _guard4934;
wire _guard4936 = early_reset_static_par0_go_out;
wire _guard4937 = early_reset_static_par0_go_out;
wire _guard4938 = early_reset_static_par0_go_out;
wire _guard4939 = early_reset_static_par0_go_out;
wire _guard4940 = early_reset_static_par0_go_out;
wire _guard4941 = early_reset_static_par0_go_out;
wire _guard4942 = ~_guard0;
wire _guard4943 = early_reset_static_par0_go_out;
wire _guard4944 = _guard4942 & _guard4943;
wire _guard4945 = early_reset_static_par0_go_out;
wire _guard4946 = ~_guard0;
wire _guard4947 = early_reset_static_par0_go_out;
wire _guard4948 = _guard4946 & _guard4947;
wire _guard4949 = early_reset_static_par0_go_out;
wire _guard4950 = ~_guard0;
wire _guard4951 = early_reset_static_par0_go_out;
wire _guard4952 = _guard4950 & _guard4951;
wire _guard4953 = early_reset_static_par0_go_out;
wire _guard4954 = ~_guard0;
wire _guard4955 = early_reset_static_par0_go_out;
wire _guard4956 = _guard4954 & _guard4955;
wire _guard4957 = early_reset_static_par0_go_out;
wire _guard4958 = early_reset_static_par0_go_out;
wire _guard4959 = early_reset_static_par0_go_out;
wire _guard4960 = early_reset_static_par0_go_out;
wire _guard4961 = early_reset_static_par0_go_out;
wire _guard4962 = early_reset_static_par0_go_out;
wire _guard4963 = cond_wire9_out;
wire _guard4964 = early_reset_static_par0_go_out;
wire _guard4965 = _guard4963 & _guard4964;
wire _guard4966 = cond_wire9_out;
wire _guard4967 = early_reset_static_par0_go_out;
wire _guard4968 = _guard4966 & _guard4967;
wire _guard4969 = cond_wire6_out;
wire _guard4970 = early_reset_static_par0_go_out;
wire _guard4971 = _guard4969 & _guard4970;
wire _guard4972 = cond_wire6_out;
wire _guard4973 = early_reset_static_par0_go_out;
wire _guard4974 = _guard4972 & _guard4973;
wire _guard4975 = cond_wire111_out;
wire _guard4976 = early_reset_static_par0_go_out;
wire _guard4977 = _guard4975 & _guard4976;
wire _guard4978 = cond_wire111_out;
wire _guard4979 = early_reset_static_par0_go_out;
wire _guard4980 = _guard4978 & _guard4979;
wire _guard4981 = cond_wire119_out;
wire _guard4982 = early_reset_static_par0_go_out;
wire _guard4983 = _guard4981 & _guard4982;
wire _guard4984 = cond_wire119_out;
wire _guard4985 = early_reset_static_par0_go_out;
wire _guard4986 = _guard4984 & _guard4985;
wire _guard4987 = cond_wire111_out;
wire _guard4988 = early_reset_static_par0_go_out;
wire _guard4989 = _guard4987 & _guard4988;
wire _guard4990 = cond_wire111_out;
wire _guard4991 = early_reset_static_par0_go_out;
wire _guard4992 = _guard4990 & _guard4991;
wire _guard4993 = cond_wire115_out;
wire _guard4994 = early_reset_static_par0_go_out;
wire _guard4995 = _guard4993 & _guard4994;
wire _guard4996 = cond_wire115_out;
wire _guard4997 = early_reset_static_par0_go_out;
wire _guard4998 = _guard4996 & _guard4997;
wire _guard4999 = cond_wire189_out;
wire _guard5000 = early_reset_static_par0_go_out;
wire _guard5001 = _guard4999 & _guard5000;
wire _guard5002 = cond_wire189_out;
wire _guard5003 = early_reset_static_par0_go_out;
wire _guard5004 = _guard5002 & _guard5003;
wire _guard5005 = cond_wire193_out;
wire _guard5006 = early_reset_static_par0_go_out;
wire _guard5007 = _guard5005 & _guard5006;
wire _guard5008 = cond_wire193_out;
wire _guard5009 = early_reset_static_par0_go_out;
wire _guard5010 = _guard5008 & _guard5009;
wire _guard5011 = cond_wire226_out;
wire _guard5012 = early_reset_static_par0_go_out;
wire _guard5013 = _guard5011 & _guard5012;
wire _guard5014 = cond_wire226_out;
wire _guard5015 = early_reset_static_par0_go_out;
wire _guard5016 = _guard5014 & _guard5015;
wire _guard5017 = cond_wire243_out;
wire _guard5018 = early_reset_static_par0_go_out;
wire _guard5019 = _guard5017 & _guard5018;
wire _guard5020 = cond_wire243_out;
wire _guard5021 = early_reset_static_par0_go_out;
wire _guard5022 = _guard5020 & _guard5021;
wire _guard5023 = cond_wire260_out;
wire _guard5024 = early_reset_static_par0_go_out;
wire _guard5025 = _guard5023 & _guard5024;
wire _guard5026 = cond_wire258_out;
wire _guard5027 = early_reset_static_par0_go_out;
wire _guard5028 = _guard5026 & _guard5027;
wire _guard5029 = fsm_out == 1'd0;
wire _guard5030 = cond_wire258_out;
wire _guard5031 = _guard5029 & _guard5030;
wire _guard5032 = fsm_out == 1'd0;
wire _guard5033 = _guard5031 & _guard5032;
wire _guard5034 = fsm_out == 1'd0;
wire _guard5035 = cond_wire260_out;
wire _guard5036 = _guard5034 & _guard5035;
wire _guard5037 = fsm_out == 1'd0;
wire _guard5038 = _guard5036 & _guard5037;
wire _guard5039 = _guard5033 | _guard5038;
wire _guard5040 = early_reset_static_par0_go_out;
wire _guard5041 = _guard5039 & _guard5040;
wire _guard5042 = fsm_out == 1'd0;
wire _guard5043 = cond_wire258_out;
wire _guard5044 = _guard5042 & _guard5043;
wire _guard5045 = fsm_out == 1'd0;
wire _guard5046 = _guard5044 & _guard5045;
wire _guard5047 = fsm_out == 1'd0;
wire _guard5048 = cond_wire260_out;
wire _guard5049 = _guard5047 & _guard5048;
wire _guard5050 = fsm_out == 1'd0;
wire _guard5051 = _guard5049 & _guard5050;
wire _guard5052 = _guard5046 | _guard5051;
wire _guard5053 = early_reset_static_par0_go_out;
wire _guard5054 = _guard5052 & _guard5053;
wire _guard5055 = fsm_out == 1'd0;
wire _guard5056 = cond_wire258_out;
wire _guard5057 = _guard5055 & _guard5056;
wire _guard5058 = fsm_out == 1'd0;
wire _guard5059 = _guard5057 & _guard5058;
wire _guard5060 = fsm_out == 1'd0;
wire _guard5061 = cond_wire260_out;
wire _guard5062 = _guard5060 & _guard5061;
wire _guard5063 = fsm_out == 1'd0;
wire _guard5064 = _guard5062 & _guard5063;
wire _guard5065 = _guard5059 | _guard5064;
wire _guard5066 = early_reset_static_par0_go_out;
wire _guard5067 = _guard5065 & _guard5066;
wire _guard5068 = cond_wire264_out;
wire _guard5069 = early_reset_static_par0_go_out;
wire _guard5070 = _guard5068 & _guard5069;
wire _guard5071 = cond_wire262_out;
wire _guard5072 = early_reset_static_par0_go_out;
wire _guard5073 = _guard5071 & _guard5072;
wire _guard5074 = fsm_out == 1'd0;
wire _guard5075 = cond_wire262_out;
wire _guard5076 = _guard5074 & _guard5075;
wire _guard5077 = fsm_out == 1'd0;
wire _guard5078 = _guard5076 & _guard5077;
wire _guard5079 = fsm_out == 1'd0;
wire _guard5080 = cond_wire264_out;
wire _guard5081 = _guard5079 & _guard5080;
wire _guard5082 = fsm_out == 1'd0;
wire _guard5083 = _guard5081 & _guard5082;
wire _guard5084 = _guard5078 | _guard5083;
wire _guard5085 = early_reset_static_par0_go_out;
wire _guard5086 = _guard5084 & _guard5085;
wire _guard5087 = fsm_out == 1'd0;
wire _guard5088 = cond_wire262_out;
wire _guard5089 = _guard5087 & _guard5088;
wire _guard5090 = fsm_out == 1'd0;
wire _guard5091 = _guard5089 & _guard5090;
wire _guard5092 = fsm_out == 1'd0;
wire _guard5093 = cond_wire264_out;
wire _guard5094 = _guard5092 & _guard5093;
wire _guard5095 = fsm_out == 1'd0;
wire _guard5096 = _guard5094 & _guard5095;
wire _guard5097 = _guard5091 | _guard5096;
wire _guard5098 = early_reset_static_par0_go_out;
wire _guard5099 = _guard5097 & _guard5098;
wire _guard5100 = fsm_out == 1'd0;
wire _guard5101 = cond_wire262_out;
wire _guard5102 = _guard5100 & _guard5101;
wire _guard5103 = fsm_out == 1'd0;
wire _guard5104 = _guard5102 & _guard5103;
wire _guard5105 = fsm_out == 1'd0;
wire _guard5106 = cond_wire264_out;
wire _guard5107 = _guard5105 & _guard5106;
wire _guard5108 = fsm_out == 1'd0;
wire _guard5109 = _guard5107 & _guard5108;
wire _guard5110 = _guard5104 | _guard5109;
wire _guard5111 = early_reset_static_par0_go_out;
wire _guard5112 = _guard5110 & _guard5111;
wire _guard5113 = cond_wire_out;
wire _guard5114 = early_reset_static_par0_go_out;
wire _guard5115 = _guard5113 & _guard5114;
wire _guard5116 = cond_wire_out;
wire _guard5117 = early_reset_static_par0_go_out;
wire _guard5118 = _guard5116 & _guard5117;
wire _guard5119 = cond_wire_out;
wire _guard5120 = early_reset_static_par0_go_out;
wire _guard5121 = _guard5119 & _guard5120;
wire _guard5122 = cond_wire_out;
wire _guard5123 = early_reset_static_par0_go_out;
wire _guard5124 = _guard5122 & _guard5123;
wire _guard5125 = early_reset_static_par_go_out;
wire _guard5126 = early_reset_static_par0_go_out;
wire _guard5127 = _guard5125 | _guard5126;
wire _guard5128 = early_reset_static_par0_go_out;
wire _guard5129 = early_reset_static_par_go_out;
wire _guard5130 = early_reset_static_par0_go_out;
wire _guard5131 = early_reset_static_par0_go_out;
wire _guard5132 = early_reset_static_par0_go_out;
wire _guard5133 = early_reset_static_par0_go_out;
wire _guard5134 = early_reset_static_par0_go_out;
wire _guard5135 = early_reset_static_par0_go_out;
wire _guard5136 = early_reset_static_par0_go_out;
wire _guard5137 = early_reset_static_par0_go_out;
wire _guard5138 = early_reset_static_par0_go_out;
wire _guard5139 = early_reset_static_par0_go_out;
wire _guard5140 = ~_guard0;
wire _guard5141 = early_reset_static_par0_go_out;
wire _guard5142 = _guard5140 & _guard5141;
wire _guard5143 = early_reset_static_par0_go_out;
wire _guard5144 = ~_guard0;
wire _guard5145 = early_reset_static_par0_go_out;
wire _guard5146 = _guard5144 & _guard5145;
wire _guard5147 = early_reset_static_par0_go_out;
wire _guard5148 = early_reset_static_par0_go_out;
wire _guard5149 = early_reset_static_par0_go_out;
wire _guard5150 = ~_guard0;
wire _guard5151 = early_reset_static_par0_go_out;
wire _guard5152 = _guard5150 & _guard5151;
wire _guard5153 = early_reset_static_par0_go_out;
wire _guard5154 = early_reset_static_par0_go_out;
wire _guard5155 = early_reset_static_par0_go_out;
wire _guard5156 = early_reset_static_par0_go_out;
wire _guard5157 = early_reset_static_par0_go_out;
wire _guard5158 = early_reset_static_par0_go_out;
wire _guard5159 = early_reset_static_par0_go_out;
wire _guard5160 = early_reset_static_par0_go_out;
wire _guard5161 = early_reset_static_par0_go_out;
wire _guard5162 = ~_guard0;
wire _guard5163 = early_reset_static_par0_go_out;
wire _guard5164 = _guard5162 & _guard5163;
wire _guard5165 = early_reset_static_par0_go_out;
wire _guard5166 = ~_guard0;
wire _guard5167 = early_reset_static_par0_go_out;
wire _guard5168 = _guard5166 & _guard5167;
wire _guard5169 = early_reset_static_par0_go_out;
wire _guard5170 = early_reset_static_par0_go_out;
wire _guard5171 = early_reset_static_par0_go_out;
wire _guard5172 = ~_guard0;
wire _guard5173 = early_reset_static_par0_go_out;
wire _guard5174 = _guard5172 & _guard5173;
wire _guard5175 = early_reset_static_par0_go_out;
wire _guard5176 = ~_guard0;
wire _guard5177 = early_reset_static_par0_go_out;
wire _guard5178 = _guard5176 & _guard5177;
wire _guard5179 = early_reset_static_par0_go_out;
wire _guard5180 = early_reset_static_par0_go_out;
wire _guard5181 = early_reset_static_par0_go_out;
wire _guard5182 = early_reset_static_par0_go_out;
wire _guard5183 = early_reset_static_par0_go_out;
wire _guard5184 = early_reset_static_par0_go_out;
wire _guard5185 = ~_guard0;
wire _guard5186 = early_reset_static_par0_go_out;
wire _guard5187 = _guard5185 & _guard5186;
wire _guard5188 = early_reset_static_par0_go_out;
wire _guard5189 = early_reset_static_par0_go_out;
wire _guard5190 = early_reset_static_par0_go_out;
wire _guard5191 = early_reset_static_par0_go_out;
wire _guard5192 = ~_guard0;
wire _guard5193 = early_reset_static_par0_go_out;
wire _guard5194 = _guard5192 & _guard5193;
wire _guard5195 = early_reset_static_par0_go_out;
wire _guard5196 = early_reset_static_par0_go_out;
wire _guard5197 = early_reset_static_par0_go_out;
wire _guard5198 = early_reset_static_par0_go_out;
wire _guard5199 = early_reset_static_par0_go_out;
wire _guard5200 = ~_guard0;
wire _guard5201 = early_reset_static_par0_go_out;
wire _guard5202 = _guard5200 & _guard5201;
wire _guard5203 = early_reset_static_par0_go_out;
wire _guard5204 = early_reset_static_par0_go_out;
wire _guard5205 = ~_guard0;
wire _guard5206 = early_reset_static_par0_go_out;
wire _guard5207 = _guard5205 & _guard5206;
wire _guard5208 = early_reset_static_par0_go_out;
wire _guard5209 = ~_guard0;
wire _guard5210 = early_reset_static_par0_go_out;
wire _guard5211 = _guard5209 & _guard5210;
wire _guard5212 = early_reset_static_par0_go_out;
wire _guard5213 = early_reset_static_par0_go_out;
wire _guard5214 = early_reset_static_par0_go_out;
wire _guard5215 = ~_guard0;
wire _guard5216 = early_reset_static_par0_go_out;
wire _guard5217 = _guard5215 & _guard5216;
wire _guard5218 = early_reset_static_par0_go_out;
wire _guard5219 = ~_guard0;
wire _guard5220 = early_reset_static_par0_go_out;
wire _guard5221 = _guard5219 & _guard5220;
wire _guard5222 = early_reset_static_par0_go_out;
wire _guard5223 = early_reset_static_par0_go_out;
wire _guard5224 = early_reset_static_par0_go_out;
wire _guard5225 = ~_guard0;
wire _guard5226 = early_reset_static_par0_go_out;
wire _guard5227 = _guard5225 & _guard5226;
wire _guard5228 = early_reset_static_par0_go_out;
wire _guard5229 = early_reset_static_par0_go_out;
wire _guard5230 = ~_guard0;
wire _guard5231 = early_reset_static_par0_go_out;
wire _guard5232 = _guard5230 & _guard5231;
wire _guard5233 = early_reset_static_par0_go_out;
wire _guard5234 = early_reset_static_par0_go_out;
wire _guard5235 = early_reset_static_par0_go_out;
wire _guard5236 = early_reset_static_par0_go_out;
wire _guard5237 = ~_guard0;
wire _guard5238 = early_reset_static_par0_go_out;
wire _guard5239 = _guard5237 & _guard5238;
wire _guard5240 = early_reset_static_par0_go_out;
wire _guard5241 = ~_guard0;
wire _guard5242 = early_reset_static_par0_go_out;
wire _guard5243 = _guard5241 & _guard5242;
wire _guard5244 = early_reset_static_par0_go_out;
wire _guard5245 = early_reset_static_par0_go_out;
wire _guard5246 = ~_guard0;
wire _guard5247 = early_reset_static_par0_go_out;
wire _guard5248 = _guard5246 & _guard5247;
wire _guard5249 = early_reset_static_par0_go_out;
wire _guard5250 = early_reset_static_par0_go_out;
wire _guard5251 = ~_guard0;
wire _guard5252 = early_reset_static_par0_go_out;
wire _guard5253 = _guard5251 & _guard5252;
wire _guard5254 = early_reset_static_par0_go_out;
wire _guard5255 = ~_guard0;
wire _guard5256 = early_reset_static_par0_go_out;
wire _guard5257 = _guard5255 & _guard5256;
wire _guard5258 = early_reset_static_par0_go_out;
wire _guard5259 = early_reset_static_par0_go_out;
wire _guard5260 = fsm_out == 1'd0;
wire _guard5261 = signal_reg_out;
wire _guard5262 = _guard5260 & _guard5261;
wire _guard5263 = fsm_out == 1'd0;
wire _guard5264 = signal_reg_out;
wire _guard5265 = ~_guard5264;
wire _guard5266 = _guard5263 & _guard5265;
wire _guard5267 = wrapper_early_reset_static_par_go_out;
wire _guard5268 = _guard5266 & _guard5267;
wire _guard5269 = _guard5262 | _guard5268;
wire _guard5270 = fsm_out == 1'd0;
wire _guard5271 = signal_reg_out;
wire _guard5272 = ~_guard5271;
wire _guard5273 = _guard5270 & _guard5272;
wire _guard5274 = wrapper_early_reset_static_par_go_out;
wire _guard5275 = _guard5273 & _guard5274;
wire _guard5276 = fsm_out == 1'd0;
wire _guard5277 = signal_reg_out;
wire _guard5278 = _guard5276 & _guard5277;
wire _guard5279 = early_reset_static_par0_go_out;
wire _guard5280 = early_reset_static_par0_go_out;
wire _guard5281 = early_reset_static_par0_go_out;
wire _guard5282 = early_reset_static_par0_go_out;
wire _guard5283 = early_reset_static_par0_go_out;
wire _guard5284 = early_reset_static_par0_go_out;
wire _guard5285 = cond_wire19_out;
wire _guard5286 = early_reset_static_par0_go_out;
wire _guard5287 = _guard5285 & _guard5286;
wire _guard5288 = cond_wire19_out;
wire _guard5289 = early_reset_static_par0_go_out;
wire _guard5290 = _guard5288 & _guard5289;
wire _guard5291 = cond_wire21_out;
wire _guard5292 = early_reset_static_par0_go_out;
wire _guard5293 = _guard5291 & _guard5292;
wire _guard5294 = cond_wire21_out;
wire _guard5295 = early_reset_static_par0_go_out;
wire _guard5296 = _guard5294 & _guard5295;
wire _guard5297 = cond_wire75_out;
wire _guard5298 = early_reset_static_par0_go_out;
wire _guard5299 = _guard5297 & _guard5298;
wire _guard5300 = cond_wire73_out;
wire _guard5301 = early_reset_static_par0_go_out;
wire _guard5302 = _guard5300 & _guard5301;
wire _guard5303 = fsm_out == 1'd0;
wire _guard5304 = cond_wire73_out;
wire _guard5305 = _guard5303 & _guard5304;
wire _guard5306 = fsm_out == 1'd0;
wire _guard5307 = _guard5305 & _guard5306;
wire _guard5308 = fsm_out == 1'd0;
wire _guard5309 = cond_wire75_out;
wire _guard5310 = _guard5308 & _guard5309;
wire _guard5311 = fsm_out == 1'd0;
wire _guard5312 = _guard5310 & _guard5311;
wire _guard5313 = _guard5307 | _guard5312;
wire _guard5314 = early_reset_static_par0_go_out;
wire _guard5315 = _guard5313 & _guard5314;
wire _guard5316 = fsm_out == 1'd0;
wire _guard5317 = cond_wire73_out;
wire _guard5318 = _guard5316 & _guard5317;
wire _guard5319 = fsm_out == 1'd0;
wire _guard5320 = _guard5318 & _guard5319;
wire _guard5321 = fsm_out == 1'd0;
wire _guard5322 = cond_wire75_out;
wire _guard5323 = _guard5321 & _guard5322;
wire _guard5324 = fsm_out == 1'd0;
wire _guard5325 = _guard5323 & _guard5324;
wire _guard5326 = _guard5320 | _guard5325;
wire _guard5327 = early_reset_static_par0_go_out;
wire _guard5328 = _guard5326 & _guard5327;
wire _guard5329 = fsm_out == 1'd0;
wire _guard5330 = cond_wire73_out;
wire _guard5331 = _guard5329 & _guard5330;
wire _guard5332 = fsm_out == 1'd0;
wire _guard5333 = _guard5331 & _guard5332;
wire _guard5334 = fsm_out == 1'd0;
wire _guard5335 = cond_wire75_out;
wire _guard5336 = _guard5334 & _guard5335;
wire _guard5337 = fsm_out == 1'd0;
wire _guard5338 = _guard5336 & _guard5337;
wire _guard5339 = _guard5333 | _guard5338;
wire _guard5340 = early_reset_static_par0_go_out;
wire _guard5341 = _guard5339 & _guard5340;
wire _guard5342 = cond_wire74_out;
wire _guard5343 = early_reset_static_par0_go_out;
wire _guard5344 = _guard5342 & _guard5343;
wire _guard5345 = cond_wire74_out;
wire _guard5346 = early_reset_static_par0_go_out;
wire _guard5347 = _guard5345 & _guard5346;
wire _guard5348 = cond_wire49_out;
wire _guard5349 = early_reset_static_par0_go_out;
wire _guard5350 = _guard5348 & _guard5349;
wire _guard5351 = cond_wire49_out;
wire _guard5352 = early_reset_static_par0_go_out;
wire _guard5353 = _guard5351 & _guard5352;
wire _guard5354 = cond_wire90_out;
wire _guard5355 = early_reset_static_par0_go_out;
wire _guard5356 = _guard5354 & _guard5355;
wire _guard5357 = cond_wire90_out;
wire _guard5358 = early_reset_static_par0_go_out;
wire _guard5359 = _guard5357 & _guard5358;
wire _guard5360 = cond_wire127_out;
wire _guard5361 = early_reset_static_par0_go_out;
wire _guard5362 = _guard5360 & _guard5361;
wire _guard5363 = cond_wire127_out;
wire _guard5364 = early_reset_static_par0_go_out;
wire _guard5365 = _guard5363 & _guard5364;
wire _guard5366 = cond_wire157_out;
wire _guard5367 = early_reset_static_par0_go_out;
wire _guard5368 = _guard5366 & _guard5367;
wire _guard5369 = cond_wire155_out;
wire _guard5370 = early_reset_static_par0_go_out;
wire _guard5371 = _guard5369 & _guard5370;
wire _guard5372 = fsm_out == 1'd0;
wire _guard5373 = cond_wire155_out;
wire _guard5374 = _guard5372 & _guard5373;
wire _guard5375 = fsm_out == 1'd0;
wire _guard5376 = _guard5374 & _guard5375;
wire _guard5377 = fsm_out == 1'd0;
wire _guard5378 = cond_wire157_out;
wire _guard5379 = _guard5377 & _guard5378;
wire _guard5380 = fsm_out == 1'd0;
wire _guard5381 = _guard5379 & _guard5380;
wire _guard5382 = _guard5376 | _guard5381;
wire _guard5383 = early_reset_static_par0_go_out;
wire _guard5384 = _guard5382 & _guard5383;
wire _guard5385 = fsm_out == 1'd0;
wire _guard5386 = cond_wire155_out;
wire _guard5387 = _guard5385 & _guard5386;
wire _guard5388 = fsm_out == 1'd0;
wire _guard5389 = _guard5387 & _guard5388;
wire _guard5390 = fsm_out == 1'd0;
wire _guard5391 = cond_wire157_out;
wire _guard5392 = _guard5390 & _guard5391;
wire _guard5393 = fsm_out == 1'd0;
wire _guard5394 = _guard5392 & _guard5393;
wire _guard5395 = _guard5389 | _guard5394;
wire _guard5396 = early_reset_static_par0_go_out;
wire _guard5397 = _guard5395 & _guard5396;
wire _guard5398 = fsm_out == 1'd0;
wire _guard5399 = cond_wire155_out;
wire _guard5400 = _guard5398 & _guard5399;
wire _guard5401 = fsm_out == 1'd0;
wire _guard5402 = _guard5400 & _guard5401;
wire _guard5403 = fsm_out == 1'd0;
wire _guard5404 = cond_wire157_out;
wire _guard5405 = _guard5403 & _guard5404;
wire _guard5406 = fsm_out == 1'd0;
wire _guard5407 = _guard5405 & _guard5406;
wire _guard5408 = _guard5402 | _guard5407;
wire _guard5409 = early_reset_static_par0_go_out;
wire _guard5410 = _guard5408 & _guard5409;
wire _guard5411 = cond_wire152_out;
wire _guard5412 = early_reset_static_par0_go_out;
wire _guard5413 = _guard5411 & _guard5412;
wire _guard5414 = cond_wire152_out;
wire _guard5415 = early_reset_static_par0_go_out;
wire _guard5416 = _guard5414 & _guard5415;
wire _guard5417 = cond_wire169_out;
wire _guard5418 = early_reset_static_par0_go_out;
wire _guard5419 = _guard5417 & _guard5418;
wire _guard5420 = cond_wire167_out;
wire _guard5421 = early_reset_static_par0_go_out;
wire _guard5422 = _guard5420 & _guard5421;
wire _guard5423 = fsm_out == 1'd0;
wire _guard5424 = cond_wire167_out;
wire _guard5425 = _guard5423 & _guard5424;
wire _guard5426 = fsm_out == 1'd0;
wire _guard5427 = _guard5425 & _guard5426;
wire _guard5428 = fsm_out == 1'd0;
wire _guard5429 = cond_wire169_out;
wire _guard5430 = _guard5428 & _guard5429;
wire _guard5431 = fsm_out == 1'd0;
wire _guard5432 = _guard5430 & _guard5431;
wire _guard5433 = _guard5427 | _guard5432;
wire _guard5434 = early_reset_static_par0_go_out;
wire _guard5435 = _guard5433 & _guard5434;
wire _guard5436 = fsm_out == 1'd0;
wire _guard5437 = cond_wire167_out;
wire _guard5438 = _guard5436 & _guard5437;
wire _guard5439 = fsm_out == 1'd0;
wire _guard5440 = _guard5438 & _guard5439;
wire _guard5441 = fsm_out == 1'd0;
wire _guard5442 = cond_wire169_out;
wire _guard5443 = _guard5441 & _guard5442;
wire _guard5444 = fsm_out == 1'd0;
wire _guard5445 = _guard5443 & _guard5444;
wire _guard5446 = _guard5440 | _guard5445;
wire _guard5447 = early_reset_static_par0_go_out;
wire _guard5448 = _guard5446 & _guard5447;
wire _guard5449 = fsm_out == 1'd0;
wire _guard5450 = cond_wire167_out;
wire _guard5451 = _guard5449 & _guard5450;
wire _guard5452 = fsm_out == 1'd0;
wire _guard5453 = _guard5451 & _guard5452;
wire _guard5454 = fsm_out == 1'd0;
wire _guard5455 = cond_wire169_out;
wire _guard5456 = _guard5454 & _guard5455;
wire _guard5457 = fsm_out == 1'd0;
wire _guard5458 = _guard5456 & _guard5457;
wire _guard5459 = _guard5453 | _guard5458;
wire _guard5460 = early_reset_static_par0_go_out;
wire _guard5461 = _guard5459 & _guard5460;
wire _guard5462 = cond_wire189_out;
wire _guard5463 = early_reset_static_par0_go_out;
wire _guard5464 = _guard5462 & _guard5463;
wire _guard5465 = cond_wire189_out;
wire _guard5466 = early_reset_static_par0_go_out;
wire _guard5467 = _guard5465 & _guard5466;
wire _guard5468 = cond_wire237_out;
wire _guard5469 = early_reset_static_par0_go_out;
wire _guard5470 = _guard5468 & _guard5469;
wire _guard5471 = cond_wire237_out;
wire _guard5472 = early_reset_static_par0_go_out;
wire _guard5473 = _guard5471 & _guard5472;
wire _guard5474 = cond_wire218_out;
wire _guard5475 = early_reset_static_par0_go_out;
wire _guard5476 = _guard5474 & _guard5475;
wire _guard5477 = cond_wire218_out;
wire _guard5478 = early_reset_static_par0_go_out;
wire _guard5479 = _guard5477 & _guard5478;
wire _guard5480 = cond_wire230_out;
wire _guard5481 = early_reset_static_par0_go_out;
wire _guard5482 = _guard5480 & _guard5481;
wire _guard5483 = cond_wire230_out;
wire _guard5484 = early_reset_static_par0_go_out;
wire _guard5485 = _guard5483 & _guard5484;
wire _guard5486 = cond_wire4_out;
wire _guard5487 = early_reset_static_par0_go_out;
wire _guard5488 = _guard5486 & _guard5487;
wire _guard5489 = cond_wire4_out;
wire _guard5490 = early_reset_static_par0_go_out;
wire _guard5491 = _guard5489 & _guard5490;
wire _guard5492 = early_reset_static_par_go_out;
wire _guard5493 = cond_wire14_out;
wire _guard5494 = early_reset_static_par0_go_out;
wire _guard5495 = _guard5493 & _guard5494;
wire _guard5496 = _guard5492 | _guard5495;
wire _guard5497 = cond_wire14_out;
wire _guard5498 = early_reset_static_par0_go_out;
wire _guard5499 = _guard5497 & _guard5498;
wire _guard5500 = early_reset_static_par_go_out;
wire _guard5501 = cond_wire138_out;
wire _guard5502 = early_reset_static_par0_go_out;
wire _guard5503 = _guard5501 & _guard5502;
wire _guard5504 = cond_wire138_out;
wire _guard5505 = early_reset_static_par0_go_out;
wire _guard5506 = _guard5504 & _guard5505;
wire _guard5507 = early_reset_static_par0_go_out;
wire _guard5508 = early_reset_static_par0_go_out;
wire _guard5509 = early_reset_static_par0_go_out;
wire _guard5510 = early_reset_static_par0_go_out;
wire _guard5511 = early_reset_static_par0_go_out;
wire _guard5512 = early_reset_static_par0_go_out;
wire _guard5513 = early_reset_static_par0_go_out;
wire _guard5514 = early_reset_static_par0_go_out;
wire _guard5515 = early_reset_static_par0_go_out;
wire _guard5516 = early_reset_static_par0_go_out;
wire _guard5517 = early_reset_static_par0_go_out;
wire _guard5518 = early_reset_static_par0_go_out;
wire _guard5519 = early_reset_static_par0_go_out;
wire _guard5520 = early_reset_static_par0_go_out;
wire _guard5521 = early_reset_static_par0_go_out;
wire _guard5522 = early_reset_static_par0_go_out;
wire _guard5523 = early_reset_static_par_go_out;
wire _guard5524 = early_reset_static_par0_go_out;
wire _guard5525 = _guard5523 | _guard5524;
wire _guard5526 = early_reset_static_par_go_out;
wire _guard5527 = early_reset_static_par0_go_out;
wire _guard5528 = early_reset_static_par0_go_out;
wire _guard5529 = early_reset_static_par0_go_out;
wire _guard5530 = early_reset_static_par0_go_out;
wire _guard5531 = early_reset_static_par0_go_out;
wire _guard5532 = early_reset_static_par_go_out;
wire _guard5533 = early_reset_static_par0_go_out;
wire _guard5534 = _guard5532 | _guard5533;
wire _guard5535 = early_reset_static_par0_go_out;
wire _guard5536 = early_reset_static_par_go_out;
wire _guard5537 = early_reset_static_par_go_out;
wire _guard5538 = early_reset_static_par0_go_out;
wire _guard5539 = _guard5537 | _guard5538;
wire _guard5540 = early_reset_static_par_go_out;
wire _guard5541 = early_reset_static_par0_go_out;
wire _guard5542 = ~_guard0;
wire _guard5543 = early_reset_static_par0_go_out;
wire _guard5544 = _guard5542 & _guard5543;
wire _guard5545 = early_reset_static_par0_go_out;
wire _guard5546 = ~_guard0;
wire _guard5547 = early_reset_static_par0_go_out;
wire _guard5548 = _guard5546 & _guard5547;
wire _guard5549 = early_reset_static_par0_go_out;
wire _guard5550 = early_reset_static_par0_go_out;
wire _guard5551 = early_reset_static_par0_go_out;
wire _guard5552 = early_reset_static_par0_go_out;
wire _guard5553 = early_reset_static_par0_go_out;
wire _guard5554 = early_reset_static_par0_go_out;
wire _guard5555 = ~_guard0;
wire _guard5556 = early_reset_static_par0_go_out;
wire _guard5557 = _guard5555 & _guard5556;
wire _guard5558 = early_reset_static_par0_go_out;
wire _guard5559 = ~_guard0;
wire _guard5560 = early_reset_static_par0_go_out;
wire _guard5561 = _guard5559 & _guard5560;
wire _guard5562 = early_reset_static_par0_go_out;
wire _guard5563 = ~_guard0;
wire _guard5564 = early_reset_static_par0_go_out;
wire _guard5565 = _guard5563 & _guard5564;
wire _guard5566 = early_reset_static_par0_go_out;
wire _guard5567 = ~_guard0;
wire _guard5568 = early_reset_static_par0_go_out;
wire _guard5569 = _guard5567 & _guard5568;
wire _guard5570 = ~_guard0;
wire _guard5571 = early_reset_static_par0_go_out;
wire _guard5572 = _guard5570 & _guard5571;
wire _guard5573 = early_reset_static_par0_go_out;
wire _guard5574 = early_reset_static_par0_go_out;
wire _guard5575 = ~_guard0;
wire _guard5576 = early_reset_static_par0_go_out;
wire _guard5577 = _guard5575 & _guard5576;
wire _guard5578 = early_reset_static_par0_go_out;
wire _guard5579 = early_reset_static_par0_go_out;
wire _guard5580 = early_reset_static_par0_go_out;
wire _guard5581 = early_reset_static_par0_go_out;
wire _guard5582 = early_reset_static_par0_go_out;
wire _guard5583 = ~_guard0;
wire _guard5584 = early_reset_static_par0_go_out;
wire _guard5585 = _guard5583 & _guard5584;
wire _guard5586 = ~_guard0;
wire _guard5587 = early_reset_static_par0_go_out;
wire _guard5588 = _guard5586 & _guard5587;
wire _guard5589 = early_reset_static_par0_go_out;
wire _guard5590 = early_reset_static_par0_go_out;
wire _guard5591 = early_reset_static_par0_go_out;
wire _guard5592 = early_reset_static_par0_go_out;
wire _guard5593 = early_reset_static_par0_go_out;
wire _guard5594 = early_reset_static_par0_go_out;
wire _guard5595 = ~_guard0;
wire _guard5596 = early_reset_static_par0_go_out;
wire _guard5597 = _guard5595 & _guard5596;
wire _guard5598 = early_reset_static_par0_go_out;
wire _guard5599 = early_reset_static_par0_go_out;
wire _guard5600 = early_reset_static_par0_go_out;
wire _guard5601 = ~_guard0;
wire _guard5602 = early_reset_static_par0_go_out;
wire _guard5603 = _guard5601 & _guard5602;
wire _guard5604 = early_reset_static_par0_go_out;
wire _guard5605 = early_reset_static_par0_go_out;
wire _guard5606 = early_reset_static_par0_go_out;
wire _guard5607 = early_reset_static_par0_go_out;
wire _guard5608 = early_reset_static_par0_go_out;
wire _guard5609 = early_reset_static_par0_go_out;
wire _guard5610 = early_reset_static_par0_go_out;
wire _guard5611 = early_reset_static_par0_go_out;
wire _guard5612 = early_reset_static_par0_go_out;
wire _guard5613 = ~_guard0;
wire _guard5614 = early_reset_static_par0_go_out;
wire _guard5615 = _guard5613 & _guard5614;
wire _guard5616 = ~_guard0;
wire _guard5617 = early_reset_static_par0_go_out;
wire _guard5618 = _guard5616 & _guard5617;
wire _guard5619 = early_reset_static_par0_go_out;
wire _guard5620 = early_reset_static_par0_go_out;
wire _guard5621 = early_reset_static_par0_go_out;
wire _guard5622 = early_reset_static_par0_go_out;
wire _guard5623 = early_reset_static_par0_go_out;
wire _guard5624 = early_reset_static_par0_go_out;
wire _guard5625 = early_reset_static_par0_go_out;
wire _guard5626 = early_reset_static_par0_go_out;
wire _guard5627 = early_reset_static_par0_go_out;
wire _guard5628 = early_reset_static_par0_go_out;
wire _guard5629 = early_reset_static_par0_go_out;
wire _guard5630 = ~_guard0;
wire _guard5631 = early_reset_static_par0_go_out;
wire _guard5632 = _guard5630 & _guard5631;
wire _guard5633 = early_reset_static_par0_go_out;
wire _guard5634 = ~_guard0;
wire _guard5635 = early_reset_static_par0_go_out;
wire _guard5636 = _guard5634 & _guard5635;
wire _guard5637 = early_reset_static_par0_go_out;
wire _guard5638 = ~_guard0;
wire _guard5639 = early_reset_static_par0_go_out;
wire _guard5640 = _guard5638 & _guard5639;
wire _guard5641 = early_reset_static_par0_go_out;
wire _guard5642 = early_reset_static_par0_go_out;
wire _guard5643 = early_reset_static_par0_go_out;
wire _guard5644 = early_reset_static_par0_go_out;
wire _guard5645 = ~_guard0;
wire _guard5646 = early_reset_static_par0_go_out;
wire _guard5647 = _guard5645 & _guard5646;
wire _guard5648 = early_reset_static_par0_go_out;
wire _guard5649 = early_reset_static_par0_go_out;
wire _guard5650 = early_reset_static_par0_go_out;
wire _guard5651 = early_reset_static_par0_go_out;
wire _guard5652 = early_reset_static_par0_go_out;
wire _guard5653 = early_reset_static_par0_go_out;
wire _guard5654 = early_reset_static_par0_go_out;
wire _guard5655 = early_reset_static_par0_go_out;
wire _guard5656 = cond_wire2_out;
wire _guard5657 = early_reset_static_par0_go_out;
wire _guard5658 = _guard5656 & _guard5657;
wire _guard5659 = cond_wire0_out;
wire _guard5660 = early_reset_static_par0_go_out;
wire _guard5661 = _guard5659 & _guard5660;
wire _guard5662 = fsm_out == 1'd0;
wire _guard5663 = cond_wire0_out;
wire _guard5664 = _guard5662 & _guard5663;
wire _guard5665 = fsm_out == 1'd0;
wire _guard5666 = _guard5664 & _guard5665;
wire _guard5667 = fsm_out == 1'd0;
wire _guard5668 = cond_wire2_out;
wire _guard5669 = _guard5667 & _guard5668;
wire _guard5670 = fsm_out == 1'd0;
wire _guard5671 = _guard5669 & _guard5670;
wire _guard5672 = _guard5666 | _guard5671;
wire _guard5673 = early_reset_static_par0_go_out;
wire _guard5674 = _guard5672 & _guard5673;
wire _guard5675 = fsm_out == 1'd0;
wire _guard5676 = cond_wire0_out;
wire _guard5677 = _guard5675 & _guard5676;
wire _guard5678 = fsm_out == 1'd0;
wire _guard5679 = _guard5677 & _guard5678;
wire _guard5680 = fsm_out == 1'd0;
wire _guard5681 = cond_wire2_out;
wire _guard5682 = _guard5680 & _guard5681;
wire _guard5683 = fsm_out == 1'd0;
wire _guard5684 = _guard5682 & _guard5683;
wire _guard5685 = _guard5679 | _guard5684;
wire _guard5686 = early_reset_static_par0_go_out;
wire _guard5687 = _guard5685 & _guard5686;
wire _guard5688 = fsm_out == 1'd0;
wire _guard5689 = cond_wire0_out;
wire _guard5690 = _guard5688 & _guard5689;
wire _guard5691 = fsm_out == 1'd0;
wire _guard5692 = _guard5690 & _guard5691;
wire _guard5693 = fsm_out == 1'd0;
wire _guard5694 = cond_wire2_out;
wire _guard5695 = _guard5693 & _guard5694;
wire _guard5696 = fsm_out == 1'd0;
wire _guard5697 = _guard5695 & _guard5696;
wire _guard5698 = _guard5692 | _guard5697;
wire _guard5699 = early_reset_static_par0_go_out;
wire _guard5700 = _guard5698 & _guard5699;
wire _guard5701 = cond_wire61_out;
wire _guard5702 = early_reset_static_par0_go_out;
wire _guard5703 = _guard5701 & _guard5702;
wire _guard5704 = cond_wire61_out;
wire _guard5705 = early_reset_static_par0_go_out;
wire _guard5706 = _guard5704 & _guard5705;
wire _guard5707 = cond_wire120_out;
wire _guard5708 = early_reset_static_par0_go_out;
wire _guard5709 = _guard5707 & _guard5708;
wire _guard5710 = cond_wire118_out;
wire _guard5711 = early_reset_static_par0_go_out;
wire _guard5712 = _guard5710 & _guard5711;
wire _guard5713 = fsm_out == 1'd0;
wire _guard5714 = cond_wire118_out;
wire _guard5715 = _guard5713 & _guard5714;
wire _guard5716 = fsm_out == 1'd0;
wire _guard5717 = _guard5715 & _guard5716;
wire _guard5718 = fsm_out == 1'd0;
wire _guard5719 = cond_wire120_out;
wire _guard5720 = _guard5718 & _guard5719;
wire _guard5721 = fsm_out == 1'd0;
wire _guard5722 = _guard5720 & _guard5721;
wire _guard5723 = _guard5717 | _guard5722;
wire _guard5724 = early_reset_static_par0_go_out;
wire _guard5725 = _guard5723 & _guard5724;
wire _guard5726 = fsm_out == 1'd0;
wire _guard5727 = cond_wire118_out;
wire _guard5728 = _guard5726 & _guard5727;
wire _guard5729 = fsm_out == 1'd0;
wire _guard5730 = _guard5728 & _guard5729;
wire _guard5731 = fsm_out == 1'd0;
wire _guard5732 = cond_wire120_out;
wire _guard5733 = _guard5731 & _guard5732;
wire _guard5734 = fsm_out == 1'd0;
wire _guard5735 = _guard5733 & _guard5734;
wire _guard5736 = _guard5730 | _guard5735;
wire _guard5737 = early_reset_static_par0_go_out;
wire _guard5738 = _guard5736 & _guard5737;
wire _guard5739 = fsm_out == 1'd0;
wire _guard5740 = cond_wire118_out;
wire _guard5741 = _guard5739 & _guard5740;
wire _guard5742 = fsm_out == 1'd0;
wire _guard5743 = _guard5741 & _guard5742;
wire _guard5744 = fsm_out == 1'd0;
wire _guard5745 = cond_wire120_out;
wire _guard5746 = _guard5744 & _guard5745;
wire _guard5747 = fsm_out == 1'd0;
wire _guard5748 = _guard5746 & _guard5747;
wire _guard5749 = _guard5743 | _guard5748;
wire _guard5750 = early_reset_static_par0_go_out;
wire _guard5751 = _guard5749 & _guard5750;
wire _guard5752 = cond_wire86_out;
wire _guard5753 = early_reset_static_par0_go_out;
wire _guard5754 = _guard5752 & _guard5753;
wire _guard5755 = cond_wire86_out;
wire _guard5756 = early_reset_static_par0_go_out;
wire _guard5757 = _guard5755 & _guard5756;
wire _guard5758 = cond_wire119_out;
wire _guard5759 = early_reset_static_par0_go_out;
wire _guard5760 = _guard5758 & _guard5759;
wire _guard5761 = cond_wire119_out;
wire _guard5762 = early_reset_static_par0_go_out;
wire _guard5763 = _guard5761 & _guard5762;
wire _guard5764 = cond_wire131_out;
wire _guard5765 = early_reset_static_par0_go_out;
wire _guard5766 = _guard5764 & _guard5765;
wire _guard5767 = cond_wire131_out;
wire _guard5768 = early_reset_static_par0_go_out;
wire _guard5769 = _guard5767 & _guard5768;
wire _guard5770 = cond_wire198_out;
wire _guard5771 = early_reset_static_par0_go_out;
wire _guard5772 = _guard5770 & _guard5771;
wire _guard5773 = cond_wire196_out;
wire _guard5774 = early_reset_static_par0_go_out;
wire _guard5775 = _guard5773 & _guard5774;
wire _guard5776 = fsm_out == 1'd0;
wire _guard5777 = cond_wire196_out;
wire _guard5778 = _guard5776 & _guard5777;
wire _guard5779 = fsm_out == 1'd0;
wire _guard5780 = _guard5778 & _guard5779;
wire _guard5781 = fsm_out == 1'd0;
wire _guard5782 = cond_wire198_out;
wire _guard5783 = _guard5781 & _guard5782;
wire _guard5784 = fsm_out == 1'd0;
wire _guard5785 = _guard5783 & _guard5784;
wire _guard5786 = _guard5780 | _guard5785;
wire _guard5787 = early_reset_static_par0_go_out;
wire _guard5788 = _guard5786 & _guard5787;
wire _guard5789 = fsm_out == 1'd0;
wire _guard5790 = cond_wire196_out;
wire _guard5791 = _guard5789 & _guard5790;
wire _guard5792 = fsm_out == 1'd0;
wire _guard5793 = _guard5791 & _guard5792;
wire _guard5794 = fsm_out == 1'd0;
wire _guard5795 = cond_wire198_out;
wire _guard5796 = _guard5794 & _guard5795;
wire _guard5797 = fsm_out == 1'd0;
wire _guard5798 = _guard5796 & _guard5797;
wire _guard5799 = _guard5793 | _guard5798;
wire _guard5800 = early_reset_static_par0_go_out;
wire _guard5801 = _guard5799 & _guard5800;
wire _guard5802 = fsm_out == 1'd0;
wire _guard5803 = cond_wire196_out;
wire _guard5804 = _guard5802 & _guard5803;
wire _guard5805 = fsm_out == 1'd0;
wire _guard5806 = _guard5804 & _guard5805;
wire _guard5807 = fsm_out == 1'd0;
wire _guard5808 = cond_wire198_out;
wire _guard5809 = _guard5807 & _guard5808;
wire _guard5810 = fsm_out == 1'd0;
wire _guard5811 = _guard5809 & _guard5810;
wire _guard5812 = _guard5806 | _guard5811;
wire _guard5813 = early_reset_static_par0_go_out;
wire _guard5814 = _guard5812 & _guard5813;
wire _guard5815 = cond_wire164_out;
wire _guard5816 = early_reset_static_par0_go_out;
wire _guard5817 = _guard5815 & _guard5816;
wire _guard5818 = cond_wire164_out;
wire _guard5819 = early_reset_static_par0_go_out;
wire _guard5820 = _guard5818 & _guard5819;
wire _guard5821 = cond_wire181_out;
wire _guard5822 = early_reset_static_par0_go_out;
wire _guard5823 = _guard5821 & _guard5822;
wire _guard5824 = cond_wire181_out;
wire _guard5825 = early_reset_static_par0_go_out;
wire _guard5826 = _guard5824 & _guard5825;
wire _guard5827 = cond_wire244_out;
wire _guard5828 = early_reset_static_par0_go_out;
wire _guard5829 = _guard5827 & _guard5828;
wire _guard5830 = cond_wire242_out;
wire _guard5831 = early_reset_static_par0_go_out;
wire _guard5832 = _guard5830 & _guard5831;
wire _guard5833 = fsm_out == 1'd0;
wire _guard5834 = cond_wire242_out;
wire _guard5835 = _guard5833 & _guard5834;
wire _guard5836 = fsm_out == 1'd0;
wire _guard5837 = _guard5835 & _guard5836;
wire _guard5838 = fsm_out == 1'd0;
wire _guard5839 = cond_wire244_out;
wire _guard5840 = _guard5838 & _guard5839;
wire _guard5841 = fsm_out == 1'd0;
wire _guard5842 = _guard5840 & _guard5841;
wire _guard5843 = _guard5837 | _guard5842;
wire _guard5844 = early_reset_static_par0_go_out;
wire _guard5845 = _guard5843 & _guard5844;
wire _guard5846 = fsm_out == 1'd0;
wire _guard5847 = cond_wire242_out;
wire _guard5848 = _guard5846 & _guard5847;
wire _guard5849 = fsm_out == 1'd0;
wire _guard5850 = _guard5848 & _guard5849;
wire _guard5851 = fsm_out == 1'd0;
wire _guard5852 = cond_wire244_out;
wire _guard5853 = _guard5851 & _guard5852;
wire _guard5854 = fsm_out == 1'd0;
wire _guard5855 = _guard5853 & _guard5854;
wire _guard5856 = _guard5850 | _guard5855;
wire _guard5857 = early_reset_static_par0_go_out;
wire _guard5858 = _guard5856 & _guard5857;
wire _guard5859 = fsm_out == 1'd0;
wire _guard5860 = cond_wire242_out;
wire _guard5861 = _guard5859 & _guard5860;
wire _guard5862 = fsm_out == 1'd0;
wire _guard5863 = _guard5861 & _guard5862;
wire _guard5864 = fsm_out == 1'd0;
wire _guard5865 = cond_wire244_out;
wire _guard5866 = _guard5864 & _guard5865;
wire _guard5867 = fsm_out == 1'd0;
wire _guard5868 = _guard5866 & _guard5867;
wire _guard5869 = _guard5863 | _guard5868;
wire _guard5870 = early_reset_static_par0_go_out;
wire _guard5871 = _guard5869 & _guard5870;
wire _guard5872 = cond_wire9_out;
wire _guard5873 = early_reset_static_par0_go_out;
wire _guard5874 = _guard5872 & _guard5873;
wire _guard5875 = cond_wire9_out;
wire _guard5876 = early_reset_static_par0_go_out;
wire _guard5877 = _guard5875 & _guard5876;
wire _guard5878 = cond_wire24_out;
wire _guard5879 = early_reset_static_par0_go_out;
wire _guard5880 = _guard5878 & _guard5879;
wire _guard5881 = cond_wire24_out;
wire _guard5882 = early_reset_static_par0_go_out;
wire _guard5883 = _guard5881 & _guard5882;
wire _guard5884 = early_reset_static_par0_go_out;
wire _guard5885 = early_reset_static_par0_go_out;
wire _guard5886 = early_reset_static_par_go_out;
wire _guard5887 = early_reset_static_par0_go_out;
wire _guard5888 = _guard5886 | _guard5887;
wire _guard5889 = early_reset_static_par0_go_out;
wire _guard5890 = early_reset_static_par_go_out;
wire _guard5891 = early_reset_static_par_go_out;
wire _guard5892 = early_reset_static_par0_go_out;
wire _guard5893 = _guard5891 | _guard5892;
wire _guard5894 = early_reset_static_par_go_out;
wire _guard5895 = early_reset_static_par0_go_out;
wire _guard5896 = early_reset_static_par0_go_out;
wire _guard5897 = early_reset_static_par0_go_out;
wire _guard5898 = early_reset_static_par_go_out;
wire _guard5899 = early_reset_static_par0_go_out;
wire _guard5900 = _guard5898 | _guard5899;
wire _guard5901 = early_reset_static_par0_go_out;
wire _guard5902 = early_reset_static_par_go_out;
wire _guard5903 = early_reset_static_par_go_out;
wire _guard5904 = early_reset_static_par0_go_out;
wire _guard5905 = _guard5903 | _guard5904;
wire _guard5906 = early_reset_static_par_go_out;
wire _guard5907 = early_reset_static_par0_go_out;
wire _guard5908 = early_reset_static_par0_go_out;
wire _guard5909 = early_reset_static_par0_go_out;
wire _guard5910 = early_reset_static_par_go_out;
wire _guard5911 = early_reset_static_par0_go_out;
wire _guard5912 = _guard5910 | _guard5911;
wire _guard5913 = early_reset_static_par0_go_out;
wire _guard5914 = early_reset_static_par_go_out;
wire _guard5915 = early_reset_static_par0_go_out;
wire _guard5916 = early_reset_static_par0_go_out;
wire _guard5917 = early_reset_static_par_go_out;
wire _guard5918 = early_reset_static_par0_go_out;
wire _guard5919 = _guard5917 | _guard5918;
wire _guard5920 = early_reset_static_par_go_out;
wire _guard5921 = early_reset_static_par0_go_out;
wire _guard5922 = early_reset_static_par0_go_out;
wire _guard5923 = early_reset_static_par0_go_out;
wire _guard5924 = early_reset_static_par0_go_out;
wire _guard5925 = early_reset_static_par0_go_out;
wire _guard5926 = early_reset_static_par0_go_out;
wire _guard5927 = early_reset_static_par0_go_out;
wire _guard5928 = early_reset_static_par0_go_out;
wire _guard5929 = early_reset_static_par0_go_out;
wire _guard5930 = early_reset_static_par_go_out;
wire _guard5931 = early_reset_static_par0_go_out;
wire _guard5932 = _guard5930 | _guard5931;
wire _guard5933 = early_reset_static_par0_go_out;
wire _guard5934 = early_reset_static_par_go_out;
wire _guard5935 = early_reset_static_par0_go_out;
wire _guard5936 = early_reset_static_par0_go_out;
wire _guard5937 = early_reset_static_par0_go_out;
wire _guard5938 = early_reset_static_par0_go_out;
wire _guard5939 = early_reset_static_par_go_out;
wire _guard5940 = early_reset_static_par0_go_out;
wire _guard5941 = _guard5939 | _guard5940;
wire _guard5942 = early_reset_static_par0_go_out;
wire _guard5943 = early_reset_static_par_go_out;
wire _guard5944 = early_reset_static_par_go_out;
wire _guard5945 = early_reset_static_par0_go_out;
wire _guard5946 = _guard5944 | _guard5945;
wire _guard5947 = early_reset_static_par_go_out;
wire _guard5948 = early_reset_static_par0_go_out;
wire _guard5949 = early_reset_static_par0_go_out;
wire _guard5950 = early_reset_static_par0_go_out;
wire _guard5951 = early_reset_static_par0_go_out;
wire _guard5952 = early_reset_static_par0_go_out;
wire _guard5953 = early_reset_static_par0_go_out;
wire _guard5954 = early_reset_static_par0_go_out;
wire _guard5955 = early_reset_static_par0_go_out;
wire _guard5956 = early_reset_static_par0_go_out;
wire _guard5957 = ~_guard0;
wire _guard5958 = early_reset_static_par0_go_out;
wire _guard5959 = _guard5957 & _guard5958;
wire _guard5960 = early_reset_static_par0_go_out;
wire _guard5961 = early_reset_static_par0_go_out;
wire _guard5962 = ~_guard0;
wire _guard5963 = early_reset_static_par0_go_out;
wire _guard5964 = _guard5962 & _guard5963;
wire _guard5965 = early_reset_static_par0_go_out;
wire _guard5966 = ~_guard0;
wire _guard5967 = early_reset_static_par0_go_out;
wire _guard5968 = _guard5966 & _guard5967;
wire _guard5969 = ~_guard0;
wire _guard5970 = early_reset_static_par0_go_out;
wire _guard5971 = _guard5969 & _guard5970;
wire _guard5972 = early_reset_static_par0_go_out;
wire _guard5973 = ~_guard0;
wire _guard5974 = early_reset_static_par0_go_out;
wire _guard5975 = _guard5973 & _guard5974;
wire _guard5976 = early_reset_static_par0_go_out;
wire _guard5977 = early_reset_static_par0_go_out;
wire _guard5978 = ~_guard0;
wire _guard5979 = early_reset_static_par0_go_out;
wire _guard5980 = _guard5978 & _guard5979;
wire _guard5981 = early_reset_static_par0_go_out;
wire _guard5982 = ~_guard0;
wire _guard5983 = early_reset_static_par0_go_out;
wire _guard5984 = _guard5982 & _guard5983;
wire _guard5985 = early_reset_static_par0_go_out;
wire _guard5986 = early_reset_static_par0_go_out;
wire _guard5987 = early_reset_static_par0_go_out;
wire _guard5988 = ~_guard0;
wire _guard5989 = early_reset_static_par0_go_out;
wire _guard5990 = _guard5988 & _guard5989;
wire _guard5991 = early_reset_static_par0_go_out;
wire _guard5992 = early_reset_static_par0_go_out;
wire _guard5993 = early_reset_static_par0_go_out;
wire _guard5994 = early_reset_static_par0_go_out;
wire _guard5995 = early_reset_static_par0_go_out;
wire _guard5996 = early_reset_static_par0_go_out;
wire _guard5997 = ~_guard0;
wire _guard5998 = early_reset_static_par0_go_out;
wire _guard5999 = _guard5997 & _guard5998;
wire _guard6000 = early_reset_static_par0_go_out;
wire _guard6001 = ~_guard0;
wire _guard6002 = early_reset_static_par0_go_out;
wire _guard6003 = _guard6001 & _guard6002;
wire _guard6004 = early_reset_static_par0_go_out;
wire _guard6005 = early_reset_static_par0_go_out;
wire _guard6006 = early_reset_static_par0_go_out;
wire _guard6007 = early_reset_static_par0_go_out;
wire _guard6008 = early_reset_static_par0_go_out;
wire _guard6009 = ~_guard0;
wire _guard6010 = early_reset_static_par0_go_out;
wire _guard6011 = _guard6009 & _guard6010;
wire _guard6012 = early_reset_static_par0_go_out;
wire _guard6013 = early_reset_static_par0_go_out;
wire _guard6014 = early_reset_static_par0_go_out;
wire _guard6015 = early_reset_static_par0_go_out;
wire _guard6016 = ~_guard0;
wire _guard6017 = early_reset_static_par0_go_out;
wire _guard6018 = _guard6016 & _guard6017;
wire _guard6019 = early_reset_static_par0_go_out;
wire _guard6020 = early_reset_static_par0_go_out;
wire _guard6021 = early_reset_static_par0_go_out;
wire _guard6022 = ~_guard0;
wire _guard6023 = early_reset_static_par0_go_out;
wire _guard6024 = _guard6022 & _guard6023;
wire _guard6025 = early_reset_static_par0_go_out;
wire _guard6026 = early_reset_static_par0_go_out;
wire _guard6027 = early_reset_static_par0_go_out;
wire _guard6028 = early_reset_static_par0_go_out;
wire _guard6029 = early_reset_static_par0_go_out;
wire _guard6030 = ~_guard0;
wire _guard6031 = early_reset_static_par0_go_out;
wire _guard6032 = _guard6030 & _guard6031;
wire _guard6033 = early_reset_static_par0_go_out;
wire _guard6034 = ~_guard0;
wire _guard6035 = early_reset_static_par0_go_out;
wire _guard6036 = _guard6034 & _guard6035;
wire _guard6037 = early_reset_static_par0_go_out;
wire _guard6038 = early_reset_static_par0_go_out;
wire _guard6039 = ~_guard0;
wire _guard6040 = early_reset_static_par0_go_out;
wire _guard6041 = _guard6039 & _guard6040;
wire _guard6042 = early_reset_static_par0_go_out;
wire _guard6043 = ~_guard0;
wire _guard6044 = early_reset_static_par0_go_out;
wire _guard6045 = _guard6043 & _guard6044;
wire _guard6046 = early_reset_static_par0_go_out;
wire _guard6047 = early_reset_static_par0_go_out;
wire _guard6048 = ~_guard0;
wire _guard6049 = early_reset_static_par0_go_out;
wire _guard6050 = _guard6048 & _guard6049;
wire _guard6051 = early_reset_static_par0_go_out;
wire _guard6052 = early_reset_static_par0_go_out;
wire _guard6053 = early_reset_static_par0_go_out;
wire _guard6054 = early_reset_static_par0_go_out;
wire _guard6055 = early_reset_static_par0_go_out;
wire _guard6056 = early_reset_static_par0_go_out;
wire _guard6057 = ~_guard0;
wire _guard6058 = early_reset_static_par0_go_out;
wire _guard6059 = _guard6057 & _guard6058;
wire _guard6060 = early_reset_static_par0_go_out;
wire _guard6061 = early_reset_static_par0_go_out;
wire _guard6062 = ~_guard0;
wire _guard6063 = early_reset_static_par0_go_out;
wire _guard6064 = _guard6062 & _guard6063;
wire _guard6065 = fsm0_out == 2'd2;
wire _guard6066 = cond_wire14_out;
wire _guard6067 = early_reset_static_par0_go_out;
wire _guard6068 = _guard6066 & _guard6067;
wire _guard6069 = cond_wire14_out;
wire _guard6070 = early_reset_static_par0_go_out;
wire _guard6071 = _guard6069 & _guard6070;
wire _guard6072 = cond_wire32_out;
wire _guard6073 = early_reset_static_par0_go_out;
wire _guard6074 = _guard6072 & _guard6073;
wire _guard6075 = cond_wire30_out;
wire _guard6076 = early_reset_static_par0_go_out;
wire _guard6077 = _guard6075 & _guard6076;
wire _guard6078 = fsm_out == 1'd0;
wire _guard6079 = cond_wire30_out;
wire _guard6080 = _guard6078 & _guard6079;
wire _guard6081 = fsm_out == 1'd0;
wire _guard6082 = _guard6080 & _guard6081;
wire _guard6083 = fsm_out == 1'd0;
wire _guard6084 = cond_wire32_out;
wire _guard6085 = _guard6083 & _guard6084;
wire _guard6086 = fsm_out == 1'd0;
wire _guard6087 = _guard6085 & _guard6086;
wire _guard6088 = _guard6082 | _guard6087;
wire _guard6089 = early_reset_static_par0_go_out;
wire _guard6090 = _guard6088 & _guard6089;
wire _guard6091 = fsm_out == 1'd0;
wire _guard6092 = cond_wire30_out;
wire _guard6093 = _guard6091 & _guard6092;
wire _guard6094 = fsm_out == 1'd0;
wire _guard6095 = _guard6093 & _guard6094;
wire _guard6096 = fsm_out == 1'd0;
wire _guard6097 = cond_wire32_out;
wire _guard6098 = _guard6096 & _guard6097;
wire _guard6099 = fsm_out == 1'd0;
wire _guard6100 = _guard6098 & _guard6099;
wire _guard6101 = _guard6095 | _guard6100;
wire _guard6102 = early_reset_static_par0_go_out;
wire _guard6103 = _guard6101 & _guard6102;
wire _guard6104 = fsm_out == 1'd0;
wire _guard6105 = cond_wire30_out;
wire _guard6106 = _guard6104 & _guard6105;
wire _guard6107 = fsm_out == 1'd0;
wire _guard6108 = _guard6106 & _guard6107;
wire _guard6109 = fsm_out == 1'd0;
wire _guard6110 = cond_wire32_out;
wire _guard6111 = _guard6109 & _guard6110;
wire _guard6112 = fsm_out == 1'd0;
wire _guard6113 = _guard6111 & _guard6112;
wire _guard6114 = _guard6108 | _guard6113;
wire _guard6115 = early_reset_static_par0_go_out;
wire _guard6116 = _guard6114 & _guard6115;
wire _guard6117 = cond_wire36_out;
wire _guard6118 = early_reset_static_par0_go_out;
wire _guard6119 = _guard6117 & _guard6118;
wire _guard6120 = cond_wire36_out;
wire _guard6121 = early_reset_static_par0_go_out;
wire _guard6122 = _guard6120 & _guard6121;
wire _guard6123 = cond_wire45_out;
wire _guard6124 = early_reset_static_par0_go_out;
wire _guard6125 = _guard6123 & _guard6124;
wire _guard6126 = cond_wire45_out;
wire _guard6127 = early_reset_static_par0_go_out;
wire _guard6128 = _guard6126 & _guard6127;
wire _guard6129 = cond_wire115_out;
wire _guard6130 = early_reset_static_par0_go_out;
wire _guard6131 = _guard6129 & _guard6130;
wire _guard6132 = cond_wire115_out;
wire _guard6133 = early_reset_static_par0_go_out;
wire _guard6134 = _guard6132 & _guard6133;
wire _guard6135 = cond_wire102_out;
wire _guard6136 = early_reset_static_par0_go_out;
wire _guard6137 = _guard6135 & _guard6136;
wire _guard6138 = cond_wire102_out;
wire _guard6139 = early_reset_static_par0_go_out;
wire _guard6140 = _guard6138 & _guard6139;
wire _guard6141 = cond_wire140_out;
wire _guard6142 = early_reset_static_par0_go_out;
wire _guard6143 = _guard6141 & _guard6142;
wire _guard6144 = cond_wire140_out;
wire _guard6145 = early_reset_static_par0_go_out;
wire _guard6146 = _guard6144 & _guard6145;
wire _guard6147 = cond_wire153_out;
wire _guard6148 = early_reset_static_par0_go_out;
wire _guard6149 = _guard6147 & _guard6148;
wire _guard6150 = cond_wire151_out;
wire _guard6151 = early_reset_static_par0_go_out;
wire _guard6152 = _guard6150 & _guard6151;
wire _guard6153 = fsm_out == 1'd0;
wire _guard6154 = cond_wire151_out;
wire _guard6155 = _guard6153 & _guard6154;
wire _guard6156 = fsm_out == 1'd0;
wire _guard6157 = _guard6155 & _guard6156;
wire _guard6158 = fsm_out == 1'd0;
wire _guard6159 = cond_wire153_out;
wire _guard6160 = _guard6158 & _guard6159;
wire _guard6161 = fsm_out == 1'd0;
wire _guard6162 = _guard6160 & _guard6161;
wire _guard6163 = _guard6157 | _guard6162;
wire _guard6164 = early_reset_static_par0_go_out;
wire _guard6165 = _guard6163 & _guard6164;
wire _guard6166 = fsm_out == 1'd0;
wire _guard6167 = cond_wire151_out;
wire _guard6168 = _guard6166 & _guard6167;
wire _guard6169 = fsm_out == 1'd0;
wire _guard6170 = _guard6168 & _guard6169;
wire _guard6171 = fsm_out == 1'd0;
wire _guard6172 = cond_wire153_out;
wire _guard6173 = _guard6171 & _guard6172;
wire _guard6174 = fsm_out == 1'd0;
wire _guard6175 = _guard6173 & _guard6174;
wire _guard6176 = _guard6170 | _guard6175;
wire _guard6177 = early_reset_static_par0_go_out;
wire _guard6178 = _guard6176 & _guard6177;
wire _guard6179 = fsm_out == 1'd0;
wire _guard6180 = cond_wire151_out;
wire _guard6181 = _guard6179 & _guard6180;
wire _guard6182 = fsm_out == 1'd0;
wire _guard6183 = _guard6181 & _guard6182;
wire _guard6184 = fsm_out == 1'd0;
wire _guard6185 = cond_wire153_out;
wire _guard6186 = _guard6184 & _guard6185;
wire _guard6187 = fsm_out == 1'd0;
wire _guard6188 = _guard6186 & _guard6187;
wire _guard6189 = _guard6183 | _guard6188;
wire _guard6190 = early_reset_static_par0_go_out;
wire _guard6191 = _guard6189 & _guard6190;
wire _guard6192 = cond_wire171_out;
wire _guard6193 = early_reset_static_par0_go_out;
wire _guard6194 = _guard6192 & _guard6193;
wire _guard6195 = cond_wire171_out;
wire _guard6196 = early_reset_static_par0_go_out;
wire _guard6197 = _guard6195 & _guard6196;
wire _guard6198 = cond_wire231_out;
wire _guard6199 = early_reset_static_par0_go_out;
wire _guard6200 = _guard6198 & _guard6199;
wire _guard6201 = cond_wire229_out;
wire _guard6202 = early_reset_static_par0_go_out;
wire _guard6203 = _guard6201 & _guard6202;
wire _guard6204 = fsm_out == 1'd0;
wire _guard6205 = cond_wire229_out;
wire _guard6206 = _guard6204 & _guard6205;
wire _guard6207 = fsm_out == 1'd0;
wire _guard6208 = _guard6206 & _guard6207;
wire _guard6209 = fsm_out == 1'd0;
wire _guard6210 = cond_wire231_out;
wire _guard6211 = _guard6209 & _guard6210;
wire _guard6212 = fsm_out == 1'd0;
wire _guard6213 = _guard6211 & _guard6212;
wire _guard6214 = _guard6208 | _guard6213;
wire _guard6215 = early_reset_static_par0_go_out;
wire _guard6216 = _guard6214 & _guard6215;
wire _guard6217 = fsm_out == 1'd0;
wire _guard6218 = cond_wire229_out;
wire _guard6219 = _guard6217 & _guard6218;
wire _guard6220 = fsm_out == 1'd0;
wire _guard6221 = _guard6219 & _guard6220;
wire _guard6222 = fsm_out == 1'd0;
wire _guard6223 = cond_wire231_out;
wire _guard6224 = _guard6222 & _guard6223;
wire _guard6225 = fsm_out == 1'd0;
wire _guard6226 = _guard6224 & _guard6225;
wire _guard6227 = _guard6221 | _guard6226;
wire _guard6228 = early_reset_static_par0_go_out;
wire _guard6229 = _guard6227 & _guard6228;
wire _guard6230 = fsm_out == 1'd0;
wire _guard6231 = cond_wire229_out;
wire _guard6232 = _guard6230 & _guard6231;
wire _guard6233 = fsm_out == 1'd0;
wire _guard6234 = _guard6232 & _guard6233;
wire _guard6235 = fsm_out == 1'd0;
wire _guard6236 = cond_wire231_out;
wire _guard6237 = _guard6235 & _guard6236;
wire _guard6238 = fsm_out == 1'd0;
wire _guard6239 = _guard6237 & _guard6238;
wire _guard6240 = _guard6234 | _guard6239;
wire _guard6241 = early_reset_static_par0_go_out;
wire _guard6242 = _guard6240 & _guard6241;
wire _guard6243 = cond_wire248_out;
wire _guard6244 = early_reset_static_par0_go_out;
wire _guard6245 = _guard6243 & _guard6244;
wire _guard6246 = cond_wire246_out;
wire _guard6247 = early_reset_static_par0_go_out;
wire _guard6248 = _guard6246 & _guard6247;
wire _guard6249 = fsm_out == 1'd0;
wire _guard6250 = cond_wire246_out;
wire _guard6251 = _guard6249 & _guard6250;
wire _guard6252 = fsm_out == 1'd0;
wire _guard6253 = _guard6251 & _guard6252;
wire _guard6254 = fsm_out == 1'd0;
wire _guard6255 = cond_wire248_out;
wire _guard6256 = _guard6254 & _guard6255;
wire _guard6257 = fsm_out == 1'd0;
wire _guard6258 = _guard6256 & _guard6257;
wire _guard6259 = _guard6253 | _guard6258;
wire _guard6260 = early_reset_static_par0_go_out;
wire _guard6261 = _guard6259 & _guard6260;
wire _guard6262 = fsm_out == 1'd0;
wire _guard6263 = cond_wire246_out;
wire _guard6264 = _guard6262 & _guard6263;
wire _guard6265 = fsm_out == 1'd0;
wire _guard6266 = _guard6264 & _guard6265;
wire _guard6267 = fsm_out == 1'd0;
wire _guard6268 = cond_wire248_out;
wire _guard6269 = _guard6267 & _guard6268;
wire _guard6270 = fsm_out == 1'd0;
wire _guard6271 = _guard6269 & _guard6270;
wire _guard6272 = _guard6266 | _guard6271;
wire _guard6273 = early_reset_static_par0_go_out;
wire _guard6274 = _guard6272 & _guard6273;
wire _guard6275 = fsm_out == 1'd0;
wire _guard6276 = cond_wire246_out;
wire _guard6277 = _guard6275 & _guard6276;
wire _guard6278 = fsm_out == 1'd0;
wire _guard6279 = _guard6277 & _guard6278;
wire _guard6280 = fsm_out == 1'd0;
wire _guard6281 = cond_wire248_out;
wire _guard6282 = _guard6280 & _guard6281;
wire _guard6283 = fsm_out == 1'd0;
wire _guard6284 = _guard6282 & _guard6283;
wire _guard6285 = _guard6279 | _guard6284;
wire _guard6286 = early_reset_static_par0_go_out;
wire _guard6287 = _guard6285 & _guard6286;
wire _guard6288 = cond_wire267_out;
wire _guard6289 = early_reset_static_par0_go_out;
wire _guard6290 = _guard6288 & _guard6289;
wire _guard6291 = cond_wire266_out;
wire _guard6292 = early_reset_static_par0_go_out;
wire _guard6293 = _guard6291 & _guard6292;
wire _guard6294 = fsm_out == 1'd0;
wire _guard6295 = cond_wire266_out;
wire _guard6296 = _guard6294 & _guard6295;
wire _guard6297 = fsm_out == 1'd0;
wire _guard6298 = _guard6296 & _guard6297;
wire _guard6299 = fsm_out == 1'd0;
wire _guard6300 = cond_wire267_out;
wire _guard6301 = _guard6299 & _guard6300;
wire _guard6302 = fsm_out == 1'd0;
wire _guard6303 = _guard6301 & _guard6302;
wire _guard6304 = _guard6298 | _guard6303;
wire _guard6305 = early_reset_static_par0_go_out;
wire _guard6306 = _guard6304 & _guard6305;
wire _guard6307 = fsm_out == 1'd0;
wire _guard6308 = cond_wire266_out;
wire _guard6309 = _guard6307 & _guard6308;
wire _guard6310 = fsm_out == 1'd0;
wire _guard6311 = _guard6309 & _guard6310;
wire _guard6312 = fsm_out == 1'd0;
wire _guard6313 = cond_wire267_out;
wire _guard6314 = _guard6312 & _guard6313;
wire _guard6315 = fsm_out == 1'd0;
wire _guard6316 = _guard6314 & _guard6315;
wire _guard6317 = _guard6311 | _guard6316;
wire _guard6318 = early_reset_static_par0_go_out;
wire _guard6319 = _guard6317 & _guard6318;
wire _guard6320 = fsm_out == 1'd0;
wire _guard6321 = cond_wire266_out;
wire _guard6322 = _guard6320 & _guard6321;
wire _guard6323 = fsm_out == 1'd0;
wire _guard6324 = _guard6322 & _guard6323;
wire _guard6325 = fsm_out == 1'd0;
wire _guard6326 = cond_wire267_out;
wire _guard6327 = _guard6325 & _guard6326;
wire _guard6328 = fsm_out == 1'd0;
wire _guard6329 = _guard6327 & _guard6328;
wire _guard6330 = _guard6324 | _guard6329;
wire _guard6331 = early_reset_static_par0_go_out;
wire _guard6332 = _guard6330 & _guard6331;
wire _guard6333 = early_reset_static_par_go_out;
wire _guard6334 = cond_wire9_out;
wire _guard6335 = early_reset_static_par0_go_out;
wire _guard6336 = _guard6334 & _guard6335;
wire _guard6337 = _guard6333 | _guard6336;
wire _guard6338 = early_reset_static_par_go_out;
wire _guard6339 = cond_wire9_out;
wire _guard6340 = early_reset_static_par0_go_out;
wire _guard6341 = _guard6339 & _guard6340;
wire _guard6342 = early_reset_static_par_go_out;
wire _guard6343 = cond_wire72_out;
wire _guard6344 = early_reset_static_par0_go_out;
wire _guard6345 = _guard6343 & _guard6344;
wire _guard6346 = _guard6342 | _guard6345;
wire _guard6347 = early_reset_static_par_go_out;
wire _guard6348 = cond_wire72_out;
wire _guard6349 = early_reset_static_par0_go_out;
wire _guard6350 = _guard6348 & _guard6349;
wire _guard6351 = early_reset_static_par_go_out;
wire _guard6352 = cond_wire204_out;
wire _guard6353 = early_reset_static_par0_go_out;
wire _guard6354 = _guard6352 & _guard6353;
wire _guard6355 = _guard6351 | _guard6354;
wire _guard6356 = early_reset_static_par_go_out;
wire _guard6357 = cond_wire204_out;
wire _guard6358 = early_reset_static_par0_go_out;
wire _guard6359 = _guard6357 & _guard6358;
wire _guard6360 = early_reset_static_par0_go_out;
wire _guard6361 = early_reset_static_par0_go_out;
wire _guard6362 = early_reset_static_par0_go_out;
wire _guard6363 = early_reset_static_par0_go_out;
wire _guard6364 = early_reset_static_par0_go_out;
wire _guard6365 = early_reset_static_par0_go_out;
wire _guard6366 = early_reset_static_par0_go_out;
wire _guard6367 = early_reset_static_par0_go_out;
wire _guard6368 = early_reset_static_par0_go_out;
wire _guard6369 = early_reset_static_par0_go_out;
wire _guard6370 = early_reset_static_par_go_out;
wire _guard6371 = early_reset_static_par0_go_out;
wire _guard6372 = _guard6370 | _guard6371;
wire _guard6373 = early_reset_static_par0_go_out;
wire _guard6374 = early_reset_static_par_go_out;
wire _guard6375 = early_reset_static_par0_go_out;
wire _guard6376 = early_reset_static_par0_go_out;
wire _guard6377 = early_reset_static_par0_go_out;
wire _guard6378 = early_reset_static_par0_go_out;
wire _guard6379 = ~_guard0;
wire _guard6380 = early_reset_static_par0_go_out;
wire _guard6381 = _guard6379 & _guard6380;
wire _guard6382 = early_reset_static_par0_go_out;
wire _guard6383 = early_reset_static_par0_go_out;
wire _guard6384 = early_reset_static_par0_go_out;
wire _guard6385 = early_reset_static_par0_go_out;
wire _guard6386 = early_reset_static_par0_go_out;
wire _guard6387 = ~_guard0;
wire _guard6388 = early_reset_static_par0_go_out;
wire _guard6389 = _guard6387 & _guard6388;
wire _guard6390 = early_reset_static_par0_go_out;
wire _guard6391 = early_reset_static_par0_go_out;
wire _guard6392 = early_reset_static_par0_go_out;
wire _guard6393 = early_reset_static_par0_go_out;
wire _guard6394 = early_reset_static_par0_go_out;
wire _guard6395 = ~_guard0;
wire _guard6396 = early_reset_static_par0_go_out;
wire _guard6397 = _guard6395 & _guard6396;
wire _guard6398 = early_reset_static_par0_go_out;
wire _guard6399 = ~_guard0;
wire _guard6400 = early_reset_static_par0_go_out;
wire _guard6401 = _guard6399 & _guard6400;
wire _guard6402 = early_reset_static_par0_go_out;
wire _guard6403 = ~_guard0;
wire _guard6404 = early_reset_static_par0_go_out;
wire _guard6405 = _guard6403 & _guard6404;
wire _guard6406 = early_reset_static_par0_go_out;
wire _guard6407 = early_reset_static_par0_go_out;
wire _guard6408 = ~_guard0;
wire _guard6409 = early_reset_static_par0_go_out;
wire _guard6410 = _guard6408 & _guard6409;
wire _guard6411 = early_reset_static_par0_go_out;
wire _guard6412 = early_reset_static_par0_go_out;
wire _guard6413 = early_reset_static_par0_go_out;
wire _guard6414 = early_reset_static_par0_go_out;
wire _guard6415 = early_reset_static_par0_go_out;
wire _guard6416 = ~_guard0;
wire _guard6417 = early_reset_static_par0_go_out;
wire _guard6418 = _guard6416 & _guard6417;
wire _guard6419 = early_reset_static_par0_go_out;
wire _guard6420 = early_reset_static_par0_go_out;
wire _guard6421 = early_reset_static_par0_go_out;
wire _guard6422 = early_reset_static_par0_go_out;
wire _guard6423 = early_reset_static_par0_go_out;
wire _guard6424 = early_reset_static_par0_go_out;
wire _guard6425 = early_reset_static_par0_go_out;
wire _guard6426 = early_reset_static_par0_go_out;
wire _guard6427 = early_reset_static_par0_go_out;
wire _guard6428 = early_reset_static_par0_go_out;
wire _guard6429 = early_reset_static_par0_go_out;
wire _guard6430 = early_reset_static_par0_go_out;
wire _guard6431 = early_reset_static_par0_go_out;
wire _guard6432 = ~_guard0;
wire _guard6433 = early_reset_static_par0_go_out;
wire _guard6434 = _guard6432 & _guard6433;
wire _guard6435 = early_reset_static_par0_go_out;
wire _guard6436 = early_reset_static_par0_go_out;
wire _guard6437 = early_reset_static_par0_go_out;
wire _guard6438 = early_reset_static_par0_go_out;
wire _guard6439 = early_reset_static_par0_go_out;
wire _guard6440 = ~_guard0;
wire _guard6441 = early_reset_static_par0_go_out;
wire _guard6442 = _guard6440 & _guard6441;
wire _guard6443 = early_reset_static_par0_go_out;
wire _guard6444 = early_reset_static_par0_go_out;
wire _guard6445 = early_reset_static_par0_go_out;
wire _guard6446 = early_reset_static_par0_go_out;
wire _guard6447 = early_reset_static_par0_go_out;
wire _guard6448 = early_reset_static_par0_go_out;
wire _guard6449 = early_reset_static_par0_go_out;
wire _guard6450 = ~_guard0;
wire _guard6451 = early_reset_static_par0_go_out;
wire _guard6452 = _guard6450 & _guard6451;
wire _guard6453 = ~_guard0;
wire _guard6454 = early_reset_static_par0_go_out;
wire _guard6455 = _guard6453 & _guard6454;
wire _guard6456 = early_reset_static_par0_go_out;
wire _guard6457 = early_reset_static_par0_go_out;
wire _guard6458 = early_reset_static_par0_go_out;
wire _guard6459 = ~_guard0;
wire _guard6460 = early_reset_static_par0_go_out;
wire _guard6461 = _guard6459 & _guard6460;
wire _guard6462 = early_reset_static_par0_go_out;
wire _guard6463 = early_reset_static_par0_go_out;
wire _guard6464 = early_reset_static_par0_go_out;
wire _guard6465 = early_reset_static_par0_go_out;
wire _guard6466 = ~_guard0;
wire _guard6467 = early_reset_static_par0_go_out;
wire _guard6468 = _guard6466 & _guard6467;
wire _guard6469 = ~_guard0;
wire _guard6470 = early_reset_static_par0_go_out;
wire _guard6471 = _guard6469 & _guard6470;
wire _guard6472 = early_reset_static_par0_go_out;
wire _guard6473 = ~_guard0;
wire _guard6474 = early_reset_static_par0_go_out;
wire _guard6475 = _guard6473 & _guard6474;
wire _guard6476 = early_reset_static_par0_go_out;
wire _guard6477 = early_reset_static_par0_go_out;
wire _guard6478 = early_reset_static_par0_go_out;
wire _guard6479 = early_reset_static_par0_go_out;
wire _guard6480 = ~_guard0;
wire _guard6481 = early_reset_static_par0_go_out;
wire _guard6482 = _guard6480 & _guard6481;
wire _guard6483 = early_reset_static_par0_go_out;
wire _guard6484 = early_reset_static_par0_go_out;
wire _guard6485 = wrapper_early_reset_static_par_go_out;
wire _guard6486 = early_reset_static_par_go_out;
wire _guard6487 = early_reset_static_par_go_out;
wire _guard6488 = early_reset_static_par0_go_out;
wire _guard6489 = early_reset_static_par0_go_out;
wire _guard6490 = early_reset_static_par0_go_out;
wire _guard6491 = early_reset_static_par0_go_out;
wire _guard6492 = early_reset_static_par0_go_out;
wire _guard6493 = early_reset_static_par0_go_out;
wire _guard6494 = early_reset_static_par0_go_out;
wire _guard6495 = early_reset_static_par0_go_out;
wire _guard6496 = early_reset_static_par0_go_out;
wire _guard6497 = early_reset_static_par0_go_out;
wire _guard6498 = early_reset_static_par0_go_out;
wire _guard6499 = early_reset_static_par0_go_out;
wire _guard6500 = cond_wire_out;
wire _guard6501 = early_reset_static_par0_go_out;
wire _guard6502 = _guard6500 & _guard6501;
wire _guard6503 = cond_wire_out;
wire _guard6504 = early_reset_static_par0_go_out;
wire _guard6505 = _guard6503 & _guard6504;
wire _guard6506 = cond_wire24_out;
wire _guard6507 = early_reset_static_par0_go_out;
wire _guard6508 = _guard6506 & _guard6507;
wire _guard6509 = cond_wire24_out;
wire _guard6510 = early_reset_static_par0_go_out;
wire _guard6511 = _guard6509 & _guard6510;
wire _guard6512 = cond_wire46_out;
wire _guard6513 = early_reset_static_par0_go_out;
wire _guard6514 = _guard6512 & _guard6513;
wire _guard6515 = cond_wire44_out;
wire _guard6516 = early_reset_static_par0_go_out;
wire _guard6517 = _guard6515 & _guard6516;
wire _guard6518 = fsm_out == 1'd0;
wire _guard6519 = cond_wire44_out;
wire _guard6520 = _guard6518 & _guard6519;
wire _guard6521 = fsm_out == 1'd0;
wire _guard6522 = _guard6520 & _guard6521;
wire _guard6523 = fsm_out == 1'd0;
wire _guard6524 = cond_wire46_out;
wire _guard6525 = _guard6523 & _guard6524;
wire _guard6526 = fsm_out == 1'd0;
wire _guard6527 = _guard6525 & _guard6526;
wire _guard6528 = _guard6522 | _guard6527;
wire _guard6529 = early_reset_static_par0_go_out;
wire _guard6530 = _guard6528 & _guard6529;
wire _guard6531 = fsm_out == 1'd0;
wire _guard6532 = cond_wire44_out;
wire _guard6533 = _guard6531 & _guard6532;
wire _guard6534 = fsm_out == 1'd0;
wire _guard6535 = _guard6533 & _guard6534;
wire _guard6536 = fsm_out == 1'd0;
wire _guard6537 = cond_wire46_out;
wire _guard6538 = _guard6536 & _guard6537;
wire _guard6539 = fsm_out == 1'd0;
wire _guard6540 = _guard6538 & _guard6539;
wire _guard6541 = _guard6535 | _guard6540;
wire _guard6542 = early_reset_static_par0_go_out;
wire _guard6543 = _guard6541 & _guard6542;
wire _guard6544 = fsm_out == 1'd0;
wire _guard6545 = cond_wire44_out;
wire _guard6546 = _guard6544 & _guard6545;
wire _guard6547 = fsm_out == 1'd0;
wire _guard6548 = _guard6546 & _guard6547;
wire _guard6549 = fsm_out == 1'd0;
wire _guard6550 = cond_wire46_out;
wire _guard6551 = _guard6549 & _guard6550;
wire _guard6552 = fsm_out == 1'd0;
wire _guard6553 = _guard6551 & _guard6552;
wire _guard6554 = _guard6548 | _guard6553;
wire _guard6555 = early_reset_static_par0_go_out;
wire _guard6556 = _guard6554 & _guard6555;
wire _guard6557 = cond_wire69_out;
wire _guard6558 = early_reset_static_par0_go_out;
wire _guard6559 = _guard6557 & _guard6558;
wire _guard6560 = cond_wire69_out;
wire _guard6561 = early_reset_static_par0_go_out;
wire _guard6562 = _guard6560 & _guard6561;
wire _guard6563 = cond_wire177_out;
wire _guard6564 = early_reset_static_par0_go_out;
wire _guard6565 = _guard6563 & _guard6564;
wire _guard6566 = cond_wire177_out;
wire _guard6567 = early_reset_static_par0_go_out;
wire _guard6568 = _guard6566 & _guard6567;
wire _guard6569 = cond_wire168_out;
wire _guard6570 = early_reset_static_par0_go_out;
wire _guard6571 = _guard6569 & _guard6570;
wire _guard6572 = cond_wire168_out;
wire _guard6573 = early_reset_static_par0_go_out;
wire _guard6574 = _guard6572 & _guard6573;
wire _guard6575 = cond_wire197_out;
wire _guard6576 = early_reset_static_par0_go_out;
wire _guard6577 = _guard6575 & _guard6576;
wire _guard6578 = cond_wire197_out;
wire _guard6579 = early_reset_static_par0_go_out;
wire _guard6580 = _guard6578 & _guard6579;
wire _guard6581 = cond_wire204_out;
wire _guard6582 = early_reset_static_par0_go_out;
wire _guard6583 = _guard6581 & _guard6582;
wire _guard6584 = cond_wire204_out;
wire _guard6585 = early_reset_static_par0_go_out;
wire _guard6586 = _guard6584 & _guard6585;
wire _guard6587 = cond_wire210_out;
wire _guard6588 = early_reset_static_par0_go_out;
wire _guard6589 = _guard6587 & _guard6588;
wire _guard6590 = cond_wire210_out;
wire _guard6591 = early_reset_static_par0_go_out;
wire _guard6592 = _guard6590 & _guard6591;
wire _guard6593 = early_reset_static_par0_go_out;
wire _guard6594 = early_reset_static_par0_go_out;
wire _guard6595 = early_reset_static_par0_go_out;
wire _guard6596 = early_reset_static_par0_go_out;
wire _guard6597 = early_reset_static_par_go_out;
wire _guard6598 = early_reset_static_par0_go_out;
wire _guard6599 = _guard6597 | _guard6598;
wire _guard6600 = early_reset_static_par0_go_out;
wire _guard6601 = early_reset_static_par_go_out;
wire _guard6602 = early_reset_static_par0_go_out;
wire _guard6603 = early_reset_static_par0_go_out;
wire _guard6604 = early_reset_static_par0_go_out;
wire _guard6605 = early_reset_static_par0_go_out;
wire _guard6606 = early_reset_static_par0_go_out;
wire _guard6607 = early_reset_static_par0_go_out;
wire _guard6608 = early_reset_static_par0_go_out;
wire _guard6609 = early_reset_static_par0_go_out;
wire _guard6610 = early_reset_static_par_go_out;
wire _guard6611 = early_reset_static_par0_go_out;
wire _guard6612 = _guard6610 | _guard6611;
wire _guard6613 = early_reset_static_par_go_out;
wire _guard6614 = early_reset_static_par0_go_out;
wire _guard6615 = early_reset_static_par0_go_out;
wire _guard6616 = early_reset_static_par0_go_out;
wire _guard6617 = early_reset_static_par0_go_out;
wire _guard6618 = early_reset_static_par0_go_out;
wire _guard6619 = early_reset_static_par0_go_out;
wire _guard6620 = early_reset_static_par0_go_out;
wire _guard6621 = early_reset_static_par0_go_out;
wire _guard6622 = ~_guard0;
wire _guard6623 = early_reset_static_par0_go_out;
wire _guard6624 = _guard6622 & _guard6623;
wire _guard6625 = early_reset_static_par0_go_out;
wire _guard6626 = early_reset_static_par0_go_out;
wire _guard6627 = early_reset_static_par0_go_out;
wire _guard6628 = early_reset_static_par0_go_out;
wire _guard6629 = early_reset_static_par0_go_out;
wire _guard6630 = early_reset_static_par0_go_out;
wire _guard6631 = early_reset_static_par0_go_out;
wire _guard6632 = ~_guard0;
wire _guard6633 = early_reset_static_par0_go_out;
wire _guard6634 = _guard6632 & _guard6633;
wire _guard6635 = ~_guard0;
wire _guard6636 = early_reset_static_par0_go_out;
wire _guard6637 = _guard6635 & _guard6636;
wire _guard6638 = early_reset_static_par0_go_out;
wire _guard6639 = early_reset_static_par0_go_out;
wire _guard6640 = early_reset_static_par0_go_out;
wire _guard6641 = ~_guard0;
wire _guard6642 = early_reset_static_par0_go_out;
wire _guard6643 = _guard6641 & _guard6642;
wire _guard6644 = early_reset_static_par0_go_out;
wire _guard6645 = early_reset_static_par0_go_out;
wire _guard6646 = early_reset_static_par0_go_out;
wire _guard6647 = early_reset_static_par0_go_out;
wire _guard6648 = ~_guard0;
wire _guard6649 = early_reset_static_par0_go_out;
wire _guard6650 = _guard6648 & _guard6649;
wire _guard6651 = ~_guard0;
wire _guard6652 = early_reset_static_par0_go_out;
wire _guard6653 = _guard6651 & _guard6652;
wire _guard6654 = early_reset_static_par0_go_out;
wire _guard6655 = early_reset_static_par0_go_out;
wire _guard6656 = ~_guard0;
wire _guard6657 = early_reset_static_par0_go_out;
wire _guard6658 = _guard6656 & _guard6657;
wire _guard6659 = early_reset_static_par0_go_out;
wire _guard6660 = ~_guard0;
wire _guard6661 = early_reset_static_par0_go_out;
wire _guard6662 = _guard6660 & _guard6661;
wire _guard6663 = ~_guard0;
wire _guard6664 = early_reset_static_par0_go_out;
wire _guard6665 = _guard6663 & _guard6664;
wire _guard6666 = early_reset_static_par0_go_out;
wire _guard6667 = early_reset_static_par0_go_out;
wire _guard6668 = early_reset_static_par0_go_out;
wire _guard6669 = early_reset_static_par0_go_out;
wire _guard6670 = ~_guard0;
wire _guard6671 = early_reset_static_par0_go_out;
wire _guard6672 = _guard6670 & _guard6671;
wire _guard6673 = early_reset_static_par0_go_out;
wire _guard6674 = early_reset_static_par0_go_out;
wire _guard6675 = early_reset_static_par0_go_out;
wire _guard6676 = early_reset_static_par0_go_out;
wire _guard6677 = early_reset_static_par0_go_out;
wire _guard6678 = ~_guard0;
wire _guard6679 = early_reset_static_par0_go_out;
wire _guard6680 = _guard6678 & _guard6679;
wire _guard6681 = early_reset_static_par0_go_out;
wire _guard6682 = early_reset_static_par0_go_out;
wire _guard6683 = ~_guard0;
wire _guard6684 = early_reset_static_par0_go_out;
wire _guard6685 = _guard6683 & _guard6684;
wire _guard6686 = early_reset_static_par0_go_out;
wire _guard6687 = ~_guard0;
wire _guard6688 = early_reset_static_par0_go_out;
wire _guard6689 = _guard6687 & _guard6688;
wire _guard6690 = early_reset_static_par0_go_out;
wire _guard6691 = ~_guard0;
wire _guard6692 = early_reset_static_par0_go_out;
wire _guard6693 = _guard6691 & _guard6692;
wire _guard6694 = early_reset_static_par0_go_out;
wire _guard6695 = early_reset_static_par0_go_out;
wire _guard6696 = early_reset_static_par0_go_out;
wire _guard6697 = early_reset_static_par0_go_out;
wire _guard6698 = early_reset_static_par0_go_out;
wire _guard6699 = early_reset_static_par0_go_out;
wire _guard6700 = ~_guard0;
wire _guard6701 = early_reset_static_par0_go_out;
wire _guard6702 = _guard6700 & _guard6701;
wire _guard6703 = early_reset_static_par0_go_out;
wire _guard6704 = ~_guard0;
wire _guard6705 = early_reset_static_par0_go_out;
wire _guard6706 = _guard6704 & _guard6705;
wire _guard6707 = early_reset_static_par0_go_out;
wire _guard6708 = early_reset_static_par0_go_out;
wire _guard6709 = early_reset_static_par0_go_out;
wire _guard6710 = early_reset_static_par0_go_out;
wire _guard6711 = early_reset_static_par0_go_out;
wire _guard6712 = ~_guard0;
wire _guard6713 = early_reset_static_par0_go_out;
wire _guard6714 = _guard6712 & _guard6713;
wire _guard6715 = early_reset_static_par0_go_out;
wire _guard6716 = early_reset_static_par0_go_out;
wire _guard6717 = ~_guard0;
wire _guard6718 = early_reset_static_par0_go_out;
wire _guard6719 = _guard6717 & _guard6718;
wire _guard6720 = early_reset_static_par0_go_out;
wire _guard6721 = early_reset_static_par0_go_out;
wire _guard6722 = early_reset_static_par0_go_out;
wire _guard6723 = early_reset_static_par0_go_out;
wire _guard6724 = early_reset_static_par0_go_out;
wire _guard6725 = cond_wire1_out;
wire _guard6726 = early_reset_static_par0_go_out;
wire _guard6727 = _guard6725 & _guard6726;
wire _guard6728 = cond_wire1_out;
wire _guard6729 = early_reset_static_par0_go_out;
wire _guard6730 = _guard6728 & _guard6729;
wire _guard6731 = cond_wire34_out;
wire _guard6732 = early_reset_static_par0_go_out;
wire _guard6733 = _guard6731 & _guard6732;
wire _guard6734 = cond_wire34_out;
wire _guard6735 = early_reset_static_par0_go_out;
wire _guard6736 = _guard6734 & _guard6735;
wire _guard6737 = cond_wire65_out;
wire _guard6738 = early_reset_static_par0_go_out;
wire _guard6739 = _guard6737 & _guard6738;
wire _guard6740 = cond_wire65_out;
wire _guard6741 = early_reset_static_par0_go_out;
wire _guard6742 = _guard6740 & _guard6741;
wire _guard6743 = cond_wire83_out;
wire _guard6744 = early_reset_static_par0_go_out;
wire _guard6745 = _guard6743 & _guard6744;
wire _guard6746 = cond_wire81_out;
wire _guard6747 = early_reset_static_par0_go_out;
wire _guard6748 = _guard6746 & _guard6747;
wire _guard6749 = fsm_out == 1'd0;
wire _guard6750 = cond_wire81_out;
wire _guard6751 = _guard6749 & _guard6750;
wire _guard6752 = fsm_out == 1'd0;
wire _guard6753 = _guard6751 & _guard6752;
wire _guard6754 = fsm_out == 1'd0;
wire _guard6755 = cond_wire83_out;
wire _guard6756 = _guard6754 & _guard6755;
wire _guard6757 = fsm_out == 1'd0;
wire _guard6758 = _guard6756 & _guard6757;
wire _guard6759 = _guard6753 | _guard6758;
wire _guard6760 = early_reset_static_par0_go_out;
wire _guard6761 = _guard6759 & _guard6760;
wire _guard6762 = fsm_out == 1'd0;
wire _guard6763 = cond_wire81_out;
wire _guard6764 = _guard6762 & _guard6763;
wire _guard6765 = fsm_out == 1'd0;
wire _guard6766 = _guard6764 & _guard6765;
wire _guard6767 = fsm_out == 1'd0;
wire _guard6768 = cond_wire83_out;
wire _guard6769 = _guard6767 & _guard6768;
wire _guard6770 = fsm_out == 1'd0;
wire _guard6771 = _guard6769 & _guard6770;
wire _guard6772 = _guard6766 | _guard6771;
wire _guard6773 = early_reset_static_par0_go_out;
wire _guard6774 = _guard6772 & _guard6773;
wire _guard6775 = fsm_out == 1'd0;
wire _guard6776 = cond_wire81_out;
wire _guard6777 = _guard6775 & _guard6776;
wire _guard6778 = fsm_out == 1'd0;
wire _guard6779 = _guard6777 & _guard6778;
wire _guard6780 = fsm_out == 1'd0;
wire _guard6781 = cond_wire83_out;
wire _guard6782 = _guard6780 & _guard6781;
wire _guard6783 = fsm_out == 1'd0;
wire _guard6784 = _guard6782 & _guard6783;
wire _guard6785 = _guard6779 | _guard6784;
wire _guard6786 = early_reset_static_par0_go_out;
wire _guard6787 = _guard6785 & _guard6786;
wire _guard6788 = cond_wire145_out;
wire _guard6789 = early_reset_static_par0_go_out;
wire _guard6790 = _guard6788 & _guard6789;
wire _guard6791 = cond_wire143_out;
wire _guard6792 = early_reset_static_par0_go_out;
wire _guard6793 = _guard6791 & _guard6792;
wire _guard6794 = fsm_out == 1'd0;
wire _guard6795 = cond_wire143_out;
wire _guard6796 = _guard6794 & _guard6795;
wire _guard6797 = fsm_out == 1'd0;
wire _guard6798 = _guard6796 & _guard6797;
wire _guard6799 = fsm_out == 1'd0;
wire _guard6800 = cond_wire145_out;
wire _guard6801 = _guard6799 & _guard6800;
wire _guard6802 = fsm_out == 1'd0;
wire _guard6803 = _guard6801 & _guard6802;
wire _guard6804 = _guard6798 | _guard6803;
wire _guard6805 = early_reset_static_par0_go_out;
wire _guard6806 = _guard6804 & _guard6805;
wire _guard6807 = fsm_out == 1'd0;
wire _guard6808 = cond_wire143_out;
wire _guard6809 = _guard6807 & _guard6808;
wire _guard6810 = fsm_out == 1'd0;
wire _guard6811 = _guard6809 & _guard6810;
wire _guard6812 = fsm_out == 1'd0;
wire _guard6813 = cond_wire145_out;
wire _guard6814 = _guard6812 & _guard6813;
wire _guard6815 = fsm_out == 1'd0;
wire _guard6816 = _guard6814 & _guard6815;
wire _guard6817 = _guard6811 | _guard6816;
wire _guard6818 = early_reset_static_par0_go_out;
wire _guard6819 = _guard6817 & _guard6818;
wire _guard6820 = fsm_out == 1'd0;
wire _guard6821 = cond_wire143_out;
wire _guard6822 = _guard6820 & _guard6821;
wire _guard6823 = fsm_out == 1'd0;
wire _guard6824 = _guard6822 & _guard6823;
wire _guard6825 = fsm_out == 1'd0;
wire _guard6826 = cond_wire145_out;
wire _guard6827 = _guard6825 & _guard6826;
wire _guard6828 = fsm_out == 1'd0;
wire _guard6829 = _guard6827 & _guard6828;
wire _guard6830 = _guard6824 | _guard6829;
wire _guard6831 = early_reset_static_par0_go_out;
wire _guard6832 = _guard6830 & _guard6831;
wire _guard6833 = cond_wire148_out;
wire _guard6834 = early_reset_static_par0_go_out;
wire _guard6835 = _guard6833 & _guard6834;
wire _guard6836 = cond_wire148_out;
wire _guard6837 = early_reset_static_par0_go_out;
wire _guard6838 = _guard6836 & _guard6837;
wire _guard6839 = cond_wire214_out;
wire _guard6840 = early_reset_static_par0_go_out;
wire _guard6841 = _guard6839 & _guard6840;
wire _guard6842 = cond_wire214_out;
wire _guard6843 = early_reset_static_par0_go_out;
wire _guard6844 = _guard6842 & _guard6843;
wire _guard6845 = cond_wire72_out;
wire _guard6846 = early_reset_static_par0_go_out;
wire _guard6847 = _guard6845 & _guard6846;
wire _guard6848 = cond_wire72_out;
wire _guard6849 = early_reset_static_par0_go_out;
wire _guard6850 = _guard6848 & _guard6849;
wire _guard6851 = early_reset_static_par_go_out;
wire _guard6852 = cond_wire171_out;
wire _guard6853 = early_reset_static_par0_go_out;
wire _guard6854 = _guard6852 & _guard6853;
wire _guard6855 = _guard6851 | _guard6854;
wire _guard6856 = early_reset_static_par_go_out;
wire _guard6857 = cond_wire171_out;
wire _guard6858 = early_reset_static_par0_go_out;
wire _guard6859 = _guard6857 & _guard6858;
wire _guard6860 = cond_wire204_out;
wire _guard6861 = early_reset_static_par0_go_out;
wire _guard6862 = _guard6860 & _guard6861;
wire _guard6863 = cond_wire204_out;
wire _guard6864 = early_reset_static_par0_go_out;
wire _guard6865 = _guard6863 & _guard6864;
wire _guard6866 = early_reset_static_par_go_out;
wire _guard6867 = early_reset_static_par0_go_out;
wire _guard6868 = _guard6866 | _guard6867;
wire _guard6869 = early_reset_static_par_go_out;
wire _guard6870 = early_reset_static_par0_go_out;
wire _guard6871 = early_reset_static_par_go_out;
wire _guard6872 = early_reset_static_par0_go_out;
wire _guard6873 = _guard6871 | _guard6872;
wire _guard6874 = early_reset_static_par0_go_out;
wire _guard6875 = early_reset_static_par_go_out;
wire _guard6876 = early_reset_static_par0_go_out;
wire _guard6877 = early_reset_static_par0_go_out;
wire _guard6878 = early_reset_static_par0_go_out;
wire _guard6879 = early_reset_static_par0_go_out;
wire _guard6880 = early_reset_static_par0_go_out;
wire _guard6881 = early_reset_static_par0_go_out;
wire _guard6882 = early_reset_static_par0_go_out;
wire _guard6883 = early_reset_static_par0_go_out;
wire _guard6884 = early_reset_static_par0_go_out;
wire _guard6885 = early_reset_static_par0_go_out;
wire _guard6886 = early_reset_static_par0_go_out;
wire _guard6887 = early_reset_static_par0_go_out;
wire _guard6888 = early_reset_static_par_go_out;
wire _guard6889 = early_reset_static_par0_go_out;
wire _guard6890 = _guard6888 | _guard6889;
wire _guard6891 = early_reset_static_par0_go_out;
wire _guard6892 = early_reset_static_par_go_out;
wire _guard6893 = early_reset_static_par_go_out;
wire _guard6894 = early_reset_static_par0_go_out;
wire _guard6895 = _guard6893 | _guard6894;
wire _guard6896 = early_reset_static_par0_go_out;
wire _guard6897 = early_reset_static_par_go_out;
wire _guard6898 = early_reset_static_par0_go_out;
wire _guard6899 = early_reset_static_par0_go_out;
wire _guard6900 = early_reset_static_par0_go_out;
wire _guard6901 = early_reset_static_par0_go_out;
wire _guard6902 = early_reset_static_par0_go_out;
wire _guard6903 = early_reset_static_par0_go_out;
wire _guard6904 = early_reset_static_par_go_out;
wire _guard6905 = early_reset_static_par0_go_out;
wire _guard6906 = _guard6904 | _guard6905;
wire _guard6907 = early_reset_static_par0_go_out;
wire _guard6908 = early_reset_static_par_go_out;
wire _guard6909 = ~_guard0;
wire _guard6910 = early_reset_static_par0_go_out;
wire _guard6911 = _guard6909 & _guard6910;
wire _guard6912 = early_reset_static_par0_go_out;
wire _guard6913 = ~_guard0;
wire _guard6914 = early_reset_static_par0_go_out;
wire _guard6915 = _guard6913 & _guard6914;
wire _guard6916 = early_reset_static_par0_go_out;
wire _guard6917 = early_reset_static_par0_go_out;
wire _guard6918 = early_reset_static_par0_go_out;
wire _guard6919 = early_reset_static_par0_go_out;
wire _guard6920 = early_reset_static_par0_go_out;
wire _guard6921 = early_reset_static_par0_go_out;
wire _guard6922 = ~_guard0;
wire _guard6923 = early_reset_static_par0_go_out;
wire _guard6924 = _guard6922 & _guard6923;
wire _guard6925 = early_reset_static_par0_go_out;
wire _guard6926 = early_reset_static_par0_go_out;
wire _guard6927 = ~_guard0;
wire _guard6928 = early_reset_static_par0_go_out;
wire _guard6929 = _guard6927 & _guard6928;
wire _guard6930 = early_reset_static_par0_go_out;
wire _guard6931 = early_reset_static_par0_go_out;
wire _guard6932 = ~_guard0;
wire _guard6933 = early_reset_static_par0_go_out;
wire _guard6934 = _guard6932 & _guard6933;
wire _guard6935 = early_reset_static_par0_go_out;
wire _guard6936 = early_reset_static_par0_go_out;
wire _guard6937 = early_reset_static_par0_go_out;
wire _guard6938 = ~_guard0;
wire _guard6939 = early_reset_static_par0_go_out;
wire _guard6940 = _guard6938 & _guard6939;
wire _guard6941 = early_reset_static_par0_go_out;
wire _guard6942 = early_reset_static_par0_go_out;
wire _guard6943 = early_reset_static_par0_go_out;
wire _guard6944 = ~_guard0;
wire _guard6945 = early_reset_static_par0_go_out;
wire _guard6946 = _guard6944 & _guard6945;
wire _guard6947 = early_reset_static_par0_go_out;
wire _guard6948 = early_reset_static_par0_go_out;
wire _guard6949 = early_reset_static_par0_go_out;
wire _guard6950 = early_reset_static_par0_go_out;
wire _guard6951 = ~_guard0;
wire _guard6952 = early_reset_static_par0_go_out;
wire _guard6953 = _guard6951 & _guard6952;
wire _guard6954 = early_reset_static_par0_go_out;
wire _guard6955 = early_reset_static_par0_go_out;
wire _guard6956 = ~_guard0;
wire _guard6957 = early_reset_static_par0_go_out;
wire _guard6958 = _guard6956 & _guard6957;
wire _guard6959 = ~_guard0;
wire _guard6960 = early_reset_static_par0_go_out;
wire _guard6961 = _guard6959 & _guard6960;
wire _guard6962 = early_reset_static_par0_go_out;
wire _guard6963 = ~_guard0;
wire _guard6964 = early_reset_static_par0_go_out;
wire _guard6965 = _guard6963 & _guard6964;
wire _guard6966 = early_reset_static_par0_go_out;
wire _guard6967 = early_reset_static_par0_go_out;
wire _guard6968 = early_reset_static_par0_go_out;
wire _guard6969 = ~_guard0;
wire _guard6970 = early_reset_static_par0_go_out;
wire _guard6971 = _guard6969 & _guard6970;
wire _guard6972 = early_reset_static_par0_go_out;
wire _guard6973 = early_reset_static_par0_go_out;
wire _guard6974 = ~_guard0;
wire _guard6975 = early_reset_static_par0_go_out;
wire _guard6976 = _guard6974 & _guard6975;
wire _guard6977 = early_reset_static_par0_go_out;
wire _guard6978 = ~_guard0;
wire _guard6979 = early_reset_static_par0_go_out;
wire _guard6980 = _guard6978 & _guard6979;
wire _guard6981 = early_reset_static_par0_go_out;
wire _guard6982 = ~_guard0;
wire _guard6983 = early_reset_static_par0_go_out;
wire _guard6984 = _guard6982 & _guard6983;
wire _guard6985 = ~_guard0;
wire _guard6986 = early_reset_static_par0_go_out;
wire _guard6987 = _guard6985 & _guard6986;
wire _guard6988 = early_reset_static_par0_go_out;
wire _guard6989 = early_reset_static_par0_go_out;
wire _guard6990 = early_reset_static_par0_go_out;
wire _guard6991 = early_reset_static_par0_go_out;
wire _guard6992 = early_reset_static_par0_go_out;
wire _guard6993 = early_reset_static_par0_go_out;
wire _guard6994 = ~_guard0;
wire _guard6995 = early_reset_static_par0_go_out;
wire _guard6996 = _guard6994 & _guard6995;
wire _guard6997 = while_wrapper_early_reset_static_par0_done_out;
wire _guard6998 = ~_guard6997;
wire _guard6999 = fsm0_out == 2'd1;
wire _guard7000 = _guard6998 & _guard6999;
wire _guard7001 = tdcc_go_out;
wire _guard7002 = _guard7000 & _guard7001;
wire _guard7003 = cond_reg_out;
wire _guard7004 = ~_guard7003;
wire _guard7005 = fsm_out == 1'd0;
wire _guard7006 = _guard7004 & _guard7005;
assign depth_plus_20_left = depth;
assign depth_plus_20_right = 32'd20;
assign min_depth_4_plus_5_left = min_depth_4_out;
assign min_depth_4_plus_5_right = 32'd5;
assign pe_1_4_mul_ready =
  _guard7 ? 1'd1 :
  _guard10 ? 1'd0 :
  1'd0;
assign pe_1_4_clk = clk;
assign pe_1_4_top =
  _guard23 ? top_1_4_out :
  32'd0;
assign pe_1_4_left =
  _guard36 ? left_1_4_out :
  32'd0;
assign pe_1_4_reset = reset;
assign pe_1_4_go = _guard49;
assign pe_1_7_mul_ready =
  _guard52 ? 1'd1 :
  _guard55 ? 1'd0 :
  1'd0;
assign pe_1_7_clk = clk;
assign pe_1_7_top =
  _guard68 ? top_1_7_out :
  32'd0;
assign pe_1_7_left =
  _guard81 ? left_1_7_out :
  32'd0;
assign pe_1_7_reset = reset;
assign pe_1_7_go = _guard94;
assign top_2_4_write_en = _guard97;
assign top_2_4_clk = clk;
assign top_2_4_reset = reset;
assign top_2_4_in = top_1_4_out;
assign left_2_4_write_en = _guard103;
assign left_2_4_clk = clk;
assign left_2_4_reset = reset;
assign left_2_4_in = left_2_3_out;
assign top_3_5_write_en = _guard109;
assign top_3_5_clk = clk;
assign top_3_5_reset = reset;
assign top_3_5_in = top_2_5_out;
assign top_3_6_write_en = _guard115;
assign top_3_6_clk = clk;
assign top_3_6_reset = reset;
assign top_3_6_in = top_2_6_out;
assign left_4_0_write_en = _guard121;
assign left_4_0_clk = clk;
assign left_4_0_reset = reset;
assign left_4_0_in = l4_read_data;
assign top_4_4_write_en = _guard127;
assign top_4_4_clk = clk;
assign top_4_4_reset = reset;
assign top_4_4_in = top_3_4_out;
assign pe_5_2_mul_ready =
  _guard133 ? 1'd1 :
  _guard136 ? 1'd0 :
  1'd0;
assign pe_5_2_clk = clk;
assign pe_5_2_top =
  _guard149 ? top_5_2_out :
  32'd0;
assign pe_5_2_left =
  _guard162 ? left_5_2_out :
  32'd0;
assign pe_5_2_reset = reset;
assign pe_5_2_go = _guard175;
assign top_6_1_write_en = _guard178;
assign top_6_1_clk = clk;
assign top_6_1_reset = reset;
assign top_6_1_in = top_5_1_out;
assign left_6_2_write_en = _guard184;
assign left_6_2_clk = clk;
assign left_6_2_reset = reset;
assign left_6_2_in = left_6_1_out;
assign top_6_3_write_en = _guard190;
assign top_6_3_clk = clk;
assign top_6_3_reset = reset;
assign top_6_3_in = top_5_3_out;
assign left_6_4_write_en = _guard196;
assign left_6_4_clk = clk;
assign left_6_4_reset = reset;
assign left_6_4_in = left_6_3_out;
assign top_7_0_write_en = _guard202;
assign top_7_0_clk = clk;
assign top_7_0_reset = reset;
assign top_7_0_in = top_6_0_out;
assign t3_add_left = 4'd1;
assign t3_add_right = t3_idx_out;
assign l1_add_left = 4'd1;
assign l1_add_right = l1_idx_out;
assign idx_between_depth_plus_8_depth_plus_9_reg_write_en = _guard220;
assign idx_between_depth_plus_8_depth_plus_9_reg_clk = clk;
assign idx_between_depth_plus_8_depth_plus_9_reg_reset = reset;
assign idx_between_depth_plus_8_depth_plus_9_reg_in =
  _guard221 ? idx_between_depth_plus_8_depth_plus_9_comb_out :
  _guard222 ? 1'd0 :
  'x;
assign idx_between_11_depth_plus_11_reg_write_en = _guard225;
assign idx_between_11_depth_plus_11_reg_clk = clk;
assign idx_between_11_depth_plus_11_reg_reset = reset;
assign idx_between_11_depth_plus_11_reg_in =
  _guard226 ? idx_between_11_depth_plus_11_comb_out :
  _guard227 ? 1'd0 :
  'x;
assign idx_between_depth_plus_18_depth_plus_19_comb_left = index_ge_depth_plus_18_out;
assign idx_between_depth_plus_18_depth_plus_19_comb_right = index_lt_depth_plus_19_out;
assign index_lt_min_depth_4_plus_8_left = idx_add_out;
assign index_lt_min_depth_4_plus_8_right = min_depth_4_plus_8_out;
assign index_ge_15_left = idx_add_out;
assign index_ge_15_right = 32'd15;
assign cond_wire3_in =
  _guard234 ? idx_between_depth_plus_5_depth_plus_6_reg_out :
  _guard237 ? cond3_out :
  1'd0;
assign cond_wire30_in =
  _guard240 ? cond30_out :
  _guard241 ? idx_between_7_min_depth_4_plus_7_reg_out :
  1'd0;
assign cond_wire38_in =
  _guard242 ? idx_between_depth_plus_12_depth_plus_13_reg_out :
  _guard245 ? cond38_out :
  1'd0;
assign cond_wire39_in =
  _guard246 ? idx_between_1_depth_plus_1_reg_out :
  _guard249 ? cond39_out :
  1'd0;
assign cond_wire47_in =
  _guard250 ? idx_between_depth_plus_7_depth_plus_8_reg_out :
  _guard253 ? cond47_out :
  1'd0;
assign cond53_write_en = _guard254;
assign cond53_clk = clk;
assign cond53_reset = reset;
assign cond53_in =
  _guard255 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond_wire54_in =
  _guard258 ? cond54_out :
  _guard259 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond65_write_en = _guard260;
assign cond65_clk = clk;
assign cond65_reset = reset;
assign cond65_in =
  _guard261 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond70_write_en = _guard262;
assign cond70_clk = clk;
assign cond70_reset = reset;
assign cond70_in =
  _guard263 ? idx_between_13_depth_plus_13_reg_out :
  1'd0;
assign cond71_write_en = _guard264;
assign cond71_clk = clk;
assign cond71_reset = reset;
assign cond71_in =
  _guard265 ? idx_between_depth_plus_13_depth_plus_14_reg_out :
  1'd0;
assign cond_wire89_in =
  _guard266 ? idx_between_7_min_depth_4_plus_7_reg_out :
  _guard269 ? cond89_out :
  1'd0;
assign cond_wire90_in =
  _guard270 ? idx_between_7_depth_plus_7_reg_out :
  _guard273 ? cond90_out :
  1'd0;
assign cond_wire103_in =
  _guard276 ? cond103_out :
  _guard277 ? idx_between_14_depth_plus_14_reg_out :
  1'd0;
assign cond_wire131_in =
  _guard280 ? cond131_out :
  _guard281 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond_wire164_in =
  _guard282 ? idx_between_11_depth_plus_11_reg_out :
  _guard285 ? cond164_out :
  1'd0;
assign cond167_write_en = _guard286;
assign cond167_clk = clk;
assign cond167_reset = reset;
assign cond167_in =
  _guard287 ? idx_between_12_min_depth_4_plus_12_reg_out :
  1'd0;
assign cond181_write_en = _guard288;
assign cond181_clk = clk;
assign cond181_reset = reset;
assign cond181_in =
  _guard289 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire185_in =
  _guard290 ? idx_between_9_depth_plus_9_reg_out :
  _guard293 ? cond185_out :
  1'd0;
assign cond_wire193_in =
  _guard294 ? idx_between_11_depth_plus_11_reg_out :
  _guard297 ? cond193_out :
  1'd0;
assign cond202_write_en = _guard298;
assign cond202_clk = clk;
assign cond202_reset = reset;
assign cond202_in =
  _guard299 ? idx_between_17_depth_plus_17_reg_out :
  1'd0;
assign cond_wire204_in =
  _guard302 ? cond204_out :
  _guard303 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire224_in =
  _guard306 ? cond224_out :
  _guard307 ? idx_between_depth_plus_15_depth_plus_16_reg_out :
  1'd0;
assign cond227_write_en = _guard308;
assign cond227_clk = clk;
assign cond227_reset = reset;
assign cond227_in =
  _guard309 ? idx_between_16_depth_plus_16_reg_out :
  1'd0;
assign cond230_write_en = _guard310;
assign cond230_clk = clk;
assign cond230_reset = reset;
assign cond230_in =
  _guard311 ? idx_between_13_depth_plus_13_reg_out :
  1'd0;
assign cond_wire234_in =
  _guard312 ? idx_between_14_depth_plus_14_reg_out :
  _guard315 ? cond234_out :
  1'd0;
assign cond239_write_en = _guard316;
assign cond239_clk = clk;
assign cond239_reset = reset;
assign cond239_in =
  _guard317 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire240_in =
  _guard320 ? cond240_out :
  _guard321 ? idx_between_12_depth_plus_12_reg_out :
  1'd0;
assign cond263_write_en = _guard322;
assign cond263_clk = clk;
assign cond263_reset = reset;
assign cond263_in =
  _guard323 ? idx_between_14_depth_plus_14_reg_out :
  1'd0;
assign depth_plus_16_left =
  _guard324 ? depth :
  _guard325 ? 32'd20 :
  'x;
assign depth_plus_16_right =
  _guard326 ? depth :
  _guard327 ? 32'd16 :
  'x;
assign min_depth_4_plus_10_left = min_depth_4_out;
assign min_depth_4_plus_10_right = 32'd10;
assign left_0_3_write_en = _guard332;
assign left_0_3_clk = clk;
assign left_0_3_reset = reset;
assign left_0_3_in = left_0_2_out;
assign left_0_4_write_en = _guard338;
assign left_0_4_clk = clk;
assign left_0_4_reset = reset;
assign left_0_4_in = left_0_3_out;
assign top_1_0_write_en = _guard344;
assign top_1_0_clk = clk;
assign top_1_0_reset = reset;
assign top_1_0_in = top_0_0_out;
assign pe_1_2_mul_ready =
  _guard350 ? 1'd1 :
  _guard353 ? 1'd0 :
  1'd0;
assign pe_1_2_clk = clk;
assign pe_1_2_top =
  _guard366 ? top_1_2_out :
  32'd0;
assign pe_1_2_left =
  _guard379 ? left_1_2_out :
  32'd0;
assign pe_1_2_reset = reset;
assign pe_1_2_go = _guard392;
assign pe_1_3_mul_ready =
  _guard395 ? 1'd1 :
  _guard398 ? 1'd0 :
  1'd0;
assign pe_1_3_clk = clk;
assign pe_1_3_top =
  _guard411 ? top_1_3_out :
  32'd0;
assign pe_1_3_left =
  _guard424 ? left_1_3_out :
  32'd0;
assign pe_1_3_reset = reset;
assign pe_1_3_go = _guard437;
assign left_1_3_write_en = _guard440;
assign left_1_3_clk = clk;
assign left_1_3_reset = reset;
assign left_1_3_in = left_1_2_out;
assign left_2_6_write_en = _guard446;
assign left_2_6_clk = clk;
assign left_2_6_reset = reset;
assign left_2_6_in = left_2_5_out;
assign top_4_7_write_en = _guard452;
assign top_4_7_clk = clk;
assign top_4_7_reset = reset;
assign top_4_7_in = top_3_7_out;
assign left_5_1_write_en = _guard458;
assign left_5_1_clk = clk;
assign left_5_1_reset = reset;
assign left_5_1_in = left_5_0_out;
assign left_5_3_write_en = _guard464;
assign left_5_3_clk = clk;
assign left_5_3_reset = reset;
assign left_5_3_in = left_5_2_out;
assign pe_6_4_mul_ready =
  _guard470 ? 1'd1 :
  _guard473 ? 1'd0 :
  1'd0;
assign pe_6_4_clk = clk;
assign pe_6_4_top =
  _guard486 ? top_6_4_out :
  32'd0;
assign pe_6_4_left =
  _guard499 ? left_6_4_out :
  32'd0;
assign pe_6_4_reset = reset;
assign pe_6_4_go = _guard512;
assign top_6_7_write_en = _guard515;
assign top_6_7_clk = clk;
assign top_6_7_reset = reset;
assign top_6_7_in = top_5_7_out;
assign pe_7_3_mul_ready =
  _guard521 ? 1'd1 :
  _guard524 ? 1'd0 :
  1'd0;
assign pe_7_3_clk = clk;
assign pe_7_3_top =
  _guard537 ? top_7_3_out :
  32'd0;
assign pe_7_3_left =
  _guard550 ? left_7_3_out :
  32'd0;
assign pe_7_3_reset = reset;
assign pe_7_3_go = _guard563;
assign left_7_4_write_en = _guard566;
assign left_7_4_clk = clk;
assign left_7_4_reset = reset;
assign left_7_4_in = left_7_3_out;
assign left_7_6_write_en = _guard572;
assign left_7_6_clk = clk;
assign left_7_6_reset = reset;
assign left_7_6_in = left_7_5_out;
assign top_7_7_write_en = _guard578;
assign top_7_7_clk = clk;
assign top_7_7_reset = reset;
assign top_7_7_in = top_6_7_out;
assign l3_idx_write_en = _guard586;
assign l3_idx_clk = clk;
assign l3_idx_reset = reset;
assign l3_idx_in =
  _guard589 ? l3_add_out :
  _guard590 ? 4'd0 :
  'x;
assign l7_idx_write_en = _guard595;
assign l7_idx_clk = clk;
assign l7_idx_reset = reset;
assign l7_idx_in =
  _guard596 ? 4'd0 :
  _guard599 ? l7_add_out :
  'x;
assign idx_between_depth_plus_12_depth_plus_13_comb_left = index_ge_depth_plus_12_out;
assign idx_between_depth_plus_12_depth_plus_13_comb_right = index_lt_depth_plus_13_out;
assign index_lt_depth_plus_9_left = idx_add_out;
assign index_lt_depth_plus_9_right = depth_plus_9_out;
assign index_lt_min_depth_4_plus_2_left = idx_add_out;
assign index_lt_min_depth_4_plus_2_right = min_depth_4_plus_2_out;
assign index_lt_min_depth_4_plus_3_left = idx_add_out;
assign index_lt_min_depth_4_plus_3_right = min_depth_4_plus_3_out;
assign index_lt_depth_plus_6_left = idx_add_out;
assign index_lt_depth_plus_6_right = depth_plus_6_out;
assign index_ge_8_left = idx_add_out;
assign index_ge_8_right = 32'd8;
assign idx_between_8_min_depth_4_plus_8_reg_write_en = _guard614;
assign idx_between_8_min_depth_4_plus_8_reg_clk = clk;
assign idx_between_8_min_depth_4_plus_8_reg_reset = reset;
assign idx_between_8_min_depth_4_plus_8_reg_in =
  _guard615 ? idx_between_8_min_depth_4_plus_8_comb_out :
  _guard616 ? 1'd0 :
  'x;
assign index_lt_depth_plus_20_left = idx_add_out;
assign index_lt_depth_plus_20_right = depth_plus_20_out;
assign idx_between_depth_plus_6_depth_plus_7_reg_write_en = _guard621;
assign idx_between_depth_plus_6_depth_plus_7_reg_clk = clk;
assign idx_between_depth_plus_6_depth_plus_7_reg_reset = reset;
assign idx_between_depth_plus_6_depth_plus_7_reg_in =
  _guard622 ? idx_between_depth_plus_6_depth_plus_7_comb_out :
  _guard623 ? 1'd0 :
  'x;
assign idx_between_depth_plus_15_depth_plus_16_comb_left = index_ge_depth_plus_15_out;
assign idx_between_depth_plus_15_depth_plus_16_comb_right = index_lt_depth_plus_16_out;
assign index_ge_14_left = idx_add_out;
assign index_ge_14_right = 32'd14;
assign t2_addr0 =
  _guard630 ? t2_idx_out :
  4'd0;
assign out_mem_4_write_data =
  _guard633 ? pe_4_0_out :
  _guard636 ? pe_4_5_out :
  _guard639 ? pe_4_6_out :
  _guard642 ? pe_4_2_out :
  _guard645 ? pe_4_4_out :
  _guard648 ? pe_4_7_out :
  _guard651 ? pe_4_3_out :
  _guard654 ? pe_4_1_out :
  32'd0;
assign done = _guard655;
assign l5_addr0 =
  _guard658 ? l5_idx_out :
  4'd0;
assign l0_addr0 =
  _guard661 ? l0_idx_out :
  4'd0;
assign out_mem_1_addr0 =
  _guard664 ? 32'd5 :
  _guard667 ? 32'd0 :
  _guard670 ? 32'd7 :
  _guard673 ? 32'd6 :
  _guard676 ? 32'd2 :
  _guard679 ? 32'd1 :
  _guard682 ? 32'd3 :
  _guard685 ? 32'd4 :
  32'd0;
assign out_mem_5_addr0 =
  _guard688 ? 32'd5 :
  _guard691 ? 32'd0 :
  _guard694 ? 32'd7 :
  _guard697 ? 32'd6 :
  _guard700 ? 32'd2 :
  _guard703 ? 32'd1 :
  _guard706 ? 32'd3 :
  _guard709 ? 32'd4 :
  32'd0;
assign out_mem_5_write_data =
  _guard712 ? pe_5_2_out :
  _guard715 ? pe_5_0_out :
  _guard718 ? pe_5_4_out :
  _guard721 ? pe_5_1_out :
  _guard724 ? pe_5_7_out :
  _guard727 ? pe_5_3_out :
  _guard730 ? pe_5_5_out :
  _guard733 ? pe_5_6_out :
  32'd0;
assign l6_addr0 =
  _guard736 ? l6_idx_out :
  4'd0;
assign out_mem_0_write_data =
  _guard739 ? pe_0_1_out :
  _guard742 ? pe_0_7_out :
  _guard745 ? pe_0_3_out :
  _guard748 ? pe_0_5_out :
  _guard751 ? pe_0_2_out :
  _guard754 ? pe_0_4_out :
  _guard757 ? pe_0_0_out :
  _guard760 ? pe_0_6_out :
  32'd0;
assign out_mem_6_addr0 =
  _guard763 ? 32'd5 :
  _guard766 ? 32'd0 :
  _guard769 ? 32'd7 :
  _guard772 ? 32'd6 :
  _guard775 ? 32'd2 :
  _guard778 ? 32'd1 :
  _guard781 ? 32'd3 :
  _guard784 ? 32'd4 :
  32'd0;
assign out_mem_3_write_data =
  _guard787 ? pe_3_4_out :
  _guard790 ? pe_3_7_out :
  _guard793 ? pe_3_2_out :
  _guard796 ? pe_3_5_out :
  _guard799 ? pe_3_6_out :
  _guard802 ? pe_3_0_out :
  _guard805 ? pe_3_1_out :
  _guard808 ? pe_3_3_out :
  32'd0;
assign t5_addr0 =
  _guard811 ? t5_idx_out :
  4'd0;
assign l1_addr0 =
  _guard814 ? l1_idx_out :
  4'd0;
assign out_mem_5_write_en = _guard863;
assign out_mem_7_addr0 =
  _guard866 ? 32'd5 :
  _guard869 ? 32'd0 :
  _guard872 ? 32'd7 :
  _guard875 ? 32'd6 :
  _guard878 ? 32'd2 :
  _guard881 ? 32'd1 :
  _guard884 ? 32'd3 :
  _guard887 ? 32'd4 :
  32'd0;
assign t4_addr0 =
  _guard890 ? t4_idx_out :
  4'd0;
assign t6_addr0 =
  _guard893 ? t6_idx_out :
  4'd0;
assign out_mem_7_write_en = _guard942;
assign out_mem_4_addr0 =
  _guard945 ? 32'd5 :
  _guard948 ? 32'd0 :
  _guard951 ? 32'd7 :
  _guard954 ? 32'd6 :
  _guard957 ? 32'd2 :
  _guard960 ? 32'd1 :
  _guard963 ? 32'd3 :
  _guard966 ? 32'd4 :
  32'd0;
assign l3_addr0 =
  _guard969 ? l3_idx_out :
  4'd0;
assign out_mem_2_write_data =
  _guard972 ? pe_2_7_out :
  _guard975 ? pe_2_4_out :
  _guard978 ? pe_2_1_out :
  _guard981 ? pe_2_3_out :
  _guard984 ? pe_2_5_out :
  _guard987 ? pe_2_6_out :
  _guard990 ? pe_2_0_out :
  _guard993 ? pe_2_2_out :
  32'd0;
assign l4_addr0 =
  _guard996 ? l4_idx_out :
  4'd0;
assign l7_addr0 =
  _guard999 ? l7_idx_out :
  4'd0;
assign out_mem_1_write_data =
  _guard1002 ? pe_1_4_out :
  _guard1005 ? pe_1_7_out :
  _guard1008 ? pe_1_2_out :
  _guard1011 ? pe_1_3_out :
  _guard1014 ? pe_1_0_out :
  _guard1017 ? pe_1_6_out :
  _guard1020 ? pe_1_5_out :
  _guard1023 ? pe_1_1_out :
  32'd0;
assign out_mem_1_write_en = _guard1072;
assign out_mem_4_write_en = _guard1121;
assign t0_addr0 =
  _guard1124 ? t0_idx_out :
  4'd0;
assign t1_addr0 =
  _guard1127 ? t1_idx_out :
  4'd0;
assign out_mem_0_write_en = _guard1176;
assign out_mem_2_write_en = _guard1225;
assign out_mem_3_write_en = _guard1274;
assign out_mem_6_write_data =
  _guard1277 ? pe_6_4_out :
  _guard1280 ? pe_6_0_out :
  _guard1283 ? pe_6_1_out :
  _guard1286 ? pe_6_5_out :
  _guard1289 ? pe_6_2_out :
  _guard1292 ? pe_6_3_out :
  _guard1295 ? pe_6_7_out :
  _guard1298 ? pe_6_6_out :
  32'd0;
assign out_mem_6_write_en = _guard1347;
assign out_mem_7_write_data =
  _guard1350 ? pe_7_3_out :
  _guard1353 ? pe_7_4_out :
  _guard1356 ? pe_7_0_out :
  _guard1359 ? pe_7_5_out :
  _guard1362 ? pe_7_6_out :
  _guard1365 ? pe_7_1_out :
  _guard1368 ? pe_7_2_out :
  _guard1371 ? pe_7_7_out :
  32'd0;
assign l2_addr0 =
  _guard1374 ? l2_idx_out :
  4'd0;
assign out_mem_0_addr0 =
  _guard1377 ? 32'd5 :
  _guard1380 ? 32'd0 :
  _guard1383 ? 32'd7 :
  _guard1386 ? 32'd6 :
  _guard1389 ? 32'd2 :
  _guard1392 ? 32'd1 :
  _guard1395 ? 32'd3 :
  _guard1398 ? 32'd4 :
  32'd0;
assign out_mem_3_addr0 =
  _guard1401 ? 32'd5 :
  _guard1404 ? 32'd0 :
  _guard1407 ? 32'd7 :
  _guard1410 ? 32'd6 :
  _guard1413 ? 32'd2 :
  _guard1416 ? 32'd1 :
  _guard1419 ? 32'd3 :
  _guard1422 ? 32'd4 :
  32'd0;
assign t3_addr0 =
  _guard1425 ? t3_idx_out :
  4'd0;
assign t7_addr0 =
  _guard1428 ? t7_idx_out :
  4'd0;
assign out_mem_2_addr0 =
  _guard1431 ? 32'd5 :
  _guard1434 ? 32'd0 :
  _guard1437 ? 32'd7 :
  _guard1440 ? 32'd6 :
  _guard1443 ? 32'd2 :
  _guard1446 ? 32'd1 :
  _guard1449 ? 32'd3 :
  _guard1452 ? 32'd4 :
  32'd0;
assign cond_wire0_in =
  _guard1453 ? idx_between_1_min_depth_4_plus_1_reg_out :
  _guard1456 ? cond0_out :
  1'd0;
assign cond_wire4_in =
  _guard1459 ? cond4_out :
  _guard1460 ? idx_between_1_depth_plus_1_reg_out :
  1'd0;
assign cond6_write_en = _guard1461;
assign cond6_clk = clk;
assign cond6_reset = reset;
assign cond6_in =
  _guard1462 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond_wire13_in =
  _guard1465 ? cond13_out :
  _guard1466 ? idx_between_depth_plus_7_depth_plus_8_reg_out :
  1'd0;
assign cond_wire16_in =
  _guard1469 ? cond16_out :
  _guard1470 ? idx_between_4_depth_plus_4_reg_out :
  1'd0;
assign cond30_write_en = _guard1471;
assign cond30_clk = clk;
assign cond30_reset = reset;
assign cond30_in =
  _guard1472 ? idx_between_7_min_depth_4_plus_7_reg_out :
  1'd0;
assign cond_wire32_in =
  _guard1473 ? idx_between_11_depth_plus_11_reg_out :
  _guard1476 ? cond32_out :
  1'd0;
assign cond_wire40_in =
  _guard1479 ? cond40_out :
  _guard1480 ? idx_between_2_min_depth_4_plus_2_reg_out :
  1'd0;
assign cond44_write_en = _guard1481;
assign cond44_clk = clk;
assign cond44_reset = reset;
assign cond44_in =
  _guard1482 ? idx_between_3_min_depth_4_plus_3_reg_out :
  1'd0;
assign cond45_write_en = _guard1483;
assign cond45_clk = clk;
assign cond45_reset = reset;
assign cond45_in =
  _guard1484 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond_wire73_in =
  _guard1487 ? cond73_out :
  _guard1488 ? idx_between_3_min_depth_4_plus_3_reg_out :
  1'd0;
assign cond81_write_en = _guard1489;
assign cond81_clk = clk;
assign cond81_reset = reset;
assign cond81_in =
  _guard1490 ? idx_between_5_min_depth_4_plus_5_reg_out :
  1'd0;
assign cond98_write_en = _guard1491;
assign cond98_clk = clk;
assign cond98_reset = reset;
assign cond98_in =
  _guard1492 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond100_write_en = _guard1493;
assign cond100_clk = clk;
assign cond100_reset = reset;
assign cond100_in =
  _guard1494 ? idx_between_depth_plus_13_depth_plus_14_reg_out :
  1'd0;
assign cond_wire101_in =
  _guard1495 ? idx_between_10_min_depth_4_plus_10_reg_out :
  _guard1498 ? cond101_out :
  1'd0;
assign cond107_write_en = _guard1499;
assign cond107_clk = clk;
assign cond107_reset = reset;
assign cond107_in =
  _guard1500 ? idx_between_4_depth_plus_4_reg_out :
  1'd0;
assign cond_wire107_in =
  _guard1503 ? cond107_out :
  _guard1504 ? idx_between_4_depth_plus_4_reg_out :
  1'd0;
assign cond115_write_en = _guard1505;
assign cond115_clk = clk;
assign cond115_reset = reset;
assign cond115_in =
  _guard1506 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire121_in =
  _guard1509 ? cond121_out :
  _guard1510 ? idx_between_depth_plus_11_depth_plus_12_reg_out :
  1'd0;
assign cond_wire127_in =
  _guard1511 ? idx_between_9_depth_plus_9_reg_out :
  _guard1514 ? cond127_out :
  1'd0;
assign cond_wire144_in =
  _guard1515 ? idx_between_6_depth_plus_6_reg_out :
  _guard1518 ? cond144_out :
  1'd0;
assign cond149_write_en = _guard1519;
assign cond149_clk = clk;
assign cond149_reset = reset;
assign cond149_in =
  _guard1520 ? idx_between_11_depth_plus_11_reg_out :
  1'd0;
assign cond150_write_en = _guard1521;
assign cond150_clk = clk;
assign cond150_reset = reset;
assign cond150_in =
  _guard1522 ? idx_between_depth_plus_11_depth_plus_12_reg_out :
  1'd0;
assign cond_wire160_in =
  _guard1525 ? cond160_out :
  _guard1526 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond169_write_en = _guard1527;
assign cond169_clk = clk;
assign cond169_reset = reset;
assign cond169_in =
  _guard1528 ? idx_between_16_depth_plus_16_reg_out :
  1'd0;
assign cond179_write_en = _guard1529;
assign cond179_clk = clk;
assign cond179_reset = reset;
assign cond179_in =
  _guard1530 ? idx_between_depth_plus_11_depth_plus_12_reg_out :
  1'd0;
assign cond193_write_en = _guard1531;
assign cond193_clk = clk;
assign cond193_reset = reset;
assign cond193_in =
  _guard1532 ? idx_between_11_depth_plus_11_reg_out :
  1'd0;
assign cond_wire208_in =
  _guard1535 ? cond208_out :
  _guard1536 ? idx_between_depth_plus_11_depth_plus_12_reg_out :
  1'd0;
assign cond214_write_en = _guard1537;
assign cond214_clk = clk;
assign cond214_reset = reset;
assign cond214_in =
  _guard1538 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond_wire230_in =
  _guard1541 ? cond230_out :
  _guard1542 ? idx_between_13_depth_plus_13_reg_out :
  1'd0;
assign cond236_write_en = _guard1543;
assign cond236_clk = clk;
assign cond236_reset = reset;
assign cond236_in =
  _guard1544 ? idx_between_depth_plus_18_depth_plus_19_reg_out :
  1'd0;
assign cond_wire239_in =
  _guard1547 ? cond239_out :
  _guard1548 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond245_write_en = _guard1549;
assign cond245_clk = clk;
assign cond245_reset = reset;
assign cond245_in =
  _guard1550 ? idx_between_depth_plus_13_depth_plus_14_reg_out :
  1'd0;
assign cond255_write_en = _guard1551;
assign cond255_clk = clk;
assign cond255_reset = reset;
assign cond255_in =
  _guard1552 ? idx_between_12_depth_plus_12_reg_out :
  1'd0;
assign cond_wire261_in =
  _guard1553 ? idx_between_depth_plus_17_depth_plus_18_reg_out :
  _guard1556 ? cond261_out :
  1'd0;
assign fsm_write_en = _guard1559;
assign fsm_clk = clk;
assign fsm_reset = reset;
assign fsm_in =
  _guard1562 ? adder_out :
  _guard1569 ? 1'd0 :
  _guard1572 ? adder0_out :
  1'd0;
assign adder_left =
  _guard1573 ? fsm_out :
  1'd0;
assign adder_right = _guard1574;
assign early_reset_static_par0_go_in = _guard1575;
assign depth_plus_10_left = depth;
assign depth_plus_10_right = 32'd10;
assign depth_plus_4_left = depth;
assign depth_plus_4_right = 32'd4;
assign top_0_6_write_en = _guard1582;
assign top_0_6_clk = clk;
assign top_0_6_reset = reset;
assign top_0_6_in = t6_read_data;
assign left_1_4_write_en = _guard1588;
assign left_1_4_clk = clk;
assign left_1_4_reset = reset;
assign left_1_4_in = left_1_3_out;
assign top_1_5_write_en = _guard1594;
assign top_1_5_clk = clk;
assign top_1_5_reset = reset;
assign top_1_5_in = top_0_5_out;
assign left_1_5_write_en = _guard1600;
assign left_1_5_clk = clk;
assign left_1_5_reset = reset;
assign left_1_5_in = left_1_4_out;
assign pe_3_4_mul_ready =
  _guard1606 ? 1'd1 :
  _guard1609 ? 1'd0 :
  1'd0;
assign pe_3_4_clk = clk;
assign pe_3_4_top =
  _guard1622 ? top_3_4_out :
  32'd0;
assign pe_3_4_left =
  _guard1635 ? left_3_4_out :
  32'd0;
assign pe_3_4_reset = reset;
assign pe_3_4_go = _guard1648;
assign pe_3_7_mul_ready =
  _guard1651 ? 1'd1 :
  _guard1654 ? 1'd0 :
  1'd0;
assign pe_3_7_clk = clk;
assign pe_3_7_top =
  _guard1667 ? top_3_7_out :
  32'd0;
assign pe_3_7_left =
  _guard1680 ? left_3_7_out :
  32'd0;
assign pe_3_7_reset = reset;
assign pe_3_7_go = _guard1693;
assign pe_4_0_mul_ready =
  _guard1696 ? 1'd1 :
  _guard1699 ? 1'd0 :
  1'd0;
assign pe_4_0_clk = clk;
assign pe_4_0_top =
  _guard1712 ? top_4_0_out :
  32'd0;
assign pe_4_0_left =
  _guard1725 ? left_4_0_out :
  32'd0;
assign pe_4_0_reset = reset;
assign pe_4_0_go = _guard1738;
assign left_4_2_write_en = _guard1741;
assign left_4_2_clk = clk;
assign left_4_2_reset = reset;
assign left_4_2_in = left_4_1_out;
assign pe_5_0_mul_ready =
  _guard1747 ? 1'd1 :
  _guard1750 ? 1'd0 :
  1'd0;
assign pe_5_0_clk = clk;
assign pe_5_0_top =
  _guard1763 ? top_5_0_out :
  32'd0;
assign pe_5_0_left =
  _guard1776 ? left_5_0_out :
  32'd0;
assign pe_5_0_reset = reset;
assign pe_5_0_go = _guard1789;
assign left_5_6_write_en = _guard1792;
assign left_5_6_clk = clk;
assign left_5_6_reset = reset;
assign left_5_6_in = left_5_5_out;
assign left_6_5_write_en = _guard1798;
assign left_6_5_clk = clk;
assign left_6_5_reset = reset;
assign left_6_5_in = left_6_4_out;
assign top_6_6_write_en = _guard1804;
assign top_6_6_clk = clk;
assign top_6_6_reset = reset;
assign top_6_6_in = top_5_6_out;
assign l0_idx_write_en = _guard1812;
assign l0_idx_clk = clk;
assign l0_idx_reset = reset;
assign l0_idx_in =
  _guard1813 ? 4'd0 :
  _guard1816 ? l0_add_out :
  'x;
assign idx_between_depth_plus_16_depth_plus_17_comb_left = index_ge_depth_plus_16_out;
assign idx_between_depth_plus_16_depth_plus_17_comb_right = index_lt_depth_plus_17_out;
assign index_ge_depth_plus_12_left = idx_add_out;
assign index_ge_depth_plus_12_right = depth_plus_12_out;
assign index_ge_depth_plus_17_left = idx_add_out;
assign index_ge_depth_plus_17_right = depth_plus_17_out;
assign idx_between_16_depth_plus_16_reg_write_en = _guard1825;
assign idx_between_16_depth_plus_16_reg_clk = clk;
assign idx_between_16_depth_plus_16_reg_reset = reset;
assign idx_between_16_depth_plus_16_reg_in =
  _guard1826 ? 1'd0 :
  _guard1827 ? idx_between_16_depth_plus_16_comb_out :
  'x;
assign index_lt_depth_plus_19_left = idx_add_out;
assign index_lt_depth_plus_19_right = depth_plus_19_out;
assign idx_between_3_min_depth_4_plus_3_comb_left = index_ge_3_out;
assign idx_between_3_min_depth_4_plus_3_comb_right = index_lt_min_depth_4_plus_3_out;
assign idx_between_12_min_depth_4_plus_12_comb_left = index_ge_12_out;
assign idx_between_12_min_depth_4_plus_12_comb_right = index_lt_min_depth_4_plus_12_out;
assign idx_between_depth_plus_14_depth_plus_15_comb_left = index_ge_depth_plus_14_out;
assign idx_between_depth_plus_14_depth_plus_15_comb_right = index_lt_depth_plus_15_out;
assign index_ge_depth_plus_9_left = idx_add_out;
assign index_ge_depth_plus_9_right = depth_plus_9_out;
assign idx_between_8_min_depth_4_plus_8_comb_left = index_ge_8_out;
assign idx_between_8_min_depth_4_plus_8_comb_right = index_lt_min_depth_4_plus_8_out;
assign idx_between_13_depth_plus_13_reg_write_en = _guard1842;
assign idx_between_13_depth_plus_13_reg_clk = clk;
assign idx_between_13_depth_plus_13_reg_reset = reset;
assign idx_between_13_depth_plus_13_reg_in =
  _guard1843 ? 1'd0 :
  _guard1844 ? idx_between_13_depth_plus_13_comb_out :
  'x;
assign idx_between_15_depth_plus_15_reg_write_en = _guard1847;
assign idx_between_15_depth_plus_15_reg_clk = clk;
assign idx_between_15_depth_plus_15_reg_reset = reset;
assign idx_between_15_depth_plus_15_reg_in =
  _guard1848 ? idx_between_15_depth_plus_15_comb_out :
  _guard1849 ? 1'd0 :
  'x;
assign idx_between_14_min_depth_4_plus_14_reg_write_en = _guard1852;
assign idx_between_14_min_depth_4_plus_14_reg_clk = clk;
assign idx_between_14_min_depth_4_plus_14_reg_reset = reset;
assign idx_between_14_min_depth_4_plus_14_reg_in =
  _guard1853 ? 1'd0 :
  _guard1854 ? idx_between_14_min_depth_4_plus_14_comb_out :
  'x;
assign idx_between_1_min_depth_4_plus_1_reg_write_en = _guard1857;
assign idx_between_1_min_depth_4_plus_1_reg_clk = clk;
assign idx_between_1_min_depth_4_plus_1_reg_reset = reset;
assign idx_between_1_min_depth_4_plus_1_reg_in =
  _guard1858 ? 1'd0 :
  _guard1859 ? idx_between_1_min_depth_4_plus_1_comb_out :
  'x;
assign idx_between_15_min_depth_4_plus_15_reg_write_en = _guard1862;
assign idx_between_15_min_depth_4_plus_15_reg_clk = clk;
assign idx_between_15_min_depth_4_plus_15_reg_reset = reset;
assign idx_between_15_min_depth_4_plus_15_reg_in =
  _guard1863 ? idx_between_15_min_depth_4_plus_15_comb_out :
  _guard1864 ? 1'd0 :
  'x;
assign idx_between_15_min_depth_4_plus_15_comb_left = index_ge_15_out;
assign idx_between_15_min_depth_4_plus_15_comb_right = index_lt_min_depth_4_plus_15_out;
assign cond11_write_en = _guard1867;
assign cond11_clk = clk;
assign cond11_reset = reset;
assign cond11_in =
  _guard1868 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond15_write_en = _guard1869;
assign cond15_clk = clk;
assign cond15_reset = reset;
assign cond15_in =
  _guard1870 ? idx_between_4_min_depth_4_plus_4_reg_out :
  1'd0;
assign cond_wire27_in =
  _guard1873 ? cond27_out :
  _guard1874 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond43_write_en = _guard1875;
assign cond43_clk = clk;
assign cond43_reset = reset;
assign cond43_in =
  _guard1876 ? idx_between_depth_plus_6_depth_plus_7_reg_out :
  1'd0;
assign cond_wire43_in =
  _guard1877 ? idx_between_depth_plus_6_depth_plus_7_reg_out :
  _guard1880 ? cond43_out :
  1'd0;
assign cond_wire44_in =
  _guard1883 ? cond44_out :
  _guard1884 ? idx_between_3_min_depth_4_plus_3_reg_out :
  1'd0;
assign cond62_write_en = _guard1885;
assign cond62_clk = clk;
assign cond62_reset = reset;
assign cond62_in =
  _guard1886 ? idx_between_11_depth_plus_11_reg_out :
  1'd0;
assign cond_wire63_in =
  _guard1889 ? cond63_out :
  _guard1890 ? idx_between_depth_plus_11_depth_plus_12_reg_out :
  1'd0;
assign cond_wire67_in =
  _guard1893 ? cond67_out :
  _guard1894 ? idx_between_depth_plus_12_depth_plus_13_reg_out :
  1'd0;
assign cond73_write_en = _guard1895;
assign cond73_clk = clk;
assign cond73_reset = reset;
assign cond73_in =
  _guard1896 ? idx_between_3_min_depth_4_plus_3_reg_out :
  1'd0;
assign cond_wire77_in =
  _guard1899 ? cond77_out :
  _guard1900 ? idx_between_4_min_depth_4_plus_4_reg_out :
  1'd0;
assign cond103_write_en = _guard1901;
assign cond103_clk = clk;
assign cond103_reset = reset;
assign cond103_in =
  _guard1902 ? idx_between_14_depth_plus_14_reg_out :
  1'd0;
assign cond114_write_en = _guard1903;
assign cond114_clk = clk;
assign cond114_reset = reset;
assign cond114_in =
  _guard1904 ? idx_between_6_min_depth_4_plus_6_reg_out :
  1'd0;
assign cond118_write_en = _guard1905;
assign cond118_clk = clk;
assign cond118_reset = reset;
assign cond118_in =
  _guard1906 ? idx_between_7_min_depth_4_plus_7_reg_out :
  1'd0;
assign cond121_write_en = _guard1907;
assign cond121_clk = clk;
assign cond121_reset = reset;
assign cond121_in =
  _guard1908 ? idx_between_depth_plus_11_depth_plus_12_reg_out :
  1'd0;
assign cond123_write_en = _guard1909;
assign cond123_clk = clk;
assign cond123_reset = reset;
assign cond123_in =
  _guard1910 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire126_in =
  _guard1911 ? idx_between_9_min_depth_4_plus_9_reg_out :
  _guard1914 ? cond126_out :
  1'd0;
assign cond_wire154_in =
  _guard1917 ? cond154_out :
  _guard1918 ? idx_between_depth_plus_12_depth_plus_13_reg_out :
  1'd0;
assign cond_wire195_in =
  _guard1921 ? cond195_out :
  _guard1922 ? idx_between_depth_plus_15_depth_plus_16_reg_out :
  1'd0;
assign cond206_write_en = _guard1923;
assign cond206_clk = clk;
assign cond206_reset = reset;
assign cond206_in =
  _guard1924 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond216_write_en = _guard1925;
assign cond216_clk = clk;
assign cond216_reset = reset;
assign cond216_in =
  _guard1926 ? idx_between_depth_plus_13_depth_plus_14_reg_out :
  1'd0;
assign cond_wire218_in =
  _guard1927 ? idx_between_10_depth_plus_10_reg_out :
  _guard1930 ? cond218_out :
  1'd0;
assign cond_wire238_in =
  _guard1931 ? idx_between_8_min_depth_4_plus_8_reg_out :
  _guard1934 ? cond238_out :
  1'd0;
assign cond240_write_en = _guard1935;
assign cond240_clk = clk;
assign cond240_reset = reset;
assign cond240_in =
  _guard1936 ? idx_between_12_depth_plus_12_reg_out :
  1'd0;
assign cond251_write_en = _guard1937;
assign cond251_clk = clk;
assign cond251_reset = reset;
assign cond251_in =
  _guard1938 ? idx_between_11_depth_plus_11_reg_out :
  1'd0;
assign cond264_write_en = _guard1939;
assign cond264_clk = clk;
assign cond264_reset = reset;
assign cond264_in =
  _guard1940 ? idx_between_18_depth_plus_18_reg_out :
  1'd0;
assign cond_wire265_in =
  _guard1943 ? cond265_out :
  _guard1944 ? idx_between_depth_plus_18_depth_plus_19_reg_out :
  1'd0;
assign pe_0_1_mul_ready =
  _guard1947 ? 1'd1 :
  _guard1950 ? 1'd0 :
  1'd0;
assign pe_0_1_clk = clk;
assign pe_0_1_top =
  _guard1963 ? top_0_1_out :
  32'd0;
assign pe_0_1_left =
  _guard1976 ? left_0_1_out :
  32'd0;
assign pe_0_1_reset = reset;
assign pe_0_1_go = _guard1989;
assign left_0_6_write_en = _guard1992;
assign left_0_6_clk = clk;
assign left_0_6_reset = reset;
assign left_0_6_in = left_0_5_out;
assign pe_0_7_mul_ready =
  _guard1998 ? 1'd1 :
  _guard2001 ? 1'd0 :
  1'd0;
assign pe_0_7_clk = clk;
assign pe_0_7_top =
  _guard2014 ? top_0_7_out :
  32'd0;
assign pe_0_7_left =
  _guard2027 ? left_0_7_out :
  32'd0;
assign pe_0_7_reset = reset;
assign pe_0_7_go = _guard2040;
assign left_1_2_write_en = _guard2043;
assign left_1_2_clk = clk;
assign left_1_2_reset = reset;
assign left_1_2_in = left_1_1_out;
assign left_2_2_write_en = _guard2049;
assign left_2_2_clk = clk;
assign left_2_2_reset = reset;
assign left_2_2_in = left_2_1_out;
assign top_2_5_write_en = _guard2055;
assign top_2_5_clk = clk;
assign top_2_5_reset = reset;
assign top_2_5_in = top_1_5_out;
assign pe_2_7_mul_ready =
  _guard2061 ? 1'd1 :
  _guard2064 ? 1'd0 :
  1'd0;
assign pe_2_7_clk = clk;
assign pe_2_7_top =
  _guard2077 ? top_2_7_out :
  32'd0;
assign pe_2_7_left =
  _guard2090 ? left_2_7_out :
  32'd0;
assign pe_2_7_reset = reset;
assign pe_2_7_go = _guard2103;
assign left_2_7_write_en = _guard2106;
assign left_2_7_clk = clk;
assign left_2_7_reset = reset;
assign left_2_7_in = left_2_6_out;
assign pe_4_5_mul_ready =
  _guard2112 ? 1'd1 :
  _guard2115 ? 1'd0 :
  1'd0;
assign pe_4_5_clk = clk;
assign pe_4_5_top =
  _guard2128 ? top_4_5_out :
  32'd0;
assign pe_4_5_left =
  _guard2141 ? left_4_5_out :
  32'd0;
assign pe_4_5_reset = reset;
assign pe_4_5_go = _guard2154;
assign left_4_5_write_en = _guard2157;
assign left_4_5_clk = clk;
assign left_4_5_reset = reset;
assign left_4_5_in = left_4_4_out;
assign top_5_0_write_en = _guard2163;
assign top_5_0_clk = clk;
assign top_5_0_reset = reset;
assign top_5_0_in = top_4_0_out;
assign top_5_3_write_en = _guard2169;
assign top_5_3_clk = clk;
assign top_5_3_reset = reset;
assign top_5_3_in = top_4_3_out;
assign l3_add_left = 4'd1;
assign l3_add_right = l3_idx_out;
assign idx_between_11_depth_plus_11_comb_left = index_ge_11_out;
assign idx_between_11_depth_plus_11_comb_right = index_lt_depth_plus_11_out;
assign index_lt_min_depth_4_plus_7_left = idx_add_out;
assign index_lt_min_depth_4_plus_7_right = min_depth_4_plus_7_out;
assign index_ge_3_left = idx_add_out;
assign index_ge_3_right = 32'd3;
assign idx_between_12_depth_plus_12_reg_write_en = _guard2187;
assign idx_between_12_depth_plus_12_reg_clk = clk;
assign idx_between_12_depth_plus_12_reg_reset = reset;
assign idx_between_12_depth_plus_12_reg_in =
  _guard2188 ? idx_between_12_depth_plus_12_comb_out :
  _guard2189 ? 1'd0 :
  'x;
assign index_ge_12_left = idx_add_out;
assign index_ge_12_right = 32'd12;
assign idx_between_13_min_depth_4_plus_13_comb_left = index_ge_13_out;
assign idx_between_13_min_depth_4_plus_13_comb_right = index_lt_min_depth_4_plus_13_out;
assign index_lt_depth_plus_4_left = idx_add_out;
assign index_lt_depth_plus_4_right = depth_plus_4_out;
assign idx_between_5_depth_plus_5_comb_left = index_ge_5_out;
assign idx_between_5_depth_plus_5_comb_right = index_lt_depth_plus_5_out;
assign idx_between_19_depth_plus_19_reg_write_en = _guard2200;
assign idx_between_19_depth_plus_19_reg_clk = clk;
assign idx_between_19_depth_plus_19_reg_reset = reset;
assign idx_between_19_depth_plus_19_reg_in =
  _guard2201 ? 1'd0 :
  _guard2202 ? idx_between_19_depth_plus_19_comb_out :
  'x;
assign cond_write_en = _guard2203;
assign cond_clk = clk;
assign cond_reset = reset;
assign cond_in =
  _guard2204 ? idx_between_0_depth_plus_0_reg_out :
  1'd0;
assign cond_wire26_in =
  _guard2205 ? idx_between_6_depth_plus_6_reg_out :
  _guard2208 ? cond26_out :
  1'd0;
assign cond35_write_en = _guard2209;
assign cond35_clk = clk;
assign cond35_reset = reset;
assign cond35_in =
  _guard2210 ? idx_between_8_min_depth_4_plus_8_reg_out :
  1'd0;
assign cond_wire35_in =
  _guard2211 ? idx_between_8_min_depth_4_plus_8_reg_out :
  _guard2214 ? cond35_out :
  1'd0;
assign cond_wire50_in =
  _guard2217 ? cond50_out :
  _guard2218 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire56_in =
  _guard2219 ? idx_between_6_min_depth_4_plus_6_reg_out :
  _guard2222 ? cond56_out :
  1'd0;
assign cond60_write_en = _guard2223;
assign cond60_clk = clk;
assign cond60_reset = reset;
assign cond60_in =
  _guard2224 ? idx_between_7_min_depth_4_plus_7_reg_out :
  1'd0;
assign cond69_write_en = _guard2225;
assign cond69_clk = clk;
assign cond69_reset = reset;
assign cond69_in =
  _guard2226 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond72_write_en = _guard2227;
assign cond72_clk = clk;
assign cond72_reset = reset;
assign cond72_in =
  _guard2228 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond76_write_en = _guard2229;
assign cond76_clk = clk;
assign cond76_reset = reset;
assign cond76_in =
  _guard2230 ? idx_between_depth_plus_7_depth_plus_8_reg_out :
  1'd0;
assign cond_wire85_in =
  _guard2231 ? idx_between_6_min_depth_4_plus_6_reg_out :
  _guard2234 ? cond85_out :
  1'd0;
assign cond92_write_en = _guard2235;
assign cond92_clk = clk;
assign cond92_reset = reset;
assign cond92_in =
  _guard2236 ? idx_between_depth_plus_11_depth_plus_12_reg_out :
  1'd0;
assign cond_wire116_in =
  _guard2239 ? cond116_out :
  _guard2240 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond_wire149_in =
  _guard2241 ? idx_between_11_depth_plus_11_reg_out :
  _guard2244 ? cond149_out :
  1'd0;
assign cond_wire163_in =
  _guard2245 ? idx_between_11_min_depth_4_plus_11_reg_out :
  _guard2248 ? cond163_out :
  1'd0;
assign cond_wire182_in =
  _guard2249 ? idx_between_12_depth_plus_12_reg_out :
  _guard2252 ? cond182_out :
  1'd0;
assign cond189_write_en = _guard2253;
assign cond189_clk = clk;
assign cond189_reset = reset;
assign cond189_in =
  _guard2254 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond_wire192_in =
  _guard2255 ? idx_between_11_min_depth_4_plus_11_reg_out :
  _guard2258 ? cond192_out :
  1'd0;
assign cond_wire200_in =
  _guard2259 ? idx_between_13_min_depth_4_plus_13_reg_out :
  _guard2262 ? cond200_out :
  1'd0;
assign cond_wire205_in =
  _guard2263 ? idx_between_7_min_depth_4_plus_7_reg_out :
  _guard2266 ? cond205_out :
  1'd0;
assign cond226_write_en = _guard2267;
assign cond226_clk = clk;
assign cond226_reset = reset;
assign cond226_in =
  _guard2268 ? idx_between_12_depth_plus_12_reg_out :
  1'd0;
assign cond233_write_en = _guard2269;
assign cond233_clk = clk;
assign cond233_reset = reset;
assign cond233_in =
  _guard2270 ? idx_between_14_min_depth_4_plus_14_reg_out :
  1'd0;
assign cond241_write_en = _guard2271;
assign cond241_clk = clk;
assign cond241_reset = reset;
assign cond241_in =
  _guard2272 ? idx_between_depth_plus_12_depth_plus_13_reg_out :
  1'd0;
assign cond_wire243_in =
  _guard2273 ? idx_between_9_depth_plus_9_reg_out :
  _guard2276 ? cond243_out :
  1'd0;
assign cond_wire245_in =
  _guard2279 ? cond245_out :
  _guard2280 ? idx_between_depth_plus_13_depth_plus_14_reg_out :
  1'd0;
assign cond248_write_en = _guard2281;
assign cond248_clk = clk;
assign cond248_reset = reset;
assign cond248_in =
  _guard2282 ? idx_between_14_depth_plus_14_reg_out :
  1'd0;
assign cond257_write_en = _guard2283;
assign cond257_clk = clk;
assign cond257_reset = reset;
assign cond257_in =
  _guard2284 ? idx_between_depth_plus_16_depth_plus_17_reg_out :
  1'd0;
assign cond_wire263_in =
  _guard2287 ? cond263_out :
  _guard2288 ? idx_between_14_depth_plus_14_reg_out :
  1'd0;
assign cond266_write_en = _guard2289;
assign cond266_clk = clk;
assign cond266_reset = reset;
assign cond266_in =
  _guard2290 ? idx_between_15_min_depth_4_plus_15_reg_out :
  1'd0;
assign depth_plus_18_left = depth;
assign depth_plus_18_right = 32'd18;
assign depth_plus_5_left = depth;
assign depth_plus_5_right = 32'd5;
assign pe_1_0_mul_ready =
  _guard2297 ? 1'd1 :
  _guard2300 ? 1'd0 :
  1'd0;
assign pe_1_0_clk = clk;
assign pe_1_0_top =
  _guard2313 ? top_1_0_out :
  32'd0;
assign pe_1_0_left =
  _guard2326 ? left_1_0_out :
  32'd0;
assign pe_1_0_reset = reset;
assign pe_1_0_go = _guard2339;
assign left_1_0_write_en = _guard2342;
assign left_1_0_clk = clk;
assign left_1_0_reset = reset;
assign left_1_0_in = l1_read_data;
assign left_1_1_write_en = _guard2348;
assign left_1_1_clk = clk;
assign left_1_1_reset = reset;
assign left_1_1_in = left_1_0_out;
assign top_1_2_write_en = _guard2354;
assign top_1_2_clk = clk;
assign top_1_2_reset = reset;
assign top_1_2_in = top_0_2_out;
assign left_2_0_write_en = _guard2360;
assign left_2_0_clk = clk;
assign left_2_0_reset = reset;
assign left_2_0_in = l2_read_data;
assign left_3_1_write_en = _guard2366;
assign left_3_1_clk = clk;
assign left_3_1_reset = reset;
assign left_3_1_in = left_3_0_out;
assign pe_3_2_mul_ready =
  _guard2372 ? 1'd1 :
  _guard2375 ? 1'd0 :
  1'd0;
assign pe_3_2_clk = clk;
assign pe_3_2_top =
  _guard2388 ? top_3_2_out :
  32'd0;
assign pe_3_2_left =
  _guard2401 ? left_3_2_out :
  32'd0;
assign pe_3_2_reset = reset;
assign pe_3_2_go = _guard2414;
assign pe_3_5_mul_ready =
  _guard2417 ? 1'd1 :
  _guard2420 ? 1'd0 :
  1'd0;
assign pe_3_5_clk = clk;
assign pe_3_5_top =
  _guard2433 ? top_3_5_out :
  32'd0;
assign pe_3_5_left =
  _guard2446 ? left_3_5_out :
  32'd0;
assign pe_3_5_reset = reset;
assign pe_3_5_go = _guard2459;
assign pe_3_6_mul_ready =
  _guard2462 ? 1'd1 :
  _guard2465 ? 1'd0 :
  1'd0;
assign pe_3_6_clk = clk;
assign pe_3_6_top =
  _guard2478 ? top_3_6_out :
  32'd0;
assign pe_3_6_left =
  _guard2491 ? left_3_6_out :
  32'd0;
assign pe_3_6_reset = reset;
assign pe_3_6_go = _guard2504;
assign left_3_7_write_en = _guard2507;
assign left_3_7_clk = clk;
assign left_3_7_reset = reset;
assign left_3_7_in = left_3_6_out;
assign top_4_5_write_en = _guard2513;
assign top_4_5_clk = clk;
assign top_4_5_reset = reset;
assign top_4_5_in = top_3_5_out;
assign pe_5_4_mul_ready =
  _guard2519 ? 1'd1 :
  _guard2522 ? 1'd0 :
  1'd0;
assign pe_5_4_clk = clk;
assign pe_5_4_top =
  _guard2535 ? top_5_4_out :
  32'd0;
assign pe_5_4_left =
  _guard2548 ? left_5_4_out :
  32'd0;
assign pe_5_4_reset = reset;
assign pe_5_4_go = _guard2561;
assign top_7_2_write_en = _guard2564;
assign top_7_2_clk = clk;
assign top_7_2_reset = reset;
assign top_7_2_in = top_6_2_out;
assign pe_7_4_mul_ready =
  _guard2570 ? 1'd1 :
  _guard2573 ? 1'd0 :
  1'd0;
assign pe_7_4_clk = clk;
assign pe_7_4_top =
  _guard2586 ? top_7_4_out :
  32'd0;
assign pe_7_4_left =
  _guard2599 ? left_7_4_out :
  32'd0;
assign pe_7_4_reset = reset;
assign pe_7_4_go = _guard2612;
assign t1_idx_write_en = _guard2617;
assign t1_idx_clk = clk;
assign t1_idx_reset = reset;
assign t1_idx_in =
  _guard2618 ? 4'd0 :
  _guard2621 ? t1_add_out :
  'x;
assign t7_idx_write_en = _guard2626;
assign t7_idx_clk = clk;
assign t7_idx_reset = reset;
assign t7_idx_in =
  _guard2627 ? 4'd0 :
  _guard2630 ? t7_add_out :
  'x;
assign idx_between_depth_plus_8_depth_plus_9_comb_left = index_ge_depth_plus_8_out;
assign idx_between_depth_plus_8_depth_plus_9_comb_right = index_lt_depth_plus_9_out;
assign index_lt_min_depth_4_plus_11_left = idx_add_out;
assign index_lt_min_depth_4_plus_11_right = min_depth_4_plus_11_out;
assign idx_between_7_min_depth_4_plus_7_comb_left = index_ge_7_out;
assign idx_between_7_min_depth_4_plus_7_comb_right = index_lt_min_depth_4_plus_7_out;
assign idx_between_12_depth_plus_12_comb_left = index_ge_12_out;
assign idx_between_12_depth_plus_12_comb_right = index_lt_depth_plus_12_out;
assign idx_between_depth_plus_9_depth_plus_10_reg_write_en = _guard2641;
assign idx_between_depth_plus_9_depth_plus_10_reg_clk = clk;
assign idx_between_depth_plus_9_depth_plus_10_reg_reset = reset;
assign idx_between_depth_plus_9_depth_plus_10_reg_in =
  _guard2642 ? 1'd0 :
  _guard2643 ? idx_between_depth_plus_9_depth_plus_10_comb_out :
  'x;
assign index_lt_depth_plus_10_left = idx_add_out;
assign index_lt_depth_plus_10_right = depth_plus_10_out;
assign idx_between_depth_plus_6_depth_plus_7_comb_left = index_ge_depth_plus_6_out;
assign idx_between_depth_plus_6_depth_plus_7_comb_right = index_lt_depth_plus_7_out;
assign index_ge_18_left = idx_add_out;
assign index_ge_18_right = 32'd18;
assign idx_between_15_depth_plus_15_comb_left = index_ge_15_out;
assign idx_between_15_depth_plus_15_comb_right = index_lt_depth_plus_15_out;
assign cond18_write_en = _guard2652;
assign cond18_clk = clk;
assign cond18_reset = reset;
assign cond18_in =
  _guard2653 ? idx_between_depth_plus_8_depth_plus_9_reg_out :
  1'd0;
assign cond_wire24_in =
  _guard2656 ? cond24_out :
  _guard2657 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond_wire31_in =
  _guard2658 ? idx_between_7_depth_plus_7_reg_out :
  _guard2661 ? cond31_out :
  1'd0;
assign cond_wire46_in =
  _guard2662 ? idx_between_7_depth_plus_7_reg_out :
  _guard2665 ? cond46_out :
  1'd0;
assign cond_wire48_in =
  _guard2668 ? cond48_out :
  _guard2669 ? idx_between_4_min_depth_4_plus_4_reg_out :
  1'd0;
assign cond_wire72_in =
  _guard2672 ? cond72_out :
  _guard2673 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond_wire76_in =
  _guard2676 ? cond76_out :
  _guard2677 ? idx_between_depth_plus_7_depth_plus_8_reg_out :
  1'd0;
assign cond_wire100_in =
  _guard2680 ? cond100_out :
  _guard2681 ? idx_between_depth_plus_13_depth_plus_14_reg_out :
  1'd0;
assign cond105_write_en = _guard2682;
assign cond105_clk = clk;
assign cond105_reset = reset;
assign cond105_in =
  _guard2683 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond_wire134_in =
  _guard2684 ? idx_between_11_min_depth_4_plus_11_reg_out :
  _guard2687 ? cond134_out :
  1'd0;
assign cond146_write_en = _guard2688;
assign cond146_clk = clk;
assign cond146_reset = reset;
assign cond146_in =
  _guard2689 ? idx_between_depth_plus_10_depth_plus_11_reg_out :
  1'd0;
assign cond_wire146_in =
  _guard2692 ? cond146_out :
  _guard2693 ? idx_between_depth_plus_10_depth_plus_11_reg_out :
  1'd0;
assign cond151_write_en = _guard2694;
assign cond151_clk = clk;
assign cond151_reset = reset;
assign cond151_in =
  _guard2695 ? idx_between_8_min_depth_4_plus_8_reg_out :
  1'd0;
assign cond_wire157_in =
  _guard2696 ? idx_between_13_depth_plus_13_reg_out :
  _guard2699 ? cond157_out :
  1'd0;
assign cond_wire167_in =
  _guard2702 ? cond167_out :
  _guard2703 ? idx_between_12_min_depth_4_plus_12_reg_out :
  1'd0;
assign cond_wire174_in =
  _guard2706 ? cond174_out :
  _guard2707 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond177_write_en = _guard2708;
assign cond177_clk = clk;
assign cond177_reset = reset;
assign cond177_in =
  _guard2709 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond178_write_en = _guard2710;
assign cond178_clk = clk;
assign cond178_reset = reset;
assign cond178_in =
  _guard2711 ? idx_between_11_depth_plus_11_reg_out :
  1'd0;
assign cond_wire191_in =
  _guard2714 ? cond191_out :
  _guard2715 ? idx_between_depth_plus_14_depth_plus_15_reg_out :
  1'd0;
assign cond_wire198_in =
  _guard2716 ? idx_between_16_depth_plus_16_reg_out :
  _guard2719 ? cond198_out :
  1'd0;
assign cond204_write_en = _guard2720;
assign cond204_clk = clk;
assign cond204_reset = reset;
assign cond204_in =
  _guard2721 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond215_write_en = _guard2722;
assign cond215_clk = clk;
assign cond215_reset = reset;
assign cond215_in =
  _guard2723 ? idx_between_13_depth_plus_13_reg_out :
  1'd0;
assign cond_wire216_in =
  _guard2726 ? cond216_out :
  _guard2727 ? idx_between_depth_plus_13_depth_plus_14_reg_out :
  1'd0;
assign cond_wire228_in =
  _guard2730 ? cond228_out :
  _guard2731 ? idx_between_depth_plus_16_depth_plus_17_reg_out :
  1'd0;
assign cond231_write_en = _guard2732;
assign cond231_clk = clk;
assign cond231_reset = reset;
assign cond231_in =
  _guard2733 ? idx_between_17_depth_plus_17_reg_out :
  1'd0;
assign cond_wire231_in =
  _guard2736 ? cond231_out :
  _guard2737 ? idx_between_17_depth_plus_17_reg_out :
  1'd0;
assign cond237_write_en = _guard2738;
assign cond237_clk = clk;
assign cond237_reset = reset;
assign cond237_in =
  _guard2739 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign depth_plus_12_left = depth;
assign depth_plus_12_right = 32'd12;
assign min_depth_4_plus_2_left = min_depth_4_out;
assign min_depth_4_plus_2_right = 32'd2;
assign min_depth_4_plus_14_left = min_depth_4_out;
assign min_depth_4_plus_14_right = 32'd14;
assign depth_plus_1_left = depth;
assign depth_plus_1_right = 32'd1;
assign min_depth_4_plus_15_left = min_depth_4_out;
assign min_depth_4_plus_15_right = 32'd15;
assign left_0_0_write_en = _guard2752;
assign left_0_0_clk = clk;
assign left_0_0_reset = reset;
assign left_0_0_in = l0_read_data;
assign pe_0_3_mul_ready =
  _guard2758 ? 1'd1 :
  _guard2761 ? 1'd0 :
  1'd0;
assign pe_0_3_clk = clk;
assign pe_0_3_top =
  _guard2774 ? top_0_3_out :
  32'd0;
assign pe_0_3_left =
  _guard2787 ? left_0_3_out :
  32'd0;
assign pe_0_3_reset = reset;
assign pe_0_3_go = _guard2800;
assign pe_0_5_mul_ready =
  _guard2803 ? 1'd1 :
  _guard2806 ? 1'd0 :
  1'd0;
assign pe_0_5_clk = clk;
assign pe_0_5_top =
  _guard2819 ? top_0_5_out :
  32'd0;
assign pe_0_5_left =
  _guard2832 ? left_0_5_out :
  32'd0;
assign pe_0_5_reset = reset;
assign pe_0_5_go = _guard2845;
assign top_1_3_write_en = _guard2848;
assign top_1_3_clk = clk;
assign top_1_3_reset = reset;
assign top_1_3_in = top_0_3_out;
assign top_1_4_write_en = _guard2854;
assign top_1_4_clk = clk;
assign top_1_4_reset = reset;
assign top_1_4_in = top_0_4_out;
assign left_2_3_write_en = _guard2860;
assign left_2_3_clk = clk;
assign left_2_3_reset = reset;
assign left_2_3_in = left_2_2_out;
assign pe_2_4_mul_ready =
  _guard2866 ? 1'd1 :
  _guard2869 ? 1'd0 :
  1'd0;
assign pe_2_4_clk = clk;
assign pe_2_4_top =
  _guard2882 ? top_2_4_out :
  32'd0;
assign pe_2_4_left =
  _guard2895 ? left_2_4_out :
  32'd0;
assign pe_2_4_reset = reset;
assign pe_2_4_go = _guard2908;
assign top_2_6_write_en = _guard2911;
assign top_2_6_clk = clk;
assign top_2_6_reset = reset;
assign top_2_6_in = top_1_6_out;
assign pe_3_0_mul_ready =
  _guard2917 ? 1'd1 :
  _guard2920 ? 1'd0 :
  1'd0;
assign pe_3_0_clk = clk;
assign pe_3_0_top =
  _guard2933 ? top_3_0_out :
  32'd0;
assign pe_3_0_left =
  _guard2946 ? left_3_0_out :
  32'd0;
assign pe_3_0_reset = reset;
assign pe_3_0_go = _guard2959;
assign top_3_2_write_en = _guard2962;
assign top_3_2_clk = clk;
assign top_3_2_reset = reset;
assign top_3_2_in = top_2_2_out;
assign top_4_0_write_en = _guard2968;
assign top_4_0_clk = clk;
assign top_4_0_reset = reset;
assign top_4_0_in = top_3_0_out;
assign left_4_6_write_en = _guard2974;
assign left_4_6_clk = clk;
assign left_4_6_reset = reset;
assign left_4_6_in = left_4_5_out;
assign left_4_7_write_en = _guard2980;
assign left_4_7_clk = clk;
assign left_4_7_reset = reset;
assign left_4_7_in = left_4_6_out;
assign pe_5_1_mul_ready =
  _guard2986 ? 1'd1 :
  _guard2989 ? 1'd0 :
  1'd0;
assign pe_5_1_clk = clk;
assign pe_5_1_top =
  _guard3002 ? top_5_1_out :
  32'd0;
assign pe_5_1_left =
  _guard3015 ? left_5_1_out :
  32'd0;
assign pe_5_1_reset = reset;
assign pe_5_1_go = _guard3028;
assign pe_5_7_mul_ready =
  _guard3031 ? 1'd1 :
  _guard3034 ? 1'd0 :
  1'd0;
assign pe_5_7_clk = clk;
assign pe_5_7_top =
  _guard3047 ? top_5_7_out :
  32'd0;
assign pe_5_7_left =
  _guard3060 ? left_5_7_out :
  32'd0;
assign pe_5_7_reset = reset;
assign pe_5_7_go = _guard3073;
assign pe_6_0_mul_ready =
  _guard3076 ? 1'd1 :
  _guard3079 ? 1'd0 :
  1'd0;
assign pe_6_0_clk = clk;
assign pe_6_0_top =
  _guard3092 ? top_6_0_out :
  32'd0;
assign pe_6_0_left =
  _guard3105 ? left_6_0_out :
  32'd0;
assign pe_6_0_reset = reset;
assign pe_6_0_go = _guard3118;
assign top_6_0_write_en = _guard3121;
assign top_6_0_clk = clk;
assign top_6_0_reset = reset;
assign top_6_0_in = top_5_0_out;
assign pe_6_1_mul_ready =
  _guard3127 ? 1'd1 :
  _guard3130 ? 1'd0 :
  1'd0;
assign pe_6_1_clk = clk;
assign pe_6_1_top =
  _guard3143 ? top_6_1_out :
  32'd0;
assign pe_6_1_left =
  _guard3156 ? left_6_1_out :
  32'd0;
assign pe_6_1_reset = reset;
assign pe_6_1_go = _guard3169;
assign left_7_5_write_en = _guard3172;
assign left_7_5_clk = clk;
assign left_7_5_reset = reset;
assign left_7_5_in = left_7_4_out;
assign idx_between_7_min_depth_4_plus_7_reg_write_en = _guard3178;
assign idx_between_7_min_depth_4_plus_7_reg_clk = clk;
assign idx_between_7_min_depth_4_plus_7_reg_reset = reset;
assign idx_between_7_min_depth_4_plus_7_reg_in =
  _guard3179 ? idx_between_7_min_depth_4_plus_7_comb_out :
  _guard3180 ? 1'd0 :
  'x;
assign idx_between_12_min_depth_4_plus_12_reg_write_en = _guard3183;
assign idx_between_12_min_depth_4_plus_12_reg_clk = clk;
assign idx_between_12_min_depth_4_plus_12_reg_reset = reset;
assign idx_between_12_min_depth_4_plus_12_reg_in =
  _guard3184 ? idx_between_12_min_depth_4_plus_12_comb_out :
  _guard3185 ? 1'd0 :
  'x;
assign idx_between_depth_plus_5_depth_plus_6_reg_write_en = _guard3188;
assign idx_between_depth_plus_5_depth_plus_6_reg_clk = clk;
assign idx_between_depth_plus_5_depth_plus_6_reg_reset = reset;
assign idx_between_depth_plus_5_depth_plus_6_reg_in =
  _guard3189 ? 1'd0 :
  _guard3190 ? idx_between_depth_plus_5_depth_plus_6_comb_out :
  'x;
assign index_lt_depth_plus_8_left = idx_add_out;
assign index_lt_depth_plus_8_right = depth_plus_8_out;
assign idx_between_6_min_depth_4_plus_6_comb_left = index_ge_6_out;
assign idx_between_6_min_depth_4_plus_6_comb_right = index_lt_min_depth_4_plus_6_out;
assign cond_wire18_in =
  _guard3195 ? idx_between_depth_plus_8_depth_plus_9_reg_out :
  _guard3198 ? cond18_out :
  1'd0;
assign cond19_write_en = _guard3199;
assign cond19_clk = clk;
assign cond19_reset = reset;
assign cond19_in =
  _guard3200 ? idx_between_4_depth_plus_4_reg_out :
  1'd0;
assign cond_wire29_in =
  _guard3203 ? cond29_out :
  _guard3204 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond34_write_en = _guard3205;
assign cond34_clk = clk;
assign cond34_reset = reset;
assign cond34_in =
  _guard3206 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond40_write_en = _guard3207;
assign cond40_clk = clk;
assign cond40_reset = reset;
assign cond40_in =
  _guard3208 ? idx_between_2_min_depth_4_plus_2_reg_out :
  1'd0;
assign cond57_write_en = _guard3209;
assign cond57_clk = clk;
assign cond57_reset = reset;
assign cond57_in =
  _guard3210 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire59_in =
  _guard3211 ? idx_between_depth_plus_10_depth_plus_11_reg_out :
  _guard3214 ? cond59_out :
  1'd0;
assign cond_wire61_in =
  _guard3215 ? idx_between_7_depth_plus_7_reg_out :
  _guard3218 ? cond61_out :
  1'd0;
assign cond74_write_en = _guard3219;
assign cond74_clk = clk;
assign cond74_reset = reset;
assign cond74_in =
  _guard3220 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond95_write_en = _guard3221;
assign cond95_clk = clk;
assign cond95_reset = reset;
assign cond95_in =
  _guard3222 ? idx_between_12_depth_plus_12_reg_out :
  1'd0;
assign cond109_write_en = _guard3223;
assign cond109_clk = clk;
assign cond109_reset = reset;
assign cond109_in =
  _guard3224 ? idx_between_depth_plus_8_depth_plus_9_reg_out :
  1'd0;
assign cond_wire111_in =
  _guard3225 ? idx_between_5_depth_plus_5_reg_out :
  _guard3228 ? cond111_out :
  1'd0;
assign cond_wire112_in =
  _guard3229 ? idx_between_9_depth_plus_9_reg_out :
  _guard3232 ? cond112_out :
  1'd0;
assign cond_wire118_in =
  _guard3235 ? cond118_out :
  _guard3236 ? idx_between_7_min_depth_4_plus_7_reg_out :
  1'd0;
assign cond_wire137_in =
  _guard3239 ? cond137_out :
  _guard3240 ? idx_between_depth_plus_15_depth_plus_16_reg_out :
  1'd0;
assign cond158_write_en = _guard3241;
assign cond158_clk = clk;
assign cond158_reset = reset;
assign cond158_in =
  _guard3242 ? idx_between_depth_plus_13_depth_plus_14_reg_out :
  1'd0;
assign cond159_write_en = _guard3243;
assign cond159_clk = clk;
assign cond159_reset = reset;
assign cond159_in =
  _guard3244 ? idx_between_10_min_depth_4_plus_10_reg_out :
  1'd0;
assign cond162_write_en = _guard3245;
assign cond162_clk = clk;
assign cond162_reset = reset;
assign cond162_in =
  _guard3246 ? idx_between_depth_plus_14_depth_plus_15_reg_out :
  1'd0;
assign cond164_write_en = _guard3247;
assign cond164_clk = clk;
assign cond164_reset = reset;
assign cond164_in =
  _guard3248 ? idx_between_11_depth_plus_11_reg_out :
  1'd0;
assign cond166_write_en = _guard3249;
assign cond166_clk = clk;
assign cond166_reset = reset;
assign cond166_in =
  _guard3250 ? idx_between_depth_plus_15_depth_plus_16_reg_out :
  1'd0;
assign cond_wire170_in =
  _guard3251 ? idx_between_depth_plus_16_depth_plus_17_reg_out :
  _guard3254 ? cond170_out :
  1'd0;
assign cond_wire175_in =
  _guard3255 ? idx_between_depth_plus_10_depth_plus_11_reg_out :
  _guard3258 ? cond175_out :
  1'd0;
assign cond180_write_en = _guard3259;
assign cond180_clk = clk;
assign cond180_reset = reset;
assign cond180_in =
  _guard3260 ? idx_between_8_min_depth_4_plus_8_reg_out :
  1'd0;
assign cond_wire197_in =
  _guard3261 ? idx_between_12_depth_plus_12_reg_out :
  _guard3264 ? cond197_out :
  1'd0;
assign cond198_write_en = _guard3265;
assign cond198_clk = clk;
assign cond198_reset = reset;
assign cond198_in =
  _guard3266 ? idx_between_16_depth_plus_16_reg_out :
  1'd0;
assign cond217_write_en = _guard3267;
assign cond217_clk = clk;
assign cond217_reset = reset;
assign cond217_in =
  _guard3268 ? idx_between_10_min_depth_4_plus_10_reg_out :
  1'd0;
assign cond222_write_en = _guard3269;
assign cond222_clk = clk;
assign cond222_reset = reset;
assign cond222_in =
  _guard3270 ? idx_between_11_depth_plus_11_reg_out :
  1'd0;
assign cond_wire222_in =
  _guard3271 ? idx_between_11_depth_plus_11_reg_out :
  _guard3274 ? cond222_out :
  1'd0;
assign cond_wire223_in =
  _guard3275 ? idx_between_15_depth_plus_15_reg_out :
  _guard3278 ? cond223_out :
  1'd0;
assign cond_wire225_in =
  _guard3279 ? idx_between_12_min_depth_4_plus_12_reg_out :
  _guard3282 ? cond225_out :
  1'd0;
assign cond_wire237_in =
  _guard3285 ? cond237_out :
  _guard3286 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond247_write_en = _guard3287;
assign cond247_clk = clk;
assign cond247_reset = reset;
assign cond247_in =
  _guard3288 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond_wire260_in =
  _guard3289 ? idx_between_17_depth_plus_17_reg_out :
  _guard3292 ? cond260_out :
  1'd0;
assign wrapper_early_reset_static_par_go_in = _guard3298;
assign depth_plus_7_left = depth;
assign depth_plus_7_right = 32'd7;
assign pe_0_2_mul_ready =
  _guard3303 ? 1'd1 :
  _guard3306 ? 1'd0 :
  1'd0;
assign pe_0_2_clk = clk;
assign pe_0_2_top =
  _guard3319 ? top_0_2_out :
  32'd0;
assign pe_0_2_left =
  _guard3332 ? left_0_2_out :
  32'd0;
assign pe_0_2_reset = reset;
assign pe_0_2_go = _guard3345;
assign pe_1_6_mul_ready =
  _guard3348 ? 1'd1 :
  _guard3351 ? 1'd0 :
  1'd0;
assign pe_1_6_clk = clk;
assign pe_1_6_top =
  _guard3364 ? top_1_6_out :
  32'd0;
assign pe_1_6_left =
  _guard3377 ? left_1_6_out :
  32'd0;
assign pe_1_6_reset = reset;
assign pe_1_6_go = _guard3390;
assign left_3_5_write_en = _guard3393;
assign left_3_5_clk = clk;
assign left_3_5_reset = reset;
assign left_3_5_in = left_3_4_out;
assign top_5_5_write_en = _guard3399;
assign top_5_5_clk = clk;
assign top_5_5_reset = reset;
assign top_5_5_in = top_4_5_out;
assign left_6_1_write_en = _guard3405;
assign left_6_1_clk = clk;
assign left_6_1_reset = reset;
assign left_6_1_in = left_6_0_out;
assign pe_6_5_mul_ready =
  _guard3411 ? 1'd1 :
  _guard3414 ? 1'd0 :
  1'd0;
assign pe_6_5_clk = clk;
assign pe_6_5_top =
  _guard3427 ? top_6_5_out :
  32'd0;
assign pe_6_5_left =
  _guard3440 ? left_6_5_out :
  32'd0;
assign pe_6_5_reset = reset;
assign pe_6_5_go = _guard3453;
assign left_6_7_write_en = _guard3456;
assign left_6_7_clk = clk;
assign left_6_7_reset = reset;
assign left_6_7_in = left_6_6_out;
assign pe_7_0_mul_ready =
  _guard3462 ? 1'd1 :
  _guard3465 ? 1'd0 :
  1'd0;
assign pe_7_0_clk = clk;
assign pe_7_0_top =
  _guard3478 ? top_7_0_out :
  32'd0;
assign pe_7_0_left =
  _guard3491 ? left_7_0_out :
  32'd0;
assign pe_7_0_reset = reset;
assign pe_7_0_go = _guard3504;
assign top_7_4_write_en = _guard3507;
assign top_7_4_clk = clk;
assign top_7_4_reset = reset;
assign top_7_4_in = top_6_4_out;
assign t0_idx_write_en = _guard3515;
assign t0_idx_clk = clk;
assign t0_idx_reset = reset;
assign t0_idx_in =
  _guard3516 ? 4'd0 :
  _guard3519 ? t0_add_out :
  'x;
assign t4_idx_write_en = _guard3524;
assign t4_idx_clk = clk;
assign t4_idx_reset = reset;
assign t4_idx_in =
  _guard3525 ? 4'd0 :
  _guard3528 ? t4_add_out :
  'x;
assign t6_idx_write_en = _guard3533;
assign t6_idx_clk = clk;
assign t6_idx_reset = reset;
assign t6_idx_in =
  _guard3534 ? 4'd0 :
  _guard3537 ? t6_add_out :
  'x;
assign l1_idx_write_en = _guard3542;
assign l1_idx_clk = clk;
assign l1_idx_reset = reset;
assign l1_idx_in =
  _guard3545 ? l1_add_out :
  _guard3546 ? 4'd0 :
  'x;
assign l5_add_left = 4'd1;
assign l5_add_right = l5_idx_out;
assign idx_add_left = idx_out;
assign idx_add_right = 32'd1;
assign index_lt_depth_plus_17_left = idx_add_out;
assign index_lt_depth_plus_17_right = depth_plus_17_out;
assign idx_between_2_min_depth_4_plus_2_comb_left = index_ge_2_out;
assign idx_between_2_min_depth_4_plus_2_comb_right = index_lt_min_depth_4_plus_2_out;
assign index_lt_depth_plus_18_left = idx_add_out;
assign index_lt_depth_plus_18_right = depth_plus_18_out;
assign idx_between_11_min_depth_4_plus_11_reg_write_en = _guard3563;
assign idx_between_11_min_depth_4_plus_11_reg_clk = clk;
assign idx_between_11_min_depth_4_plus_11_reg_reset = reset;
assign idx_between_11_min_depth_4_plus_11_reg_in =
  _guard3564 ? idx_between_11_min_depth_4_plus_11_comb_out :
  _guard3565 ? 1'd0 :
  'x;
assign index_ge_7_left = idx_add_out;
assign index_ge_7_right = 32'd7;
assign index_ge_depth_plus_18_left = idx_add_out;
assign index_ge_depth_plus_18_right = depth_plus_18_out;
assign idx_between_depth_plus_19_depth_plus_20_reg_write_en = _guard3572;
assign idx_between_depth_plus_19_depth_plus_20_reg_clk = clk;
assign idx_between_depth_plus_19_depth_plus_20_reg_reset = reset;
assign idx_between_depth_plus_19_depth_plus_20_reg_in =
  _guard3573 ? idx_between_depth_plus_19_depth_plus_20_comb_out :
  _guard3574 ? 1'd0 :
  'x;
assign idx_between_6_min_depth_4_plus_6_reg_write_en = _guard3577;
assign idx_between_6_min_depth_4_plus_6_reg_clk = clk;
assign idx_between_6_min_depth_4_plus_6_reg_reset = reset;
assign idx_between_6_min_depth_4_plus_6_reg_in =
  _guard3578 ? idx_between_6_min_depth_4_plus_6_comb_out :
  _guard3579 ? 1'd0 :
  'x;
assign idx_between_18_depth_plus_18_reg_write_en = _guard3582;
assign idx_between_18_depth_plus_18_reg_clk = clk;
assign idx_between_18_depth_plus_18_reg_reset = reset;
assign idx_between_18_depth_plus_18_reg_in =
  _guard3583 ? idx_between_18_depth_plus_18_comb_out :
  _guard3584 ? 1'd0 :
  'x;
assign idx_between_18_depth_plus_18_comb_left = index_ge_18_out;
assign idx_between_18_depth_plus_18_comb_right = index_lt_depth_plus_18_out;
assign cond3_write_en = _guard3587;
assign cond3_clk = clk;
assign cond3_reset = reset;
assign cond3_in =
  _guard3588 ? idx_between_depth_plus_5_depth_plus_6_reg_out :
  1'd0;
assign cond13_write_en = _guard3589;
assign cond13_clk = clk;
assign cond13_reset = reset;
assign cond13_in =
  _guard3590 ? idx_between_depth_plus_7_depth_plus_8_reg_out :
  1'd0;
assign cond29_write_en = _guard3591;
assign cond29_clk = clk;
assign cond29_reset = reset;
assign cond29_in =
  _guard3592 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond41_write_en = _guard3593;
assign cond41_clk = clk;
assign cond41_reset = reset;
assign cond41_in =
  _guard3594 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond54_write_en = _guard3595;
assign cond54_clk = clk;
assign cond54_reset = reset;
assign cond54_in =
  _guard3596 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond64_write_en = _guard3597;
assign cond64_clk = clk;
assign cond64_reset = reset;
assign cond64_in =
  _guard3598 ? idx_between_8_min_depth_4_plus_8_reg_out :
  1'd0;
assign cond67_write_en = _guard3599;
assign cond67_clk = clk;
assign cond67_reset = reset;
assign cond67_in =
  _guard3600 ? idx_between_depth_plus_12_depth_plus_13_reg_out :
  1'd0;
assign cond68_write_en = _guard3601;
assign cond68_clk = clk;
assign cond68_reset = reset;
assign cond68_in =
  _guard3602 ? idx_between_9_min_depth_4_plus_9_reg_out :
  1'd0;
assign cond77_write_en = _guard3603;
assign cond77_clk = clk;
assign cond77_reset = reset;
assign cond77_in =
  _guard3604 ? idx_between_4_min_depth_4_plus_4_reg_out :
  1'd0;
assign cond89_write_en = _guard3605;
assign cond89_clk = clk;
assign cond89_reset = reset;
assign cond89_in =
  _guard3606 ? idx_between_7_min_depth_4_plus_7_reg_out :
  1'd0;
assign cond94_write_en = _guard3607;
assign cond94_clk = clk;
assign cond94_reset = reset;
assign cond94_in =
  _guard3608 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire125_in =
  _guard3611 ? cond125_out :
  _guard3612 ? idx_between_depth_plus_12_depth_plus_13_reg_out :
  1'd0;
assign cond128_write_en = _guard3613;
assign cond128_clk = clk;
assign cond128_reset = reset;
assign cond128_in =
  _guard3614 ? idx_between_13_depth_plus_13_reg_out :
  1'd0;
assign cond131_write_en = _guard3615;
assign cond131_clk = clk;
assign cond131_reset = reset;
assign cond131_in =
  _guard3616 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond132_write_en = _guard3617;
assign cond132_clk = clk;
assign cond132_reset = reset;
assign cond132_in =
  _guard3618 ? idx_between_14_depth_plus_14_reg_out :
  1'd0;
assign cond_wire132_in =
  _guard3621 ? cond132_out :
  _guard3622 ? idx_between_14_depth_plus_14_reg_out :
  1'd0;
assign cond134_write_en = _guard3623;
assign cond134_clk = clk;
assign cond134_reset = reset;
assign cond134_in =
  _guard3624 ? idx_between_11_min_depth_4_plus_11_reg_out :
  1'd0;
assign cond136_write_en = _guard3625;
assign cond136_clk = clk;
assign cond136_reset = reset;
assign cond136_in =
  _guard3626 ? idx_between_15_depth_plus_15_reg_out :
  1'd0;
assign cond139_write_en = _guard3627;
assign cond139_clk = clk;
assign cond139_reset = reset;
assign cond139_in =
  _guard3628 ? idx_between_5_min_depth_4_plus_5_reg_out :
  1'd0;
assign cond140_write_en = _guard3629;
assign cond140_clk = clk;
assign cond140_reset = reset;
assign cond140_in =
  _guard3630 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond_wire142_in =
  _guard3631 ? idx_between_depth_plus_9_depth_plus_10_reg_out :
  _guard3634 ? cond142_out :
  1'd0;
assign cond_wire148_in =
  _guard3635 ? idx_between_7_depth_plus_7_reg_out :
  _guard3638 ? cond148_out :
  1'd0;
assign cond_wire151_in =
  _guard3639 ? idx_between_8_min_depth_4_plus_8_reg_out :
  _guard3642 ? cond151_out :
  1'd0;
assign cond_wire161_in =
  _guard3645 ? cond161_out :
  _guard3646 ? idx_between_14_depth_plus_14_reg_out :
  1'd0;
assign cond_wire162_in =
  _guard3649 ? cond162_out :
  _guard3650 ? idx_between_depth_plus_14_depth_plus_15_reg_out :
  1'd0;
assign cond_wire165_in =
  _guard3651 ? idx_between_15_depth_plus_15_reg_out :
  _guard3654 ? cond165_out :
  1'd0;
assign cond_wire171_in =
  _guard3657 ? cond171_out :
  _guard3658 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond172_write_en = _guard3659;
assign cond172_clk = clk;
assign cond172_reset = reset;
assign cond172_in =
  _guard3660 ? idx_between_6_min_depth_4_plus_6_reg_out :
  1'd0;
assign cond_wire177_in =
  _guard3663 ? cond177_out :
  _guard3664 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond183_write_en = _guard3665;
assign cond183_clk = clk;
assign cond183_reset = reset;
assign cond183_in =
  _guard3666 ? idx_between_depth_plus_12_depth_plus_13_reg_out :
  1'd0;
assign cond187_write_en = _guard3667;
assign cond187_clk = clk;
assign cond187_reset = reset;
assign cond187_in =
  _guard3668 ? idx_between_depth_plus_13_depth_plus_14_reg_out :
  1'd0;
assign cond190_write_en = _guard3669;
assign cond190_clk = clk;
assign cond190_reset = reset;
assign cond190_in =
  _guard3670 ? idx_between_14_depth_plus_14_reg_out :
  1'd0;
assign cond191_write_en = _guard3671;
assign cond191_clk = clk;
assign cond191_reset = reset;
assign cond191_in =
  _guard3672 ? idx_between_depth_plus_14_depth_plus_15_reg_out :
  1'd0;
assign cond223_write_en = _guard3673;
assign cond223_clk = clk;
assign cond223_reset = reset;
assign cond223_in =
  _guard3674 ? idx_between_15_depth_plus_15_reg_out :
  1'd0;
assign cond238_write_en = _guard3675;
assign cond238_clk = clk;
assign cond238_reset = reset;
assign cond238_in =
  _guard3676 ? idx_between_8_min_depth_4_plus_8_reg_out :
  1'd0;
assign cond244_write_en = _guard3677;
assign cond244_clk = clk;
assign cond244_reset = reset;
assign cond244_in =
  _guard3678 ? idx_between_13_depth_plus_13_reg_out :
  1'd0;
assign cond_wire252_in =
  _guard3679 ? idx_between_15_depth_plus_15_reg_out :
  _guard3682 ? cond252_out :
  1'd0;
assign cond_wire262_in =
  _guard3683 ? idx_between_14_min_depth_4_plus_14_reg_out :
  _guard3686 ? cond262_out :
  1'd0;
assign cond_wire264_in =
  _guard3689 ? cond264_out :
  _guard3690 ? idx_between_18_depth_plus_18_reg_out :
  1'd0;
assign cond265_write_en = _guard3691;
assign cond265_clk = clk;
assign cond265_reset = reset;
assign cond265_in =
  _guard3692 ? idx_between_depth_plus_18_depth_plus_19_reg_out :
  1'd0;
assign cond_wire267_in =
  _guard3693 ? idx_between_19_depth_plus_19_reg_out :
  _guard3696 ? cond267_out :
  1'd0;
assign wrapper_early_reset_static_par_done_in = _guard3699;
assign early_reset_static_par0_done_in = ud0_out;
assign tdcc_go_in = go;
assign left_0_7_write_en = _guard3702;
assign left_0_7_clk = clk;
assign left_0_7_reset = reset;
assign left_0_7_in = left_0_6_out;
assign pe_2_1_mul_ready =
  _guard3708 ? 1'd1 :
  _guard3711 ? 1'd0 :
  1'd0;
assign pe_2_1_clk = clk;
assign pe_2_1_top =
  _guard3724 ? top_2_1_out :
  32'd0;
assign pe_2_1_left =
  _guard3737 ? left_2_1_out :
  32'd0;
assign pe_2_1_reset = reset;
assign pe_2_1_go = _guard3750;
assign pe_2_3_mul_ready =
  _guard3753 ? 1'd1 :
  _guard3756 ? 1'd0 :
  1'd0;
assign pe_2_3_clk = clk;
assign pe_2_3_top =
  _guard3769 ? top_2_3_out :
  32'd0;
assign pe_2_3_left =
  _guard3782 ? left_2_3_out :
  32'd0;
assign pe_2_3_reset = reset;
assign pe_2_3_go = _guard3795;
assign pe_2_5_mul_ready =
  _guard3798 ? 1'd1 :
  _guard3801 ? 1'd0 :
  1'd0;
assign pe_2_5_clk = clk;
assign pe_2_5_top =
  _guard3814 ? top_2_5_out :
  32'd0;
assign pe_2_5_left =
  _guard3827 ? left_2_5_out :
  32'd0;
assign pe_2_5_reset = reset;
assign pe_2_5_go = _guard3840;
assign pe_3_1_mul_ready =
  _guard3843 ? 1'd1 :
  _guard3846 ? 1'd0 :
  1'd0;
assign pe_3_1_clk = clk;
assign pe_3_1_top =
  _guard3859 ? top_3_1_out :
  32'd0;
assign pe_3_1_left =
  _guard3872 ? left_3_1_out :
  32'd0;
assign pe_3_1_reset = reset;
assign pe_3_1_go = _guard3885;
assign top_3_4_write_en = _guard3888;
assign top_3_4_clk = clk;
assign top_3_4_reset = reset;
assign top_3_4_in = top_2_4_out;
assign pe_5_3_mul_ready =
  _guard3894 ? 1'd1 :
  _guard3897 ? 1'd0 :
  1'd0;
assign pe_5_3_clk = clk;
assign pe_5_3_top =
  _guard3910 ? top_5_3_out :
  32'd0;
assign pe_5_3_left =
  _guard3923 ? left_5_3_out :
  32'd0;
assign pe_5_3_reset = reset;
assign pe_5_3_go = _guard3936;
assign pe_5_5_mul_ready =
  _guard3939 ? 1'd1 :
  _guard3942 ? 1'd0 :
  1'd0;
assign pe_5_5_clk = clk;
assign pe_5_5_top =
  _guard3955 ? top_5_5_out :
  32'd0;
assign pe_5_5_left =
  _guard3968 ? left_5_5_out :
  32'd0;
assign pe_5_5_reset = reset;
assign pe_5_5_go = _guard3981;
assign pe_6_2_mul_ready =
  _guard3984 ? 1'd1 :
  _guard3987 ? 1'd0 :
  1'd0;
assign pe_6_2_clk = clk;
assign pe_6_2_top =
  _guard4000 ? top_6_2_out :
  32'd0;
assign pe_6_2_left =
  _guard4013 ? left_6_2_out :
  32'd0;
assign pe_6_2_reset = reset;
assign pe_6_2_go = _guard4026;
assign pe_6_3_mul_ready =
  _guard4029 ? 1'd1 :
  _guard4032 ? 1'd0 :
  1'd0;
assign pe_6_3_clk = clk;
assign pe_6_3_top =
  _guard4045 ? top_6_3_out :
  32'd0;
assign pe_6_3_left =
  _guard4058 ? left_6_3_out :
  32'd0;
assign pe_6_3_reset = reset;
assign pe_6_3_go = _guard4071;
assign left_7_1_write_en = _guard4074;
assign left_7_1_clk = clk;
assign left_7_1_reset = reset;
assign left_7_1_in = left_7_0_out;
assign left_7_3_write_en = _guard4080;
assign left_7_3_clk = clk;
assign left_7_3_reset = reset;
assign left_7_3_in = left_7_2_out;
assign top_7_5_write_en = _guard4086;
assign top_7_5_clk = clk;
assign top_7_5_reset = reset;
assign top_7_5_in = top_6_5_out;
assign t4_add_left = 4'd1;
assign t4_add_right = t4_idx_out;
assign t5_idx_write_en = _guard4100;
assign t5_idx_clk = clk;
assign t5_idx_reset = reset;
assign t5_idx_in =
  _guard4101 ? 4'd0 :
  _guard4104 ? t5_add_out :
  'x;
assign t6_add_left = 4'd1;
assign t6_add_right = t6_idx_out;
assign lt_iter_limit_left =
  _guard4111 ? depth :
  _guard4112 ? idx_add_out :
  'x;
assign lt_iter_limit_right =
  _guard4113 ? 32'd4 :
  _guard4114 ? iter_limit_out :
  'x;
assign idx_between_7_depth_plus_7_comb_left = index_ge_7_out;
assign idx_between_7_depth_plus_7_comb_right = index_lt_depth_plus_7_out;
assign index_lt_min_depth_4_plus_12_left = idx_add_out;
assign index_lt_min_depth_4_plus_12_right = min_depth_4_plus_12_out;
assign idx_between_17_depth_plus_17_reg_write_en = _guard4121;
assign idx_between_17_depth_plus_17_reg_clk = clk;
assign idx_between_17_depth_plus_17_reg_reset = reset;
assign idx_between_17_depth_plus_17_reg_in =
  _guard4122 ? 1'd0 :
  _guard4123 ? idx_between_17_depth_plus_17_comb_out :
  'x;
assign index_ge_17_left = idx_add_out;
assign index_ge_17_right = 32'd17;
assign idx_between_13_min_depth_4_plus_13_reg_write_en = _guard4128;
assign idx_between_13_min_depth_4_plus_13_reg_clk = clk;
assign idx_between_13_min_depth_4_plus_13_reg_reset = reset;
assign idx_between_13_min_depth_4_plus_13_reg_in =
  _guard4129 ? idx_between_13_min_depth_4_plus_13_comb_out :
  _guard4130 ? 1'd0 :
  'x;
assign index_lt_min_depth_4_plus_13_left = idx_add_out;
assign index_lt_min_depth_4_plus_13_right = min_depth_4_plus_13_out;
assign idx_between_9_min_depth_4_plus_9_reg_write_en = _guard4135;
assign idx_between_9_min_depth_4_plus_9_reg_clk = clk;
assign idx_between_9_min_depth_4_plus_9_reg_reset = reset;
assign idx_between_9_min_depth_4_plus_9_reg_in =
  _guard4136 ? idx_between_9_min_depth_4_plus_9_comb_out :
  _guard4137 ? 1'd0 :
  'x;
assign index_lt_min_depth_4_plus_9_left = idx_add_out;
assign index_lt_min_depth_4_plus_9_right = min_depth_4_plus_9_out;
assign idx_between_6_depth_plus_6_comb_left = index_ge_6_out;
assign idx_between_6_depth_plus_6_comb_right = index_lt_depth_plus_6_out;
assign index_ge_depth_plus_7_left = idx_add_out;
assign index_ge_depth_plus_7_right = depth_plus_7_out;
assign cond17_write_en = _guard4144;
assign cond17_clk = clk;
assign cond17_reset = reset;
assign cond17_in =
  _guard4145 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire22_in =
  _guard4146 ? idx_between_9_depth_plus_9_reg_out :
  _guard4149 ? cond22_out :
  1'd0;
assign cond23_write_en = _guard4150;
assign cond23_clk = clk;
assign cond23_reset = reset;
assign cond23_in =
  _guard4151 ? idx_between_depth_plus_9_depth_plus_10_reg_out :
  1'd0;
assign cond25_write_en = _guard4152;
assign cond25_clk = clk;
assign cond25_reset = reset;
assign cond25_in =
  _guard4153 ? idx_between_6_min_depth_4_plus_6_reg_out :
  1'd0;
assign cond_wire33_in =
  _guard4156 ? cond33_out :
  _guard4157 ? idx_between_depth_plus_11_depth_plus_12_reg_out :
  1'd0;
assign cond52_write_en = _guard4158;
assign cond52_clk = clk;
assign cond52_reset = reset;
assign cond52_in =
  _guard4159 ? idx_between_5_min_depth_4_plus_5_reg_out :
  1'd0;
assign cond56_write_en = _guard4160;
assign cond56_clk = clk;
assign cond56_reset = reset;
assign cond56_in =
  _guard4161 ? idx_between_6_min_depth_4_plus_6_reg_out :
  1'd0;
assign cond58_write_en = _guard4162;
assign cond58_clk = clk;
assign cond58_reset = reset;
assign cond58_in =
  _guard4163 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond75_write_en = _guard4164;
assign cond75_clk = clk;
assign cond75_reset = reset;
assign cond75_in =
  _guard4165 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond88_write_en = _guard4166;
assign cond88_clk = clk;
assign cond88_reset = reset;
assign cond88_in =
  _guard4167 ? idx_between_depth_plus_10_depth_plus_11_reg_out :
  1'd0;
assign cond93_write_en = _guard4168;
assign cond93_clk = clk;
assign cond93_reset = reset;
assign cond93_in =
  _guard4169 ? idx_between_8_min_depth_4_plus_8_reg_out :
  1'd0;
assign cond_wire98_in =
  _guard4172 ? cond98_out :
  _guard4173 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond_wire106_in =
  _guard4176 ? cond106_out :
  _guard4177 ? idx_between_4_min_depth_4_plus_4_reg_out :
  1'd0;
assign cond_wire120_in =
  _guard4178 ? idx_between_11_depth_plus_11_reg_out :
  _guard4181 ? cond120_out :
  1'd0;
assign cond124_write_en = _guard4182;
assign cond124_clk = clk;
assign cond124_reset = reset;
assign cond124_in =
  _guard4183 ? idx_between_12_depth_plus_12_reg_out :
  1'd0;
assign cond137_write_en = _guard4184;
assign cond137_clk = clk;
assign cond137_reset = reset;
assign cond137_in =
  _guard4185 ? idx_between_depth_plus_15_depth_plus_16_reg_out :
  1'd0;
assign cond155_write_en = _guard4186;
assign cond155_clk = clk;
assign cond155_reset = reset;
assign cond155_in =
  _guard4187 ? idx_between_9_min_depth_4_plus_9_reg_out :
  1'd0;
assign cond_wire176_in =
  _guard4188 ? idx_between_7_min_depth_4_plus_7_reg_out :
  _guard4191 ? cond176_out :
  1'd0;
assign cond188_write_en = _guard4192;
assign cond188_clk = clk;
assign cond188_reset = reset;
assign cond188_in =
  _guard4193 ? idx_between_10_min_depth_4_plus_10_reg_out :
  1'd0;
assign cond209_write_en = _guard4194;
assign cond209_clk = clk;
assign cond209_reset = reset;
assign cond209_in =
  _guard4195 ? idx_between_8_min_depth_4_plus_8_reg_out :
  1'd0;
assign cond_wire213_in =
  _guard4196 ? idx_between_9_min_depth_4_plus_9_reg_out :
  _guard4199 ? cond213_out :
  1'd0;
assign cond220_write_en = _guard4200;
assign cond220_clk = clk;
assign cond220_reset = reset;
assign cond220_in =
  _guard4201 ? idx_between_depth_plus_14_depth_plus_15_reg_out :
  1'd0;
assign cond_wire221_in =
  _guard4202 ? idx_between_11_min_depth_4_plus_11_reg_out :
  _guard4205 ? cond221_out :
  1'd0;
assign cond228_write_en = _guard4206;
assign cond228_clk = clk;
assign cond228_reset = reset;
assign cond228_in =
  _guard4207 ? idx_between_depth_plus_16_depth_plus_17_reg_out :
  1'd0;
assign cond232_write_en = _guard4208;
assign cond232_clk = clk;
assign cond232_reset = reset;
assign cond232_in =
  _guard4209 ? idx_between_depth_plus_17_depth_plus_18_reg_out :
  1'd0;
assign cond_wire236_in =
  _guard4212 ? cond236_out :
  _guard4213 ? idx_between_depth_plus_18_depth_plus_19_reg_out :
  1'd0;
assign cond258_write_en = _guard4214;
assign cond258_clk = clk;
assign cond258_reset = reset;
assign cond258_in =
  _guard4215 ? idx_between_13_min_depth_4_plus_13_reg_out :
  1'd0;
assign cond262_write_en = _guard4216;
assign cond262_clk = clk;
assign cond262_reset = reset;
assign cond262_in =
  _guard4217 ? idx_between_14_min_depth_4_plus_14_reg_out :
  1'd0;
assign fsm0_write_en = _guard4230;
assign fsm0_clk = clk;
assign fsm0_reset = reset;
assign fsm0_in =
  _guard4235 ? 2'd1 :
  _guard4236 ? 2'd0 :
  _guard4241 ? 2'd2 :
  2'd0;
assign depth_plus_8_left = depth;
assign depth_plus_8_right = 32'd8;
assign min_depth_4_plus_4_left = min_depth_4_out;
assign min_depth_4_plus_4_right = 32'd4;
assign depth_plus_0_left = depth;
assign depth_plus_0_right = 32'd0;
assign min_depth_4_plus_9_left = min_depth_4_out;
assign min_depth_4_plus_9_right = 32'd9;
assign pe_1_5_mul_ready =
  _guard4252 ? 1'd1 :
  _guard4255 ? 1'd0 :
  1'd0;
assign pe_1_5_clk = clk;
assign pe_1_5_top =
  _guard4268 ? top_1_5_out :
  32'd0;
assign pe_1_5_left =
  _guard4281 ? left_1_5_out :
  32'd0;
assign pe_1_5_reset = reset;
assign pe_1_5_go = _guard4294;
assign top_1_6_write_en = _guard4297;
assign top_1_6_clk = clk;
assign top_1_6_reset = reset;
assign top_1_6_in = top_0_6_out;
assign top_2_0_write_en = _guard4303;
assign top_2_0_clk = clk;
assign top_2_0_reset = reset;
assign top_2_0_in = top_1_0_out;
assign top_3_0_write_en = _guard4309;
assign top_3_0_clk = clk;
assign top_3_0_reset = reset;
assign top_3_0_in = top_2_0_out;
assign top_3_1_write_en = _guard4315;
assign top_3_1_clk = clk;
assign top_3_1_reset = reset;
assign top_3_1_in = top_2_1_out;
assign pe_4_6_mul_ready =
  _guard4321 ? 1'd1 :
  _guard4324 ? 1'd0 :
  1'd0;
assign pe_4_6_clk = clk;
assign pe_4_6_top =
  _guard4337 ? top_4_6_out :
  32'd0;
assign pe_4_6_left =
  _guard4350 ? left_4_6_out :
  32'd0;
assign pe_4_6_reset = reset;
assign pe_4_6_go = _guard4363;
assign top_5_2_write_en = _guard4366;
assign top_5_2_clk = clk;
assign top_5_2_reset = reset;
assign top_5_2_in = top_4_2_out;
assign top_5_4_write_en = _guard4372;
assign top_5_4_clk = clk;
assign top_5_4_reset = reset;
assign top_5_4_in = top_4_4_out;
assign left_7_7_write_en = _guard4378;
assign left_7_7_clk = clk;
assign left_7_7_reset = reset;
assign left_7_7_in = left_7_6_out;
assign t7_add_left = 4'd1;
assign t7_add_right = t7_idx_out;
assign l4_idx_write_en = _guard4392;
assign l4_idx_clk = clk;
assign l4_idx_reset = reset;
assign l4_idx_in =
  _guard4393 ? 4'd0 :
  _guard4396 ? l4_add_out :
  'x;
assign idx_write_en = _guard4399;
assign idx_clk = clk;
assign idx_reset = reset;
assign idx_in =
  _guard4400 ? 32'd0 :
  _guard4401 ? idx_add_out :
  'x;
assign idx_between_depth_plus_16_depth_plus_17_reg_write_en = _guard4404;
assign idx_between_depth_plus_16_depth_plus_17_reg_clk = clk;
assign idx_between_depth_plus_16_depth_plus_17_reg_reset = reset;
assign idx_between_depth_plus_16_depth_plus_17_reg_in =
  _guard4405 ? idx_between_depth_plus_16_depth_plus_17_comb_out :
  _guard4406 ? 1'd0 :
  'x;
assign idx_between_7_depth_plus_7_reg_write_en = _guard4409;
assign idx_between_7_depth_plus_7_reg_clk = clk;
assign idx_between_7_depth_plus_7_reg_reset = reset;
assign idx_between_7_depth_plus_7_reg_in =
  _guard4410 ? idx_between_7_depth_plus_7_comb_out :
  _guard4411 ? 1'd0 :
  'x;
assign index_lt_depth_plus_3_left = idx_add_out;
assign index_lt_depth_plus_3_right = depth_plus_3_out;
assign idx_between_depth_plus_10_depth_plus_11_reg_write_en = _guard4416;
assign idx_between_depth_plus_10_depth_plus_11_reg_clk = clk;
assign idx_between_depth_plus_10_depth_plus_11_reg_reset = reset;
assign idx_between_depth_plus_10_depth_plus_11_reg_in =
  _guard4417 ? 1'd0 :
  _guard4418 ? idx_between_depth_plus_10_depth_plus_11_comb_out :
  'x;
assign idx_between_depth_plus_19_depth_plus_20_comb_left = index_ge_depth_plus_19_out;
assign idx_between_depth_plus_19_depth_plus_20_comb_right = index_lt_depth_plus_20_out;
assign idx_between_4_depth_plus_4_comb_left = index_ge_4_out;
assign idx_between_4_depth_plus_4_comb_right = index_lt_depth_plus_4_out;
assign idx_between_14_depth_plus_14_comb_left = index_ge_14_out;
assign idx_between_14_depth_plus_14_comb_right = index_lt_depth_plus_14_out;
assign index_lt_min_depth_4_plus_5_left = idx_add_out;
assign index_lt_min_depth_4_plus_5_right = min_depth_4_plus_5_out;
assign index_lt_depth_plus_0_left = idx_add_out;
assign index_lt_depth_plus_0_right = depth_plus_0_out;
assign idx_between_9_depth_plus_9_reg_write_en = _guard4431;
assign idx_between_9_depth_plus_9_reg_clk = clk;
assign idx_between_9_depth_plus_9_reg_reset = reset;
assign idx_between_9_depth_plus_9_reg_in =
  _guard4432 ? 1'd0 :
  _guard4433 ? idx_between_9_depth_plus_9_comb_out :
  'x;
assign idx_between_9_min_depth_4_plus_9_comb_left = index_ge_9_out;
assign idx_between_9_min_depth_4_plus_9_comb_right = index_lt_min_depth_4_plus_9_out;
assign idx_between_1_depth_plus_1_comb_left = index_ge_1_out;
assign idx_between_1_depth_plus_1_comb_right = index_lt_depth_plus_1_out;
assign index_ge_depth_plus_11_left = idx_add_out;
assign index_ge_depth_plus_11_right = depth_plus_11_out;
assign idx_between_depth_plus_11_depth_plus_12_comb_left = index_ge_depth_plus_11_out;
assign idx_between_depth_plus_11_depth_plus_12_comb_right = index_lt_depth_plus_12_out;
assign cond7_write_en = _guard4442;
assign cond7_clk = clk;
assign cond7_reset = reset;
assign cond7_in =
  _guard4443 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire8_in =
  _guard4444 ? idx_between_depth_plus_6_depth_plus_7_reg_out :
  _guard4447 ? cond8_out :
  1'd0;
assign cond9_write_en = _guard4448;
assign cond9_clk = clk;
assign cond9_reset = reset;
assign cond9_in =
  _guard4449 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond14_write_en = _guard4450;
assign cond14_clk = clk;
assign cond14_reset = reset;
assign cond14_in =
  _guard4451 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond_wire20_in =
  _guard4452 ? idx_between_5_min_depth_4_plus_5_reg_out :
  _guard4455 ? cond20_out :
  1'd0;
assign cond27_write_en = _guard4456;
assign cond27_clk = clk;
assign cond27_reset = reset;
assign cond27_in =
  _guard4457 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond32_write_en = _guard4458;
assign cond32_clk = clk;
assign cond32_reset = reset;
assign cond32_in =
  _guard4459 ? idx_between_11_depth_plus_11_reg_out :
  1'd0;
assign cond_wire37_in =
  _guard4460 ? idx_between_12_depth_plus_12_reg_out :
  _guard4463 ? cond37_out :
  1'd0;
assign cond50_write_en = _guard4464;
assign cond50_clk = clk;
assign cond50_reset = reset;
assign cond50_in =
  _guard4465 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire60_in =
  _guard4468 ? cond60_out :
  _guard4469 ? idx_between_7_min_depth_4_plus_7_reg_out :
  1'd0;
assign cond_wire64_in =
  _guard4470 ? idx_between_8_min_depth_4_plus_8_reg_out :
  _guard4473 ? cond64_out :
  1'd0;
assign cond_wire81_in =
  _guard4476 ? cond81_out :
  _guard4477 ? idx_between_5_min_depth_4_plus_5_reg_out :
  1'd0;
assign cond_wire82_in =
  _guard4480 ? cond82_out :
  _guard4481 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond83_write_en = _guard4482;
assign cond83_clk = clk;
assign cond83_reset = reset;
assign cond83_in =
  _guard4483 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond_wire86_in =
  _guard4486 ? cond86_out :
  _guard4487 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire87_in =
  _guard4488 ? idx_between_10_depth_plus_10_reg_out :
  _guard4491 ? cond87_out :
  1'd0;
assign cond91_write_en = _guard4492;
assign cond91_clk = clk;
assign cond91_reset = reset;
assign cond91_in =
  _guard4493 ? idx_between_11_depth_plus_11_reg_out :
  1'd0;
assign cond_wire105_in =
  _guard4496 ? cond105_out :
  _guard4497 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond116_write_en = _guard4498;
assign cond116_clk = clk;
assign cond116_reset = reset;
assign cond116_in =
  _guard4499 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond_wire117_in =
  _guard4500 ? idx_between_depth_plus_10_depth_plus_11_reg_out :
  _guard4503 ? cond117_out :
  1'd0;
assign cond_wire138_in =
  _guard4504 ? idx_between_4_depth_plus_4_reg_out :
  _guard4507 ? cond138_out :
  1'd0;
assign cond_wire140_in =
  _guard4510 ? cond140_out :
  _guard4511 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond_wire156_in =
  _guard4512 ? idx_between_9_depth_plus_9_reg_out :
  _guard4515 ? cond156_out :
  1'd0;
assign cond161_write_en = _guard4516;
assign cond161_clk = clk;
assign cond161_reset = reset;
assign cond161_in =
  _guard4517 ? idx_between_14_depth_plus_14_reg_out :
  1'd0;
assign cond174_write_en = _guard4518;
assign cond174_clk = clk;
assign cond174_reset = reset;
assign cond174_in =
  _guard4519 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond176_write_en = _guard4520;
assign cond176_clk = clk;
assign cond176_reset = reset;
assign cond176_in =
  _guard4521 ? idx_between_7_min_depth_4_plus_7_reg_out :
  1'd0;
assign cond_wire187_in =
  _guard4524 ? cond187_out :
  _guard4525 ? idx_between_depth_plus_13_depth_plus_14_reg_out :
  1'd0;
assign cond_wire190_in =
  _guard4528 ? cond190_out :
  _guard4529 ? idx_between_14_depth_plus_14_reg_out :
  1'd0;
assign cond194_write_en = _guard4530;
assign cond194_clk = clk;
assign cond194_reset = reset;
assign cond194_in =
  _guard4531 ? idx_between_15_depth_plus_15_reg_out :
  1'd0;
assign cond201_write_en = _guard4532;
assign cond201_clk = clk;
assign cond201_reset = reset;
assign cond201_in =
  _guard4533 ? idx_between_13_depth_plus_13_reg_out :
  1'd0;
assign cond205_write_en = _guard4534;
assign cond205_clk = clk;
assign cond205_reset = reset;
assign cond205_in =
  _guard4535 ? idx_between_7_min_depth_4_plus_7_reg_out :
  1'd0;
assign cond_wire207_in =
  _guard4536 ? idx_between_11_depth_plus_11_reg_out :
  _guard4539 ? cond207_out :
  1'd0;
assign cond_wire209_in =
  _guard4540 ? idx_between_8_min_depth_4_plus_8_reg_out :
  _guard4543 ? cond209_out :
  1'd0;
assign cond219_write_en = _guard4544;
assign cond219_clk = clk;
assign cond219_reset = reset;
assign cond219_in =
  _guard4545 ? idx_between_14_depth_plus_14_reg_out :
  1'd0;
assign cond221_write_en = _guard4546;
assign cond221_clk = clk;
assign cond221_reset = reset;
assign cond221_in =
  _guard4547 ? idx_between_11_min_depth_4_plus_11_reg_out :
  1'd0;
assign cond225_write_en = _guard4548;
assign cond225_clk = clk;
assign cond225_reset = reset;
assign cond225_in =
  _guard4549 ? idx_between_12_min_depth_4_plus_12_reg_out :
  1'd0;
assign cond256_write_en = _guard4550;
assign cond256_clk = clk;
assign cond256_reset = reset;
assign cond256_in =
  _guard4551 ? idx_between_16_depth_plus_16_reg_out :
  1'd0;
assign min_depth_4_write_en = _guard4552;
assign min_depth_4_clk = clk;
assign min_depth_4_reset = reset;
assign min_depth_4_in =
  _guard4555 ? depth :
  _guard4559 ? 32'd4 :
  'x;
assign min_depth_4_plus_11_left = min_depth_4_out;
assign min_depth_4_plus_11_right = 32'd11;
assign depth_plus_14_left = depth;
assign depth_plus_14_right = 32'd14;
assign min_depth_4_plus_6_left = min_depth_4_out;
assign min_depth_4_plus_6_right = 32'd6;
assign top_0_1_write_en = _guard4568;
assign top_0_1_clk = clk;
assign top_0_1_reset = reset;
assign top_0_1_in = t1_read_data;
assign left_0_2_write_en = _guard4574;
assign left_0_2_clk = clk;
assign left_0_2_reset = reset;
assign left_0_2_in = left_0_1_out;
assign pe_0_4_mul_ready =
  _guard4580 ? 1'd1 :
  _guard4583 ? 1'd0 :
  1'd0;
assign pe_0_4_clk = clk;
assign pe_0_4_top =
  _guard4596 ? top_0_4_out :
  32'd0;
assign pe_0_4_left =
  _guard4609 ? left_0_4_out :
  32'd0;
assign pe_0_4_reset = reset;
assign pe_0_4_go = _guard4622;
assign top_2_3_write_en = _guard4625;
assign top_2_3_clk = clk;
assign top_2_3_reset = reset;
assign top_2_3_in = top_1_3_out;
assign pe_2_6_mul_ready =
  _guard4631 ? 1'd1 :
  _guard4634 ? 1'd0 :
  1'd0;
assign pe_2_6_clk = clk;
assign pe_2_6_top =
  _guard4647 ? top_2_6_out :
  32'd0;
assign pe_2_6_left =
  _guard4660 ? left_2_6_out :
  32'd0;
assign pe_2_6_reset = reset;
assign pe_2_6_go = _guard4673;
assign left_3_0_write_en = _guard4676;
assign left_3_0_clk = clk;
assign left_3_0_reset = reset;
assign left_3_0_in = l3_read_data;
assign pe_4_2_mul_ready =
  _guard4682 ? 1'd1 :
  _guard4685 ? 1'd0 :
  1'd0;
assign pe_4_2_clk = clk;
assign pe_4_2_top =
  _guard4698 ? top_4_2_out :
  32'd0;
assign pe_4_2_left =
  _guard4711 ? left_4_2_out :
  32'd0;
assign pe_4_2_reset = reset;
assign pe_4_2_go = _guard4724;
assign top_5_1_write_en = _guard4727;
assign top_5_1_clk = clk;
assign top_5_1_reset = reset;
assign top_5_1_in = top_4_1_out;
assign left_5_4_write_en = _guard4733;
assign left_5_4_clk = clk;
assign left_5_4_reset = reset;
assign left_5_4_in = left_5_3_out;
assign pe_6_7_mul_ready =
  _guard4739 ? 1'd1 :
  _guard4742 ? 1'd0 :
  1'd0;
assign pe_6_7_clk = clk;
assign pe_6_7_top =
  _guard4755 ? top_6_7_out :
  32'd0;
assign pe_6_7_left =
  _guard4768 ? left_6_7_out :
  32'd0;
assign pe_6_7_reset = reset;
assign pe_6_7_go = _guard4781;
assign l7_add_left = 4'd1;
assign l7_add_right = l7_idx_out;
assign idx_between_depth_plus_17_depth_plus_18_comb_left = index_ge_depth_plus_17_out;
assign idx_between_depth_plus_17_depth_plus_18_comb_right = index_lt_depth_plus_18_out;
assign idx_between_11_min_depth_4_plus_11_comb_left = index_ge_11_out;
assign idx_between_11_min_depth_4_plus_11_comb_right = index_lt_min_depth_4_plus_11_out;
assign idx_between_depth_plus_13_depth_plus_14_comb_left = index_ge_depth_plus_13_out;
assign idx_between_depth_plus_13_depth_plus_14_comb_right = index_lt_depth_plus_14_out;
assign idx_between_3_min_depth_4_plus_3_reg_write_en = _guard4796;
assign idx_between_3_min_depth_4_plus_3_reg_clk = clk;
assign idx_between_3_min_depth_4_plus_3_reg_reset = reset;
assign idx_between_3_min_depth_4_plus_3_reg_in =
  _guard4797 ? idx_between_3_min_depth_4_plus_3_comb_out :
  _guard4798 ? 1'd0 :
  'x;
assign index_lt_depth_plus_15_left = idx_add_out;
assign index_lt_depth_plus_15_right = depth_plus_15_out;
assign index_ge_4_left = idx_add_out;
assign index_ge_4_right = 32'd4;
assign idx_between_5_min_depth_4_plus_5_reg_write_en = _guard4805;
assign idx_between_5_min_depth_4_plus_5_reg_clk = clk;
assign idx_between_5_min_depth_4_plus_5_reg_reset = reset;
assign idx_between_5_min_depth_4_plus_5_reg_in =
  _guard4806 ? 1'd0 :
  _guard4807 ? idx_between_5_min_depth_4_plus_5_comb_out :
  'x;
assign index_ge_1_left = idx_add_out;
assign index_ge_1_right = 32'd1;
assign idx_between_10_min_depth_4_plus_10_reg_write_en = _guard4812;
assign idx_between_10_min_depth_4_plus_10_reg_clk = clk;
assign idx_between_10_min_depth_4_plus_10_reg_reset = reset;
assign idx_between_10_min_depth_4_plus_10_reg_in =
  _guard4813 ? 1'd0 :
  _guard4814 ? idx_between_10_min_depth_4_plus_10_comb_out :
  'x;
assign cond4_write_en = _guard4815;
assign cond4_clk = clk;
assign cond4_reset = reset;
assign cond4_in =
  _guard4816 ? idx_between_1_depth_plus_1_reg_out :
  1'd0;
assign cond5_write_en = _guard4817;
assign cond5_clk = clk;
assign cond5_reset = reset;
assign cond5_in =
  _guard4818 ? idx_between_2_min_depth_4_plus_2_reg_out :
  1'd0;
assign cond_wire6_in =
  _guard4821 ? cond6_out :
  _guard4822 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond20_write_en = _guard4823;
assign cond20_clk = clk;
assign cond20_reset = reset;
assign cond20_in =
  _guard4824 ? idx_between_5_min_depth_4_plus_5_reg_out :
  1'd0;
assign cond_wire36_in =
  _guard4827 ? cond36_out :
  _guard4828 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond46_write_en = _guard4829;
assign cond46_clk = clk;
assign cond46_reset = reset;
assign cond46_in =
  _guard4830 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond_wire62_in =
  _guard4831 ? idx_between_11_depth_plus_11_reg_out :
  _guard4834 ? cond62_out :
  1'd0;
assign cond63_write_en = _guard4835;
assign cond63_clk = clk;
assign cond63_reset = reset;
assign cond63_in =
  _guard4836 ? idx_between_depth_plus_11_depth_plus_12_reg_out :
  1'd0;
assign cond_wire66_in =
  _guard4837 ? idx_between_12_depth_plus_12_reg_out :
  _guard4840 ? cond66_out :
  1'd0;
assign cond_wire74_in =
  _guard4843 ? cond74_out :
  _guard4844 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond_wire75_in =
  _guard4847 ? cond75_out :
  _guard4848 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond78_write_en = _guard4849;
assign cond78_clk = clk;
assign cond78_reset = reset;
assign cond78_in =
  _guard4850 ? idx_between_4_depth_plus_4_reg_out :
  1'd0;
assign cond90_write_en = _guard4851;
assign cond90_clk = clk;
assign cond90_reset = reset;
assign cond90_in =
  _guard4852 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond_wire92_in =
  _guard4855 ? cond92_out :
  _guard4856 ? idx_between_depth_plus_11_depth_plus_12_reg_out :
  1'd0;
assign cond101_write_en = _guard4857;
assign cond101_clk = clk;
assign cond101_reset = reset;
assign cond101_in =
  _guard4858 ? idx_between_10_min_depth_4_plus_10_reg_out :
  1'd0;
assign cond106_write_en = _guard4859;
assign cond106_clk = clk;
assign cond106_reset = reset;
assign cond106_in =
  _guard4860 ? idx_between_4_min_depth_4_plus_4_reg_out :
  1'd0;
assign cond_wire108_in =
  _guard4861 ? idx_between_8_depth_plus_8_reg_out :
  _guard4864 ? cond108_out :
  1'd0;
assign cond112_write_en = _guard4865;
assign cond112_clk = clk;
assign cond112_reset = reset;
assign cond112_in =
  _guard4866 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond122_write_en = _guard4867;
assign cond122_clk = clk;
assign cond122_reset = reset;
assign cond122_in =
  _guard4868 ? idx_between_8_min_depth_4_plus_8_reg_out :
  1'd0;
assign cond_wire122_in =
  _guard4869 ? idx_between_8_min_depth_4_plus_8_reg_out :
  _guard4872 ? cond122_out :
  1'd0;
assign cond_wire128_in =
  _guard4873 ? idx_between_13_depth_plus_13_reg_out :
  _guard4876 ? cond128_out :
  1'd0;
assign cond_wire139_in =
  _guard4879 ? cond139_out :
  _guard4880 ? idx_between_5_min_depth_4_plus_5_reg_out :
  1'd0;
assign cond143_write_en = _guard4881;
assign cond143_clk = clk;
assign cond143_reset = reset;
assign cond143_in =
  _guard4882 ? idx_between_6_min_depth_4_plus_6_reg_out :
  1'd0;
assign cond_wire143_in =
  _guard4883 ? idx_between_6_min_depth_4_plus_6_reg_out :
  _guard4886 ? cond143_out :
  1'd0;
assign cond148_write_en = _guard4887;
assign cond148_clk = clk;
assign cond148_reset = reset;
assign cond148_in =
  _guard4888 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond152_write_en = _guard4889;
assign cond152_clk = clk;
assign cond152_reset = reset;
assign cond152_in =
  _guard4890 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire172_in =
  _guard4891 ? idx_between_6_min_depth_4_plus_6_reg_out :
  _guard4894 ? cond172_out :
  1'd0;
assign cond_wire178_in =
  _guard4895 ? idx_between_11_depth_plus_11_reg_out :
  _guard4898 ? cond178_out :
  1'd0;
assign cond_wire181_in =
  _guard4901 ? cond181_out :
  _guard4902 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire189_in =
  _guard4905 ? cond189_out :
  _guard4906 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond192_write_en = _guard4907;
assign cond192_clk = clk;
assign cond192_reset = reset;
assign cond192_in =
  _guard4908 ? idx_between_11_min_depth_4_plus_11_reg_out :
  1'd0;
assign cond196_write_en = _guard4909;
assign cond196_clk = clk;
assign cond196_reset = reset;
assign cond196_in =
  _guard4910 ? idx_between_12_min_depth_4_plus_12_reg_out :
  1'd0;
assign cond203_write_en = _guard4911;
assign cond203_clk = clk;
assign cond203_reset = reset;
assign cond203_in =
  _guard4912 ? idx_between_depth_plus_17_depth_plus_18_reg_out :
  1'd0;
assign cond_wire203_in =
  _guard4915 ? cond203_out :
  _guard4916 ? idx_between_depth_plus_17_depth_plus_18_reg_out :
  1'd0;
assign cond208_write_en = _guard4917;
assign cond208_clk = clk;
assign cond208_reset = reset;
assign cond208_in =
  _guard4918 ? idx_between_depth_plus_11_depth_plus_12_reg_out :
  1'd0;
assign cond_wire210_in =
  _guard4919 ? idx_between_8_depth_plus_8_reg_out :
  _guard4922 ? cond210_out :
  1'd0;
assign cond_wire214_in =
  _guard4925 ? cond214_out :
  _guard4926 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond_wire233_in =
  _guard4927 ? idx_between_14_min_depth_4_plus_14_reg_out :
  _guard4930 ? cond233_out :
  1'd0;
assign cond235_write_en = _guard4931;
assign cond235_clk = clk;
assign cond235_reset = reset;
assign cond235_in =
  _guard4932 ? idx_between_18_depth_plus_18_reg_out :
  1'd0;
assign cond_wire248_in =
  _guard4935 ? cond248_out :
  _guard4936 ? idx_between_14_depth_plus_14_reg_out :
  1'd0;
assign cond250_write_en = _guard4937;
assign cond250_clk = clk;
assign cond250_reset = reset;
assign cond250_in =
  _guard4938 ? idx_between_11_min_depth_4_plus_11_reg_out :
  1'd0;
assign cond252_write_en = _guard4939;
assign cond252_clk = clk;
assign cond252_reset = reset;
assign cond252_in =
  _guard4940 ? idx_between_15_depth_plus_15_reg_out :
  1'd0;
assign cond_wire253_in =
  _guard4941 ? idx_between_depth_plus_15_depth_plus_16_reg_out :
  _guard4944 ? cond253_out :
  1'd0;
assign cond_wire256_in =
  _guard4945 ? idx_between_16_depth_plus_16_reg_out :
  _guard4948 ? cond256_out :
  1'd0;
assign cond_wire258_in =
  _guard4949 ? idx_between_13_min_depth_4_plus_13_reg_out :
  _guard4952 ? cond258_out :
  1'd0;
assign cond_wire268_in =
  _guard4953 ? idx_between_depth_plus_19_depth_plus_20_reg_out :
  _guard4956 ? cond268_out :
  1'd0;
assign adder0_left =
  _guard4957 ? fsm_out :
  1'd0;
assign adder0_right = _guard4958;
assign early_reset_static_par_done_in = ud_out;
assign depth_plus_3_left = depth;
assign depth_plus_3_right = 32'd3;
assign min_depth_4_plus_13_left = min_depth_4_out;
assign min_depth_4_plus_13_right = 32'd13;
assign top_0_2_write_en = _guard4965;
assign top_0_2_clk = clk;
assign top_0_2_reset = reset;
assign top_0_2_in = t2_read_data;
assign top_1_1_write_en = _guard4971;
assign top_1_1_clk = clk;
assign top_1_1_reset = reset;
assign top_1_1_in = top_0_1_out;
assign left_3_2_write_en = _guard4977;
assign left_3_2_clk = clk;
assign left_3_2_reset = reset;
assign left_3_2_in = left_3_1_out;
assign left_3_4_write_en = _guard4983;
assign left_3_4_clk = clk;
assign left_3_4_reset = reset;
assign left_3_4_in = left_3_3_out;
assign top_4_1_write_en = _guard4989;
assign top_4_1_clk = clk;
assign top_4_1_reset = reset;
assign top_4_1_in = top_3_1_out;
assign top_4_2_write_en = _guard4995;
assign top_4_2_clk = clk;
assign top_4_2_reset = reset;
assign top_4_2_in = top_3_2_out;
assign top_6_4_write_en = _guard5001;
assign top_6_4_clk = clk;
assign top_6_4_reset = reset;
assign top_6_4_in = top_5_4_out;
assign top_6_5_write_en = _guard5007;
assign top_6_5_clk = clk;
assign top_6_5_reset = reset;
assign top_6_5_in = top_5_5_out;
assign left_6_6_write_en = _guard5013;
assign left_6_6_clk = clk;
assign left_6_6_reset = reset;
assign left_6_6_in = left_6_5_out;
assign left_7_2_write_en = _guard5019;
assign left_7_2_clk = clk;
assign left_7_2_reset = reset;
assign left_7_2_in = left_7_1_out;
assign pe_7_5_mul_ready =
  _guard5025 ? 1'd1 :
  _guard5028 ? 1'd0 :
  1'd0;
assign pe_7_5_clk = clk;
assign pe_7_5_top =
  _guard5041 ? top_7_5_out :
  32'd0;
assign pe_7_5_left =
  _guard5054 ? left_7_5_out :
  32'd0;
assign pe_7_5_reset = reset;
assign pe_7_5_go = _guard5067;
assign pe_7_6_mul_ready =
  _guard5070 ? 1'd1 :
  _guard5073 ? 1'd0 :
  1'd0;
assign pe_7_6_clk = clk;
assign pe_7_6_top =
  _guard5086 ? top_7_6_out :
  32'd0;
assign pe_7_6_left =
  _guard5099 ? left_7_6_out :
  32'd0;
assign pe_7_6_reset = reset;
assign pe_7_6_go = _guard5112;
assign t0_add_left = 4'd1;
assign t0_add_right = t0_idx_out;
assign l0_add_left = 4'd1;
assign l0_add_right = l0_idx_out;
assign idx_between_depth_plus_17_depth_plus_18_reg_write_en = _guard5127;
assign idx_between_depth_plus_17_depth_plus_18_reg_clk = clk;
assign idx_between_depth_plus_17_depth_plus_18_reg_reset = reset;
assign idx_between_depth_plus_17_depth_plus_18_reg_in =
  _guard5128 ? idx_between_depth_plus_17_depth_plus_18_comb_out :
  _guard5129 ? 1'd0 :
  'x;
assign index_ge_11_left = idx_add_out;
assign index_ge_11_right = 32'd11;
assign index_lt_min_depth_4_plus_14_left = idx_add_out;
assign index_lt_min_depth_4_plus_14_right = min_depth_4_plus_14_out;
assign index_ge_9_left = idx_add_out;
assign index_ge_9_right = 32'd9;
assign idx_between_1_min_depth_4_plus_1_comb_left = index_ge_1_out;
assign idx_between_1_min_depth_4_plus_1_comb_right = index_lt_min_depth_4_plus_1_out;
assign idx_between_depth_plus_7_depth_plus_8_comb_left = index_ge_depth_plus_7_out;
assign idx_between_depth_plus_7_depth_plus_8_comb_right = index_lt_depth_plus_8_out;
assign cond_wire2_in =
  _guard5142 ? cond2_out :
  _guard5143 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond_wire9_in =
  _guard5146 ? cond9_out :
  _guard5147 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond10_write_en = _guard5148;
assign cond10_clk = clk;
assign cond10_reset = reset;
assign cond10_in =
  _guard5149 ? idx_between_3_min_depth_4_plus_3_reg_out :
  1'd0;
assign cond_wire11_in =
  _guard5152 ? cond11_out :
  _guard5153 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond21_write_en = _guard5154;
assign cond21_clk = clk;
assign cond21_reset = reset;
assign cond21_in =
  _guard5155 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond24_write_en = _guard5156;
assign cond24_clk = clk;
assign cond24_reset = reset;
assign cond24_in =
  _guard5157 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond31_write_en = _guard5158;
assign cond31_clk = clk;
assign cond31_reset = reset;
assign cond31_in =
  _guard5159 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond36_write_en = _guard5160;
assign cond36_clk = clk;
assign cond36_reset = reset;
assign cond36_in =
  _guard5161 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire41_in =
  _guard5164 ? cond41_out :
  _guard5165 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond_wire45_in =
  _guard5168 ? cond45_out :
  _guard5169 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond51_write_en = _guard5170;
assign cond51_clk = clk;
assign cond51_reset = reset;
assign cond51_in =
  _guard5171 ? idx_between_depth_plus_8_depth_plus_9_reg_out :
  1'd0;
assign cond_wire57_in =
  _guard5174 ? cond57_out :
  _guard5175 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire58_in =
  _guard5178 ? cond58_out :
  _guard5179 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond61_write_en = _guard5180;
assign cond61_clk = clk;
assign cond61_reset = reset;
assign cond61_in =
  _guard5181 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond80_write_en = _guard5182;
assign cond80_clk = clk;
assign cond80_reset = reset;
assign cond80_in =
  _guard5183 ? idx_between_depth_plus_8_depth_plus_9_reg_out :
  1'd0;
assign cond_wire80_in =
  _guard5184 ? idx_between_depth_plus_8_depth_plus_9_reg_out :
  _guard5187 ? cond80_out :
  1'd0;
assign cond86_write_en = _guard5188;
assign cond86_clk = clk;
assign cond86_reset = reset;
assign cond86_in =
  _guard5189 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond97_write_en = _guard5190;
assign cond97_clk = clk;
assign cond97_reset = reset;
assign cond97_in =
  _guard5191 ? idx_between_9_min_depth_4_plus_9_reg_out :
  1'd0;
assign cond_wire123_in =
  _guard5194 ? cond123_out :
  _guard5195 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond127_write_en = _guard5196;
assign cond127_clk = clk;
assign cond127_reset = reset;
assign cond127_in =
  _guard5197 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond129_write_en = _guard5198;
assign cond129_clk = clk;
assign cond129_reset = reset;
assign cond129_in =
  _guard5199 ? idx_between_depth_plus_13_depth_plus_14_reg_out :
  1'd0;
assign cond_wire129_in =
  _guard5202 ? cond129_out :
  _guard5203 ? idx_between_depth_plus_13_depth_plus_14_reg_out :
  1'd0;
assign cond_wire136_in =
  _guard5204 ? idx_between_15_depth_plus_15_reg_out :
  _guard5207 ? cond136_out :
  1'd0;
assign cond_wire145_in =
  _guard5208 ? idx_between_10_depth_plus_10_reg_out :
  _guard5211 ? cond145_out :
  1'd0;
assign cond170_write_en = _guard5212;
assign cond170_clk = clk;
assign cond170_reset = reset;
assign cond170_in =
  _guard5213 ? idx_between_depth_plus_16_depth_plus_17_reg_out :
  1'd0;
assign cond_wire184_in =
  _guard5214 ? idx_between_9_min_depth_4_plus_9_reg_out :
  _guard5217 ? cond184_out :
  1'd0;
assign cond_wire194_in =
  _guard5218 ? idx_between_15_depth_plus_15_reg_out :
  _guard5221 ? cond194_out :
  1'd0;
assign cond199_write_en = _guard5222;
assign cond199_clk = clk;
assign cond199_reset = reset;
assign cond199_in =
  _guard5223 ? idx_between_depth_plus_16_depth_plus_17_reg_out :
  1'd0;
assign cond_wire201_in =
  _guard5224 ? idx_between_13_depth_plus_13_reg_out :
  _guard5227 ? cond201_out :
  1'd0;
assign cond211_write_en = _guard5228;
assign cond211_clk = clk;
assign cond211_reset = reset;
assign cond211_in =
  _guard5229 ? idx_between_12_depth_plus_12_reg_out :
  1'd0;
assign cond_wire220_in =
  _guard5232 ? cond220_out :
  _guard5233 ? idx_between_depth_plus_14_depth_plus_15_reg_out :
  1'd0;
assign cond242_write_en = _guard5234;
assign cond242_clk = clk;
assign cond242_reset = reset;
assign cond242_in =
  _guard5235 ? idx_between_9_min_depth_4_plus_9_reg_out :
  1'd0;
assign cond_wire242_in =
  _guard5236 ? idx_between_9_min_depth_4_plus_9_reg_out :
  _guard5239 ? cond242_out :
  1'd0;
assign cond_wire246_in =
  _guard5240 ? idx_between_10_min_depth_4_plus_10_reg_out :
  _guard5243 ? cond246_out :
  1'd0;
assign cond249_write_en = _guard5244;
assign cond249_clk = clk;
assign cond249_reset = reset;
assign cond249_in =
  _guard5245 ? idx_between_depth_plus_14_depth_plus_15_reg_out :
  1'd0;
assign cond_wire249_in =
  _guard5248 ? cond249_out :
  _guard5249 ? idx_between_depth_plus_14_depth_plus_15_reg_out :
  1'd0;
assign cond_wire250_in =
  _guard5250 ? idx_between_11_min_depth_4_plus_11_reg_out :
  _guard5253 ? cond250_out :
  1'd0;
assign cond_wire251_in =
  _guard5254 ? idx_between_11_depth_plus_11_reg_out :
  _guard5257 ? cond251_out :
  1'd0;
assign cond268_write_en = _guard5258;
assign cond268_clk = clk;
assign cond268_reset = reset;
assign cond268_in =
  _guard5259 ? idx_between_depth_plus_19_depth_plus_20_reg_out :
  1'd0;
assign signal_reg_write_en = _guard5269;
assign signal_reg_clk = clk;
assign signal_reg_reset = reset;
assign signal_reg_in =
  _guard5275 ? 1'd1 :
  _guard5278 ? 1'd0 :
  1'd0;
assign depth_plus_17_left = depth;
assign depth_plus_17_right = 32'd17;
assign depth_plus_9_left = depth;
assign depth_plus_9_right = 32'd9;
assign depth_plus_6_left = depth;
assign depth_plus_6_right = 32'd6;
assign top_0_4_write_en = _guard5287;
assign top_0_4_clk = clk;
assign top_0_4_reset = reset;
assign top_0_4_in = t4_read_data;
assign left_0_5_write_en = _guard5293;
assign left_0_5_clk = clk;
assign left_0_5_reset = reset;
assign left_0_5_in = left_0_4_out;
assign pe_2_0_mul_ready =
  _guard5299 ? 1'd1 :
  _guard5302 ? 1'd0 :
  1'd0;
assign pe_2_0_clk = clk;
assign pe_2_0_top =
  _guard5315 ? top_2_0_out :
  32'd0;
assign pe_2_0_left =
  _guard5328 ? left_2_0_out :
  32'd0;
assign pe_2_0_reset = reset;
assign pe_2_0_go = _guard5341;
assign left_2_1_write_en = _guard5344;
assign left_2_1_clk = clk;
assign left_2_1_reset = reset;
assign left_2_1_in = left_2_0_out;
assign top_2_2_write_en = _guard5350;
assign top_2_2_clk = clk;
assign top_2_2_reset = reset;
assign top_2_2_in = top_1_2_out;
assign left_2_5_write_en = _guard5356;
assign left_2_5_clk = clk;
assign left_2_5_reset = reset;
assign left_2_5_in = left_2_4_out;
assign left_3_6_write_en = _guard5362;
assign left_3_6_clk = clk;
assign left_3_6_reset = reset;
assign left_3_6_in = left_3_5_out;
assign pe_4_4_mul_ready =
  _guard5368 ? 1'd1 :
  _guard5371 ? 1'd0 :
  1'd0;
assign pe_4_4_clk = clk;
assign pe_4_4_top =
  _guard5384 ? top_4_4_out :
  32'd0;
assign pe_4_4_left =
  _guard5397 ? left_4_4_out :
  32'd0;
assign pe_4_4_reset = reset;
assign pe_4_4_go = _guard5410;
assign left_4_4_write_en = _guard5413;
assign left_4_4_clk = clk;
assign left_4_4_reset = reset;
assign left_4_4_in = left_4_3_out;
assign pe_4_7_mul_ready =
  _guard5419 ? 1'd1 :
  _guard5422 ? 1'd0 :
  1'd0;
assign pe_4_7_clk = clk;
assign pe_4_7_top =
  _guard5435 ? top_4_7_out :
  32'd0;
assign pe_4_7_left =
  _guard5448 ? left_4_7_out :
  32'd0;
assign pe_4_7_reset = reset;
assign pe_4_7_go = _guard5461;
assign left_5_5_write_en = _guard5464;
assign left_5_5_clk = clk;
assign left_5_5_reset = reset;
assign left_5_5_in = left_5_4_out;
assign left_7_0_write_en = _guard5470;
assign left_7_0_clk = clk;
assign left_7_0_reset = reset;
assign left_7_0_in = l7_read_data;
assign top_7_3_write_en = _guard5476;
assign top_7_3_clk = clk;
assign top_7_3_reset = reset;
assign top_7_3_in = top_6_3_out;
assign top_7_6_write_en = _guard5482;
assign top_7_6_clk = clk;
assign top_7_6_reset = reset;
assign top_7_6_in = top_6_6_out;
assign t1_add_left = 4'd1;
assign t1_add_right = t1_idx_out;
assign t3_idx_write_en = _guard5496;
assign t3_idx_clk = clk;
assign t3_idx_reset = reset;
assign t3_idx_in =
  _guard5499 ? t3_add_out :
  _guard5500 ? 4'd0 :
  'x;
assign l4_add_left = 4'd1;
assign l4_add_right = l4_idx_out;
assign index_ge_2_left = idx_add_out;
assign index_ge_2_right = 32'd2;
assign index_lt_depth_plus_11_left = idx_add_out;
assign index_lt_depth_plus_11_right = depth_plus_11_out;
assign index_lt_depth_plus_7_left = idx_add_out;
assign index_lt_depth_plus_7_right = depth_plus_7_out;
assign index_ge_16_left = idx_add_out;
assign index_ge_16_right = 32'd16;
assign idx_between_16_depth_plus_16_comb_left = index_ge_16_out;
assign idx_between_16_depth_plus_16_comb_right = index_lt_depth_plus_16_out;
assign idx_between_17_depth_plus_17_comb_left = index_ge_17_out;
assign idx_between_17_depth_plus_17_comb_right = index_lt_depth_plus_17_out;
assign idx_between_4_min_depth_4_plus_4_comb_left = index_ge_4_out;
assign idx_between_4_min_depth_4_plus_4_comb_right = index_lt_min_depth_4_plus_4_out;
assign idx_between_5_min_depth_4_plus_5_comb_left = index_ge_5_out;
assign idx_between_5_min_depth_4_plus_5_comb_right = index_lt_min_depth_4_plus_5_out;
assign idx_between_0_depth_plus_0_reg_write_en = _guard5525;
assign idx_between_0_depth_plus_0_reg_clk = clk;
assign idx_between_0_depth_plus_0_reg_reset = reset;
assign idx_between_0_depth_plus_0_reg_in =
  _guard5526 ? 1'd1 :
  _guard5527 ? index_lt_depth_plus_0_out :
  'x;
assign idx_between_10_depth_plus_10_comb_left = index_ge_10_out;
assign idx_between_10_depth_plus_10_comb_right = index_lt_depth_plus_10_out;
assign index_ge_19_left = idx_add_out;
assign index_ge_19_right = 32'd19;
assign idx_between_6_depth_plus_6_reg_write_en = _guard5534;
assign idx_between_6_depth_plus_6_reg_clk = clk;
assign idx_between_6_depth_plus_6_reg_reset = reset;
assign idx_between_6_depth_plus_6_reg_in =
  _guard5535 ? idx_between_6_depth_plus_6_comb_out :
  _guard5536 ? 1'd0 :
  'x;
assign idx_between_depth_plus_7_depth_plus_8_reg_write_en = _guard5539;
assign idx_between_depth_plus_7_depth_plus_8_reg_clk = clk;
assign idx_between_depth_plus_7_depth_plus_8_reg_reset = reset;
assign idx_between_depth_plus_7_depth_plus_8_reg_in =
  _guard5540 ? 1'd0 :
  _guard5541 ? idx_between_depth_plus_7_depth_plus_8_comb_out :
  'x;
assign cond_wire_in =
  _guard5544 ? cond_out :
  _guard5545 ? idx_between_0_depth_plus_0_reg_out :
  1'd0;
assign cond_wire15_in =
  _guard5548 ? cond15_out :
  _guard5549 ? idx_between_4_min_depth_4_plus_4_reg_out :
  1'd0;
assign cond16_write_en = _guard5550;
assign cond16_clk = clk;
assign cond16_reset = reset;
assign cond16_in =
  _guard5551 ? idx_between_4_depth_plus_4_reg_out :
  1'd0;
assign cond37_write_en = _guard5552;
assign cond37_clk = clk;
assign cond37_reset = reset;
assign cond37_in =
  _guard5553 ? idx_between_12_depth_plus_12_reg_out :
  1'd0;
assign cond_wire49_in =
  _guard5554 ? idx_between_4_depth_plus_4_reg_out :
  _guard5557 ? cond49_out :
  1'd0;
assign cond_wire55_in =
  _guard5558 ? idx_between_depth_plus_9_depth_plus_10_reg_out :
  _guard5561 ? cond55_out :
  1'd0;
assign cond_wire93_in =
  _guard5562 ? idx_between_8_min_depth_4_plus_8_reg_out :
  _guard5565 ? cond93_out :
  1'd0;
assign cond_wire95_in =
  _guard5566 ? idx_between_12_depth_plus_12_reg_out :
  _guard5569 ? cond95_out :
  1'd0;
assign cond_wire96_in =
  _guard5572 ? cond96_out :
  _guard5573 ? idx_between_depth_plus_12_depth_plus_13_reg_out :
  1'd0;
assign cond_wire99_in =
  _guard5574 ? idx_between_13_depth_plus_13_reg_out :
  _guard5577 ? cond99_out :
  1'd0;
assign cond110_write_en = _guard5578;
assign cond110_clk = clk;
assign cond110_reset = reset;
assign cond110_in =
  _guard5579 ? idx_between_5_min_depth_4_plus_5_reg_out :
  1'd0;
assign cond113_write_en = _guard5580;
assign cond113_clk = clk;
assign cond113_reset = reset;
assign cond113_in =
  _guard5581 ? idx_between_depth_plus_9_depth_plus_10_reg_out :
  1'd0;
assign cond_wire113_in =
  _guard5582 ? idx_between_depth_plus_9_depth_plus_10_reg_out :
  _guard5585 ? cond113_out :
  1'd0;
assign cond_wire114_in =
  _guard5588 ? cond114_out :
  _guard5589 ? idx_between_6_min_depth_4_plus_6_reg_out :
  1'd0;
assign cond125_write_en = _guard5590;
assign cond125_clk = clk;
assign cond125_reset = reset;
assign cond125_in =
  _guard5591 ? idx_between_depth_plus_12_depth_plus_13_reg_out :
  1'd0;
assign cond130_write_en = _guard5592;
assign cond130_clk = clk;
assign cond130_reset = reset;
assign cond130_in =
  _guard5593 ? idx_between_10_min_depth_4_plus_10_reg_out :
  1'd0;
assign cond_wire133_in =
  _guard5594 ? idx_between_depth_plus_14_depth_plus_15_reg_out :
  _guard5597 ? cond133_out :
  1'd0;
assign cond144_write_en = _guard5598;
assign cond144_clk = clk;
assign cond144_reset = reset;
assign cond144_in =
  _guard5599 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire155_in =
  _guard5600 ? idx_between_9_min_depth_4_plus_9_reg_out :
  _guard5603 ? cond155_out :
  1'd0;
assign cond160_write_en = _guard5604;
assign cond160_clk = clk;
assign cond160_reset = reset;
assign cond160_in =
  _guard5605 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond163_write_en = _guard5606;
assign cond163_clk = clk;
assign cond163_reset = reset;
assign cond163_in =
  _guard5607 ? idx_between_11_min_depth_4_plus_11_reg_out :
  1'd0;
assign cond165_write_en = _guard5608;
assign cond165_clk = clk;
assign cond165_reset = reset;
assign cond165_in =
  _guard5609 ? idx_between_15_depth_plus_15_reg_out :
  1'd0;
assign cond168_write_en = _guard5610;
assign cond168_clk = clk;
assign cond168_reset = reset;
assign cond168_in =
  _guard5611 ? idx_between_12_depth_plus_12_reg_out :
  1'd0;
assign cond_wire173_in =
  _guard5612 ? idx_between_6_depth_plus_6_reg_out :
  _guard5615 ? cond173_out :
  1'd0;
assign cond_wire179_in =
  _guard5618 ? cond179_out :
  _guard5619 ? idx_between_depth_plus_11_depth_plus_12_reg_out :
  1'd0;
assign cond184_write_en = _guard5620;
assign cond184_clk = clk;
assign cond184_reset = reset;
assign cond184_in =
  _guard5621 ? idx_between_9_min_depth_4_plus_9_reg_out :
  1'd0;
assign cond185_write_en = _guard5622;
assign cond185_clk = clk;
assign cond185_reset = reset;
assign cond185_in =
  _guard5623 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond195_write_en = _guard5624;
assign cond195_clk = clk;
assign cond195_reset = reset;
assign cond195_in =
  _guard5625 ? idx_between_depth_plus_15_depth_plus_16_reg_out :
  1'd0;
assign cond197_write_en = _guard5626;
assign cond197_clk = clk;
assign cond197_reset = reset;
assign cond197_in =
  _guard5627 ? idx_between_12_depth_plus_12_reg_out :
  1'd0;
assign cond207_write_en = _guard5628;
assign cond207_clk = clk;
assign cond207_reset = reset;
assign cond207_in =
  _guard5629 ? idx_between_11_depth_plus_11_reg_out :
  1'd0;
assign cond_wire217_in =
  _guard5632 ? cond217_out :
  _guard5633 ? idx_between_10_min_depth_4_plus_10_reg_out :
  1'd0;
assign cond_wire219_in =
  _guard5636 ? cond219_out :
  _guard5637 ? idx_between_14_depth_plus_14_reg_out :
  1'd0;
assign cond_wire241_in =
  _guard5640 ? cond241_out :
  _guard5641 ? idx_between_depth_plus_12_depth_plus_13_reg_out :
  1'd0;
assign cond243_write_en = _guard5642;
assign cond243_clk = clk;
assign cond243_reset = reset;
assign cond243_in =
  _guard5643 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond_wire244_in =
  _guard5644 ? idx_between_13_depth_plus_13_reg_out :
  _guard5647 ? cond244_out :
  1'd0;
assign cond267_write_en = _guard5648;
assign cond267_clk = clk;
assign cond267_reset = reset;
assign cond267_in =
  _guard5649 ? idx_between_19_depth_plus_19_reg_out :
  1'd0;
assign depth_plus_2_left = depth;
assign depth_plus_2_right = 32'd2;
assign depth_plus_19_left = depth;
assign depth_plus_19_right = 32'd19;
assign depth_plus_15_left = depth;
assign depth_plus_15_right = 32'd15;
assign pe_0_0_mul_ready =
  _guard5658 ? 1'd1 :
  _guard5661 ? 1'd0 :
  1'd0;
assign pe_0_0_clk = clk;
assign pe_0_0_top =
  _guard5674 ? top_0_0_out :
  32'd0;
assign pe_0_0_left =
  _guard5687 ? left_0_0_out :
  32'd0;
assign pe_0_0_reset = reset;
assign pe_0_0_go = _guard5700;
assign left_1_6_write_en = _guard5703;
assign left_1_6_clk = clk;
assign left_1_6_reset = reset;
assign left_1_6_in = left_1_5_out;
assign pe_3_3_mul_ready =
  _guard5709 ? 1'd1 :
  _guard5712 ? 1'd0 :
  1'd0;
assign pe_3_3_clk = clk;
assign pe_3_3_top =
  _guard5725 ? top_3_3_out :
  32'd0;
assign pe_3_3_left =
  _guard5738 ? left_3_3_out :
  32'd0;
assign pe_3_3_reset = reset;
assign pe_3_3_go = _guard5751;
assign top_3_3_write_en = _guard5754;
assign top_3_3_clk = clk;
assign top_3_3_reset = reset;
assign top_3_3_in = top_2_3_out;
assign top_4_3_write_en = _guard5760;
assign top_4_3_clk = clk;
assign top_4_3_reset = reset;
assign top_4_3_in = top_3_3_out;
assign top_4_6_write_en = _guard5766;
assign top_4_6_clk = clk;
assign top_4_6_reset = reset;
assign top_4_6_in = top_3_6_out;
assign pe_5_6_mul_ready =
  _guard5772 ? 1'd1 :
  _guard5775 ? 1'd0 :
  1'd0;
assign pe_5_6_clk = clk;
assign pe_5_6_top =
  _guard5788 ? top_5_6_out :
  32'd0;
assign pe_5_6_left =
  _guard5801 ? left_5_6_out :
  32'd0;
assign pe_5_6_reset = reset;
assign pe_5_6_go = _guard5814;
assign top_5_6_write_en = _guard5817;
assign top_5_6_clk = clk;
assign top_5_6_reset = reset;
assign top_5_6_in = top_4_6_out;
assign top_6_2_write_en = _guard5823;
assign top_6_2_clk = clk;
assign top_6_2_reset = reset;
assign top_6_2_in = top_5_2_out;
assign pe_7_1_mul_ready =
  _guard5829 ? 1'd1 :
  _guard5832 ? 1'd0 :
  1'd0;
assign pe_7_1_clk = clk;
assign pe_7_1_top =
  _guard5845 ? top_7_1_out :
  32'd0;
assign pe_7_1_left =
  _guard5858 ? left_7_1_out :
  32'd0;
assign pe_7_1_reset = reset;
assign pe_7_1_go = _guard5871;
assign t2_add_left = 4'd1;
assign t2_add_right = t2_idx_out;
assign t5_add_left = 4'd1;
assign t5_add_right = t5_idx_out;
assign index_lt_depth_plus_13_left = idx_add_out;
assign index_lt_depth_plus_13_right = depth_plus_13_out;
assign idx_between_2_min_depth_4_plus_2_reg_write_en = _guard5888;
assign idx_between_2_min_depth_4_plus_2_reg_clk = clk;
assign idx_between_2_min_depth_4_plus_2_reg_reset = reset;
assign idx_between_2_min_depth_4_plus_2_reg_in =
  _guard5889 ? idx_between_2_min_depth_4_plus_2_comb_out :
  _guard5890 ? 1'd0 :
  'x;
assign idx_between_2_depth_plus_2_reg_write_en = _guard5893;
assign idx_between_2_depth_plus_2_reg_clk = clk;
assign idx_between_2_depth_plus_2_reg_reset = reset;
assign idx_between_2_depth_plus_2_reg_in =
  _guard5894 ? 1'd0 :
  _guard5895 ? idx_between_2_depth_plus_2_comb_out :
  'x;
assign idx_between_2_depth_plus_2_comb_left = index_ge_2_out;
assign idx_between_2_depth_plus_2_comb_right = index_lt_depth_plus_2_out;
assign idx_between_depth_plus_13_depth_plus_14_reg_write_en = _guard5900;
assign idx_between_depth_plus_13_depth_plus_14_reg_clk = clk;
assign idx_between_depth_plus_13_depth_plus_14_reg_reset = reset;
assign idx_between_depth_plus_13_depth_plus_14_reg_in =
  _guard5901 ? idx_between_depth_plus_13_depth_plus_14_comb_out :
  _guard5902 ? 1'd0 :
  'x;
assign idx_between_3_depth_plus_3_reg_write_en = _guard5905;
assign idx_between_3_depth_plus_3_reg_clk = clk;
assign idx_between_3_depth_plus_3_reg_reset = reset;
assign idx_between_3_depth_plus_3_reg_in =
  _guard5906 ? 1'd0 :
  _guard5907 ? idx_between_3_depth_plus_3_comb_out :
  'x;
assign index_lt_depth_plus_12_left = idx_add_out;
assign index_lt_depth_plus_12_right = depth_plus_12_out;
assign idx_between_depth_plus_14_depth_plus_15_reg_write_en = _guard5912;
assign idx_between_depth_plus_14_depth_plus_15_reg_clk = clk;
assign idx_between_depth_plus_14_depth_plus_15_reg_reset = reset;
assign idx_between_depth_plus_14_depth_plus_15_reg_in =
  _guard5913 ? idx_between_depth_plus_14_depth_plus_15_comb_out :
  _guard5914 ? 1'd0 :
  'x;
assign idx_between_depth_plus_9_depth_plus_10_comb_left = index_ge_depth_plus_9_out;
assign idx_between_depth_plus_9_depth_plus_10_comb_right = index_lt_depth_plus_10_out;
assign idx_between_8_depth_plus_8_reg_write_en = _guard5919;
assign idx_between_8_depth_plus_8_reg_clk = clk;
assign idx_between_8_depth_plus_8_reg_reset = reset;
assign idx_between_8_depth_plus_8_reg_in =
  _guard5920 ? 1'd0 :
  _guard5921 ? idx_between_8_depth_plus_8_comb_out :
  'x;
assign index_ge_depth_plus_10_left = idx_add_out;
assign index_ge_depth_plus_10_right = depth_plus_10_out;
assign index_ge_depth_plus_19_left = idx_add_out;
assign index_ge_depth_plus_19_right = depth_plus_19_out;
assign index_lt_min_depth_4_plus_6_left = idx_add_out;
assign index_lt_min_depth_4_plus_6_right = min_depth_4_plus_6_out;
assign index_ge_depth_plus_6_left = idx_add_out;
assign index_ge_depth_plus_6_right = depth_plus_6_out;
assign idx_between_4_depth_plus_4_reg_write_en = _guard5932;
assign idx_between_4_depth_plus_4_reg_clk = clk;
assign idx_between_4_depth_plus_4_reg_reset = reset;
assign idx_between_4_depth_plus_4_reg_in =
  _guard5933 ? idx_between_4_depth_plus_4_comb_out :
  _guard5934 ? 1'd0 :
  'x;
assign index_lt_min_depth_4_plus_4_left = idx_add_out;
assign index_lt_min_depth_4_plus_4_right = min_depth_4_plus_4_out;
assign index_ge_5_left = idx_add_out;
assign index_ge_5_right = 32'd5;
assign idx_between_14_depth_plus_14_reg_write_en = _guard5941;
assign idx_between_14_depth_plus_14_reg_clk = clk;
assign idx_between_14_depth_plus_14_reg_reset = reset;
assign idx_between_14_depth_plus_14_reg_in =
  _guard5942 ? idx_between_14_depth_plus_14_comb_out :
  _guard5943 ? 1'd0 :
  'x;
assign idx_between_10_depth_plus_10_reg_write_en = _guard5946;
assign idx_between_10_depth_plus_10_reg_clk = clk;
assign idx_between_10_depth_plus_10_reg_reset = reset;
assign idx_between_10_depth_plus_10_reg_in =
  _guard5947 ? 1'd0 :
  _guard5948 ? idx_between_10_depth_plus_10_comb_out :
  'x;
assign index_ge_10_left = idx_add_out;
assign index_ge_10_right = 32'd10;
assign idx_between_19_depth_plus_19_comb_left = index_ge_19_out;
assign idx_between_19_depth_plus_19_comb_right = index_lt_depth_plus_19_out;
assign index_lt_min_depth_4_plus_15_left = idx_add_out;
assign index_lt_min_depth_4_plus_15_right = min_depth_4_plus_15_out;
assign cond0_write_en = _guard5955;
assign cond0_clk = clk;
assign cond0_reset = reset;
assign cond0_in =
  _guard5956 ? idx_between_1_min_depth_4_plus_1_reg_out :
  1'd0;
assign cond_wire7_in =
  _guard5959 ? cond7_out :
  _guard5960 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire10_in =
  _guard5961 ? idx_between_3_min_depth_4_plus_3_reg_out :
  _guard5964 ? cond10_out :
  1'd0;
assign cond_wire12_in =
  _guard5965 ? idx_between_7_depth_plus_7_reg_out :
  _guard5968 ? cond12_out :
  1'd0;
assign cond_wire17_in =
  _guard5971 ? cond17_out :
  _guard5972 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire19_in =
  _guard5975 ? cond19_out :
  _guard5976 ? idx_between_4_depth_plus_4_reg_out :
  1'd0;
assign cond_wire23_in =
  _guard5977 ? idx_between_depth_plus_9_depth_plus_10_reg_out :
  _guard5980 ? cond23_out :
  1'd0;
assign cond_wire25_in =
  _guard5981 ? idx_between_6_min_depth_4_plus_6_reg_out :
  _guard5984 ? cond25_out :
  1'd0;
assign cond33_write_en = _guard5985;
assign cond33_clk = clk;
assign cond33_reset = reset;
assign cond33_in =
  _guard5986 ? idx_between_depth_plus_11_depth_plus_12_reg_out :
  1'd0;
assign cond_wire42_in =
  _guard5987 ? idx_between_6_depth_plus_6_reg_out :
  _guard5990 ? cond42_out :
  1'd0;
assign cond47_write_en = _guard5991;
assign cond47_clk = clk;
assign cond47_reset = reset;
assign cond47_in =
  _guard5992 ? idx_between_depth_plus_7_depth_plus_8_reg_out :
  1'd0;
assign cond48_write_en = _guard5993;
assign cond48_clk = clk;
assign cond48_reset = reset;
assign cond48_in =
  _guard5994 ? idx_between_4_min_depth_4_plus_4_reg_out :
  1'd0;
assign cond66_write_en = _guard5995;
assign cond66_clk = clk;
assign cond66_reset = reset;
assign cond66_in =
  _guard5996 ? idx_between_12_depth_plus_12_reg_out :
  1'd0;
assign cond_wire69_in =
  _guard5999 ? cond69_out :
  _guard6000 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond_wire71_in =
  _guard6003 ? cond71_out :
  _guard6004 ? idx_between_depth_plus_13_depth_plus_14_reg_out :
  1'd0;
assign cond82_write_en = _guard6005;
assign cond82_clk = clk;
assign cond82_reset = reset;
assign cond82_in =
  _guard6006 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond84_write_en = _guard6007;
assign cond84_clk = clk;
assign cond84_reset = reset;
assign cond84_in =
  _guard6008 ? idx_between_depth_plus_9_depth_plus_10_reg_out :
  1'd0;
assign cond_wire94_in =
  _guard6011 ? cond94_out :
  _guard6012 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond102_write_en = _guard6013;
assign cond102_clk = clk;
assign cond102_reset = reset;
assign cond102_in =
  _guard6014 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond_wire104_in =
  _guard6015 ? idx_between_depth_plus_14_depth_plus_15_reg_out :
  _guard6018 ? cond104_out :
  1'd0;
assign cond108_write_en = _guard6019;
assign cond108_clk = clk;
assign cond108_reset = reset;
assign cond108_in =
  _guard6020 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire110_in =
  _guard6021 ? idx_between_5_min_depth_4_plus_5_reg_out :
  _guard6024 ? cond110_out :
  1'd0;
assign cond119_write_en = _guard6025;
assign cond119_clk = clk;
assign cond119_reset = reset;
assign cond119_in =
  _guard6026 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond120_write_en = _guard6027;
assign cond120_clk = clk;
assign cond120_reset = reset;
assign cond120_in =
  _guard6028 ? idx_between_11_depth_plus_11_reg_out :
  1'd0;
assign cond_wire130_in =
  _guard6029 ? idx_between_10_min_depth_4_plus_10_reg_out :
  _guard6032 ? cond130_out :
  1'd0;
assign cond_wire135_in =
  _guard6033 ? idx_between_11_depth_plus_11_reg_out :
  _guard6036 ? cond135_out :
  1'd0;
assign cond141_write_en = _guard6037;
assign cond141_clk = clk;
assign cond141_reset = reset;
assign cond141_in =
  _guard6038 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond_wire150_in =
  _guard6041 ? cond150_out :
  _guard6042 ? idx_between_depth_plus_11_depth_plus_12_reg_out :
  1'd0;
assign cond_wire152_in =
  _guard6045 ? cond152_out :
  _guard6046 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire153_in =
  _guard6047 ? idx_between_12_depth_plus_12_reg_out :
  _guard6050 ? cond153_out :
  1'd0;
assign cond210_write_en = _guard6051;
assign cond210_clk = clk;
assign cond210_reset = reset;
assign cond210_in =
  _guard6052 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond218_write_en = _guard6053;
assign cond218_clk = clk;
assign cond218_reset = reset;
assign cond218_in =
  _guard6054 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond229_write_en = _guard6055;
assign cond229_clk = clk;
assign cond229_reset = reset;
assign cond229_in =
  _guard6056 ? idx_between_13_min_depth_4_plus_13_reg_out :
  1'd0;
assign cond_wire255_in =
  _guard6059 ? cond255_out :
  _guard6060 ? idx_between_12_depth_plus_12_reg_out :
  1'd0;
assign cond_wire266_in =
  _guard6061 ? idx_between_15_min_depth_4_plus_15_reg_out :
  _guard6064 ? cond266_out :
  1'd0;
assign tdcc_done_in = _guard6065;
assign top_0_3_write_en = _guard6068;
assign top_0_3_clk = clk;
assign top_0_3_reset = reset;
assign top_0_3_in = t3_read_data;
assign pe_0_6_mul_ready =
  _guard6074 ? 1'd1 :
  _guard6077 ? 1'd0 :
  1'd0;
assign pe_0_6_clk = clk;
assign pe_0_6_top =
  _guard6090 ? top_0_6_out :
  32'd0;
assign pe_0_6_left =
  _guard6103 ? left_0_6_out :
  32'd0;
assign pe_0_6_reset = reset;
assign pe_0_6_go = _guard6116;
assign top_1_7_write_en = _guard6119;
assign top_1_7_clk = clk;
assign top_1_7_reset = reset;
assign top_1_7_in = top_0_7_out;
assign top_2_1_write_en = _guard6125;
assign top_2_1_clk = clk;
assign top_2_1_reset = reset;
assign top_2_1_in = top_1_1_out;
assign left_3_3_write_en = _guard6131;
assign left_3_3_clk = clk;
assign left_3_3_reset = reset;
assign left_3_3_in = left_3_2_out;
assign top_3_7_write_en = _guard6137;
assign top_3_7_clk = clk;
assign top_3_7_reset = reset;
assign top_3_7_in = top_2_7_out;
assign left_4_1_write_en = _guard6143;
assign left_4_1_clk = clk;
assign left_4_1_reset = reset;
assign left_4_1_in = left_4_0_out;
assign pe_4_3_mul_ready =
  _guard6149 ? 1'd1 :
  _guard6152 ? 1'd0 :
  1'd0;
assign pe_4_3_clk = clk;
assign pe_4_3_top =
  _guard6165 ? top_4_3_out :
  32'd0;
assign pe_4_3_left =
  _guard6178 ? left_4_3_out :
  32'd0;
assign pe_4_3_reset = reset;
assign pe_4_3_go = _guard6191;
assign left_5_0_write_en = _guard6194;
assign left_5_0_clk = clk;
assign left_5_0_reset = reset;
assign left_5_0_in = l5_read_data;
assign pe_6_6_mul_ready =
  _guard6200 ? 1'd1 :
  _guard6203 ? 1'd0 :
  1'd0;
assign pe_6_6_clk = clk;
assign pe_6_6_top =
  _guard6216 ? top_6_6_out :
  32'd0;
assign pe_6_6_left =
  _guard6229 ? left_6_6_out :
  32'd0;
assign pe_6_6_reset = reset;
assign pe_6_6_go = _guard6242;
assign pe_7_2_mul_ready =
  _guard6245 ? 1'd1 :
  _guard6248 ? 1'd0 :
  1'd0;
assign pe_7_2_clk = clk;
assign pe_7_2_top =
  _guard6261 ? top_7_2_out :
  32'd0;
assign pe_7_2_left =
  _guard6274 ? left_7_2_out :
  32'd0;
assign pe_7_2_reset = reset;
assign pe_7_2_go = _guard6287;
assign pe_7_7_mul_ready =
  _guard6290 ? 1'd1 :
  _guard6293 ? 1'd0 :
  1'd0;
assign pe_7_7_clk = clk;
assign pe_7_7_top =
  _guard6306 ? top_7_7_out :
  32'd0;
assign pe_7_7_left =
  _guard6319 ? left_7_7_out :
  32'd0;
assign pe_7_7_reset = reset;
assign pe_7_7_go = _guard6332;
assign t2_idx_write_en = _guard6337;
assign t2_idx_clk = clk;
assign t2_idx_reset = reset;
assign t2_idx_in =
  _guard6338 ? 4'd0 :
  _guard6341 ? t2_add_out :
  'x;
assign l2_idx_write_en = _guard6346;
assign l2_idx_clk = clk;
assign l2_idx_reset = reset;
assign l2_idx_in =
  _guard6347 ? 4'd0 :
  _guard6350 ? l2_add_out :
  'x;
assign l6_idx_write_en = _guard6355;
assign l6_idx_clk = clk;
assign l6_idx_reset = reset;
assign l6_idx_in =
  _guard6356 ? 4'd0 :
  _guard6359 ? l6_add_out :
  'x;
assign index_ge_depth_plus_5_left = idx_add_out;
assign index_ge_depth_plus_5_right = depth_plus_5_out;
assign index_ge_depth_plus_14_left = idx_add_out;
assign index_ge_depth_plus_14_right = depth_plus_14_out;
assign index_ge_6_left = idx_add_out;
assign index_ge_6_right = 32'd6;
assign index_ge_depth_plus_15_left = idx_add_out;
assign index_ge_depth_plus_15_right = depth_plus_15_out;
assign index_lt_depth_plus_5_left = idx_add_out;
assign index_lt_depth_plus_5_right = depth_plus_5_out;
assign idx_between_1_depth_plus_1_reg_write_en = _guard6372;
assign idx_between_1_depth_plus_1_reg_clk = clk;
assign idx_between_1_depth_plus_1_reg_reset = reset;
assign idx_between_1_depth_plus_1_reg_in =
  _guard6373 ? idx_between_1_depth_plus_1_comb_out :
  _guard6374 ? 1'd0 :
  'x;
assign cond1_write_en = _guard6375;
assign cond1_clk = clk;
assign cond1_reset = reset;
assign cond1_in =
  _guard6376 ? idx_between_1_depth_plus_1_reg_out :
  1'd0;
assign cond2_write_en = _guard6377;
assign cond2_clk = clk;
assign cond2_reset = reset;
assign cond2_in =
  _guard6378 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond_wire5_in =
  _guard6381 ? cond5_out :
  _guard6382 ? idx_between_2_min_depth_4_plus_2_reg_out :
  1'd0;
assign cond22_write_en = _guard6383;
assign cond22_clk = clk;
assign cond22_reset = reset;
assign cond22_in =
  _guard6384 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond26_write_en = _guard6385;
assign cond26_clk = clk;
assign cond26_reset = reset;
assign cond26_in =
  _guard6386 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire34_in =
  _guard6389 ? cond34_out :
  _guard6390 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond39_write_en = _guard6391;
assign cond39_clk = clk;
assign cond39_reset = reset;
assign cond39_in =
  _guard6392 ? idx_between_1_depth_plus_1_reg_out :
  1'd0;
assign cond49_write_en = _guard6393;
assign cond49_clk = clk;
assign cond49_reset = reset;
assign cond49_in =
  _guard6394 ? idx_between_4_depth_plus_4_reg_out :
  1'd0;
assign cond_wire52_in =
  _guard6397 ? cond52_out :
  _guard6398 ? idx_between_5_min_depth_4_plus_5_reg_out :
  1'd0;
assign cond_wire68_in =
  _guard6401 ? cond68_out :
  _guard6402 ? idx_between_9_min_depth_4_plus_9_reg_out :
  1'd0;
assign cond_wire70_in =
  _guard6405 ? cond70_out :
  _guard6406 ? idx_between_13_depth_plus_13_reg_out :
  1'd0;
assign cond_wire83_in =
  _guard6407 ? idx_between_9_depth_plus_9_reg_out :
  _guard6410 ? cond83_out :
  1'd0;
assign cond87_write_en = _guard6411;
assign cond87_clk = clk;
assign cond87_reset = reset;
assign cond87_in =
  _guard6412 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond96_write_en = _guard6413;
assign cond96_clk = clk;
assign cond96_reset = reset;
assign cond96_in =
  _guard6414 ? idx_between_depth_plus_12_depth_plus_13_reg_out :
  1'd0;
assign cond_wire97_in =
  _guard6415 ? idx_between_9_min_depth_4_plus_9_reg_out :
  _guard6418 ? cond97_out :
  1'd0;
assign cond99_write_en = _guard6419;
assign cond99_clk = clk;
assign cond99_reset = reset;
assign cond99_in =
  _guard6420 ? idx_between_13_depth_plus_13_reg_out :
  1'd0;
assign cond104_write_en = _guard6421;
assign cond104_clk = clk;
assign cond104_reset = reset;
assign cond104_in =
  _guard6422 ? idx_between_depth_plus_14_depth_plus_15_reg_out :
  1'd0;
assign cond133_write_en = _guard6423;
assign cond133_clk = clk;
assign cond133_reset = reset;
assign cond133_in =
  _guard6424 ? idx_between_depth_plus_14_depth_plus_15_reg_out :
  1'd0;
assign cond138_write_en = _guard6425;
assign cond138_clk = clk;
assign cond138_reset = reset;
assign cond138_in =
  _guard6426 ? idx_between_4_depth_plus_4_reg_out :
  1'd0;
assign cond145_write_en = _guard6427;
assign cond145_clk = clk;
assign cond145_reset = reset;
assign cond145_in =
  _guard6428 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond147_write_en = _guard6429;
assign cond147_clk = clk;
assign cond147_reset = reset;
assign cond147_in =
  _guard6430 ? idx_between_7_min_depth_4_plus_7_reg_out :
  1'd0;
assign cond_wire147_in =
  _guard6431 ? idx_between_7_min_depth_4_plus_7_reg_out :
  _guard6434 ? cond147_out :
  1'd0;
assign cond154_write_en = _guard6435;
assign cond154_clk = clk;
assign cond154_reset = reset;
assign cond154_in =
  _guard6436 ? idx_between_depth_plus_12_depth_plus_13_reg_out :
  1'd0;
assign cond156_write_en = _guard6437;
assign cond156_clk = clk;
assign cond156_reset = reset;
assign cond156_in =
  _guard6438 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond_wire168_in =
  _guard6439 ? idx_between_12_depth_plus_12_reg_out :
  _guard6442 ? cond168_out :
  1'd0;
assign cond173_write_en = _guard6443;
assign cond173_clk = clk;
assign cond173_reset = reset;
assign cond173_in =
  _guard6444 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond175_write_en = _guard6445;
assign cond175_clk = clk;
assign cond175_reset = reset;
assign cond175_in =
  _guard6446 ? idx_between_depth_plus_10_depth_plus_11_reg_out :
  1'd0;
assign cond182_write_en = _guard6447;
assign cond182_clk = clk;
assign cond182_reset = reset;
assign cond182_in =
  _guard6448 ? idx_between_12_depth_plus_12_reg_out :
  1'd0;
assign cond_wire199_in =
  _guard6449 ? idx_between_depth_plus_16_depth_plus_17_reg_out :
  _guard6452 ? cond199_out :
  1'd0;
assign cond_wire206_in =
  _guard6455 ? cond206_out :
  _guard6456 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond212_write_en = _guard6457;
assign cond212_clk = clk;
assign cond212_reset = reset;
assign cond212_in =
  _guard6458 ? idx_between_depth_plus_12_depth_plus_13_reg_out :
  1'd0;
assign cond_wire212_in =
  _guard6461 ? cond212_out :
  _guard6462 ? idx_between_depth_plus_12_depth_plus_13_reg_out :
  1'd0;
assign cond224_write_en = _guard6463;
assign cond224_clk = clk;
assign cond224_reset = reset;
assign cond224_in =
  _guard6464 ? idx_between_depth_plus_15_depth_plus_16_reg_out :
  1'd0;
assign cond_wire229_in =
  _guard6465 ? idx_between_13_min_depth_4_plus_13_reg_out :
  _guard6468 ? cond229_out :
  1'd0;
assign cond_wire232_in =
  _guard6471 ? cond232_out :
  _guard6472 ? idx_between_depth_plus_17_depth_plus_18_reg_out :
  1'd0;
assign cond_wire247_in =
  _guard6475 ? cond247_out :
  _guard6476 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond259_write_en = _guard6477;
assign cond259_clk = clk;
assign cond259_reset = reset;
assign cond259_in =
  _guard6478 ? idx_between_13_depth_plus_13_reg_out :
  1'd0;
assign cond_wire259_in =
  _guard6479 ? idx_between_13_depth_plus_13_reg_out :
  _guard6482 ? cond259_out :
  1'd0;
assign cond260_write_en = _guard6483;
assign cond260_clk = clk;
assign cond260_reset = reset;
assign cond260_in =
  _guard6484 ? idx_between_17_depth_plus_17_reg_out :
  1'd0;
assign early_reset_static_par_go_in = _guard6485;
assign iter_limit_write_en = _guard6486;
assign iter_limit_clk = clk;
assign iter_limit_reset = reset;
assign iter_limit_in = depth_plus_16_out;
assign depth_plus_13_left = depth;
assign depth_plus_13_right = 32'd13;
assign depth_plus_11_left = depth;
assign depth_plus_11_right = 32'd11;
assign min_depth_4_plus_7_left = min_depth_4_out;
assign min_depth_4_plus_7_right = 32'd7;
assign min_depth_4_plus_3_left = min_depth_4_out;
assign min_depth_4_plus_3_right = 32'd3;
assign min_depth_4_plus_12_left = min_depth_4_out;
assign min_depth_4_plus_12_right = 32'd12;
assign min_depth_4_plus_1_left = min_depth_4_out;
assign min_depth_4_plus_1_right = 32'd1;
assign top_0_0_write_en = _guard6502;
assign top_0_0_clk = clk;
assign top_0_0_reset = reset;
assign top_0_0_in = t0_read_data;
assign top_0_5_write_en = _guard6508;
assign top_0_5_clk = clk;
assign top_0_5_reset = reset;
assign top_0_5_in = t5_read_data;
assign pe_1_1_mul_ready =
  _guard6514 ? 1'd1 :
  _guard6517 ? 1'd0 :
  1'd0;
assign pe_1_1_clk = clk;
assign pe_1_1_top =
  _guard6530 ? top_1_1_out :
  32'd0;
assign pe_1_1_left =
  _guard6543 ? left_1_1_out :
  32'd0;
assign pe_1_1_reset = reset;
assign pe_1_1_go = _guard6556;
assign top_2_7_write_en = _guard6559;
assign top_2_7_clk = clk;
assign top_2_7_reset = reset;
assign top_2_7_in = top_1_7_out;
assign left_5_2_write_en = _guard6565;
assign left_5_2_clk = clk;
assign left_5_2_reset = reset;
assign left_5_2_in = left_5_1_out;
assign top_5_7_write_en = _guard6571;
assign top_5_7_clk = clk;
assign top_5_7_reset = reset;
assign top_5_7_in = top_4_7_out;
assign left_5_7_write_en = _guard6577;
assign left_5_7_clk = clk;
assign left_5_7_reset = reset;
assign left_5_7_in = left_5_6_out;
assign left_6_0_write_en = _guard6583;
assign left_6_0_clk = clk;
assign left_6_0_reset = reset;
assign left_6_0_in = l6_read_data;
assign top_7_1_write_en = _guard6589;
assign top_7_1_clk = clk;
assign top_7_1_reset = reset;
assign top_7_1_in = top_6_1_out;
assign index_ge_depth_plus_16_left = idx_add_out;
assign index_ge_depth_plus_16_right = depth_plus_16_out;
assign index_lt_depth_plus_2_left = idx_add_out;
assign index_lt_depth_plus_2_right = depth_plus_2_out;
assign idx_between_depth_plus_18_depth_plus_19_reg_write_en = _guard6599;
assign idx_between_depth_plus_18_depth_plus_19_reg_clk = clk;
assign idx_between_depth_plus_18_depth_plus_19_reg_reset = reset;
assign idx_between_depth_plus_18_depth_plus_19_reg_in =
  _guard6600 ? idx_between_depth_plus_18_depth_plus_19_comb_out :
  _guard6601 ? 1'd0 :
  'x;
assign idx_between_depth_plus_5_depth_plus_6_comb_left = index_ge_depth_plus_5_out;
assign idx_between_depth_plus_5_depth_plus_6_comb_right = index_lt_depth_plus_6_out;
assign idx_between_8_depth_plus_8_comb_left = index_ge_8_out;
assign idx_between_8_depth_plus_8_comb_right = index_lt_depth_plus_8_out;
assign idx_between_depth_plus_10_depth_plus_11_comb_left = index_ge_depth_plus_10_out;
assign idx_between_depth_plus_10_depth_plus_11_comb_right = index_lt_depth_plus_11_out;
assign index_ge_13_left = idx_add_out;
assign index_ge_13_right = 32'd13;
assign idx_between_4_min_depth_4_plus_4_reg_write_en = _guard6612;
assign idx_between_4_min_depth_4_plus_4_reg_clk = clk;
assign idx_between_4_min_depth_4_plus_4_reg_reset = reset;
assign idx_between_4_min_depth_4_plus_4_reg_in =
  _guard6613 ? 1'd0 :
  _guard6614 ? idx_between_4_min_depth_4_plus_4_comb_out :
  'x;
assign index_lt_min_depth_4_plus_1_left = idx_add_out;
assign index_lt_min_depth_4_plus_1_right = min_depth_4_plus_1_out;
assign index_lt_min_depth_4_plus_10_left = idx_add_out;
assign index_lt_min_depth_4_plus_10_right = min_depth_4_plus_10_out;
assign idx_between_10_min_depth_4_plus_10_comb_left = index_ge_10_out;
assign idx_between_10_min_depth_4_plus_10_comb_right = index_lt_min_depth_4_plus_10_out;
assign cond_wire1_in =
  _guard6621 ? idx_between_1_depth_plus_1_reg_out :
  _guard6624 ? cond1_out :
  1'd0;
assign cond8_write_en = _guard6625;
assign cond8_clk = clk;
assign cond8_reset = reset;
assign cond8_in =
  _guard6626 ? idx_between_depth_plus_6_depth_plus_7_reg_out :
  1'd0;
assign cond12_write_en = _guard6627;
assign cond12_clk = clk;
assign cond12_reset = reset;
assign cond12_in =
  _guard6628 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond28_write_en = _guard6629;
assign cond28_clk = clk;
assign cond28_reset = reset;
assign cond28_in =
  _guard6630 ? idx_between_depth_plus_10_depth_plus_11_reg_out :
  1'd0;
assign cond_wire28_in =
  _guard6631 ? idx_between_depth_plus_10_depth_plus_11_reg_out :
  _guard6634 ? cond28_out :
  1'd0;
assign cond_wire53_in =
  _guard6637 ? cond53_out :
  _guard6638 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond55_write_en = _guard6639;
assign cond55_clk = clk;
assign cond55_reset = reset;
assign cond55_in =
  _guard6640 ? idx_between_depth_plus_9_depth_plus_10_reg_out :
  1'd0;
assign cond_wire65_in =
  _guard6643 ? cond65_out :
  _guard6644 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond79_write_en = _guard6645;
assign cond79_clk = clk;
assign cond79_reset = reset;
assign cond79_in =
  _guard6646 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire84_in =
  _guard6647 ? idx_between_depth_plus_9_depth_plus_10_reg_out :
  _guard6650 ? cond84_out :
  1'd0;
assign cond_wire88_in =
  _guard6653 ? cond88_out :
  _guard6654 ? idx_between_depth_plus_10_depth_plus_11_reg_out :
  1'd0;
assign cond_wire91_in =
  _guard6655 ? idx_between_11_depth_plus_11_reg_out :
  _guard6658 ? cond91_out :
  1'd0;
assign cond_wire109_in =
  _guard6659 ? idx_between_depth_plus_8_depth_plus_9_reg_out :
  _guard6662 ? cond109_out :
  1'd0;
assign cond_wire115_in =
  _guard6665 ? cond115_out :
  _guard6666 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond117_write_en = _guard6667;
assign cond117_clk = clk;
assign cond117_reset = reset;
assign cond117_in =
  _guard6668 ? idx_between_depth_plus_10_depth_plus_11_reg_out :
  1'd0;
assign cond_wire119_in =
  _guard6669 ? idx_between_7_depth_plus_7_reg_out :
  _guard6672 ? cond119_out :
  1'd0;
assign cond126_write_en = _guard6673;
assign cond126_clk = clk;
assign cond126_reset = reset;
assign cond126_in =
  _guard6674 ? idx_between_9_min_depth_4_plus_9_reg_out :
  1'd0;
assign cond135_write_en = _guard6675;
assign cond135_clk = clk;
assign cond135_reset = reset;
assign cond135_in =
  _guard6676 ? idx_between_11_depth_plus_11_reg_out :
  1'd0;
assign cond_wire141_in =
  _guard6677 ? idx_between_9_depth_plus_9_reg_out :
  _guard6680 ? cond141_out :
  1'd0;
assign cond153_write_en = _guard6681;
assign cond153_clk = clk;
assign cond153_reset = reset;
assign cond153_in =
  _guard6682 ? idx_between_12_depth_plus_12_reg_out :
  1'd0;
assign cond_wire158_in =
  _guard6685 ? cond158_out :
  _guard6686 ? idx_between_depth_plus_13_depth_plus_14_reg_out :
  1'd0;
assign cond_wire159_in =
  _guard6689 ? cond159_out :
  _guard6690 ? idx_between_10_min_depth_4_plus_10_reg_out :
  1'd0;
assign cond_wire169_in =
  _guard6693 ? cond169_out :
  _guard6694 ? idx_between_16_depth_plus_16_reg_out :
  1'd0;
assign cond171_write_en = _guard6695;
assign cond171_clk = clk;
assign cond171_reset = reset;
assign cond171_in =
  _guard6696 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond186_write_en = _guard6697;
assign cond186_clk = clk;
assign cond186_reset = reset;
assign cond186_in =
  _guard6698 ? idx_between_13_depth_plus_13_reg_out :
  1'd0;
assign cond_wire186_in =
  _guard6699 ? idx_between_13_depth_plus_13_reg_out :
  _guard6702 ? cond186_out :
  1'd0;
assign cond_wire196_in =
  _guard6703 ? idx_between_12_min_depth_4_plus_12_reg_out :
  _guard6706 ? cond196_out :
  1'd0;
assign cond213_write_en = _guard6707;
assign cond213_clk = clk;
assign cond213_reset = reset;
assign cond213_in =
  _guard6708 ? idx_between_9_min_depth_4_plus_9_reg_out :
  1'd0;
assign cond234_write_en = _guard6709;
assign cond234_clk = clk;
assign cond234_reset = reset;
assign cond234_in =
  _guard6710 ? idx_between_14_depth_plus_14_reg_out :
  1'd0;
assign cond_wire235_in =
  _guard6711 ? idx_between_18_depth_plus_18_reg_out :
  _guard6714 ? cond235_out :
  1'd0;
assign cond246_write_en = _guard6715;
assign cond246_clk = clk;
assign cond246_reset = reset;
assign cond246_in =
  _guard6716 ? idx_between_10_min_depth_4_plus_10_reg_out :
  1'd0;
assign cond_wire257_in =
  _guard6719 ? cond257_out :
  _guard6720 ? idx_between_depth_plus_16_depth_plus_17_reg_out :
  1'd0;
assign cond261_write_en = _guard6721;
assign cond261_clk = clk;
assign cond261_reset = reset;
assign cond261_in =
  _guard6722 ? idx_between_depth_plus_17_depth_plus_18_reg_out :
  1'd0;
assign min_depth_4_plus_8_left = min_depth_4_out;
assign min_depth_4_plus_8_right = 32'd8;
assign left_0_1_write_en = _guard6727;
assign left_0_1_clk = clk;
assign left_0_1_reset = reset;
assign left_0_1_in = left_0_0_out;
assign top_0_7_write_en = _guard6733;
assign top_0_7_clk = clk;
assign top_0_7_reset = reset;
assign top_0_7_in = t7_read_data;
assign left_1_7_write_en = _guard6739;
assign left_1_7_clk = clk;
assign left_1_7_reset = reset;
assign left_1_7_in = left_1_6_out;
assign pe_2_2_mul_ready =
  _guard6745 ? 1'd1 :
  _guard6748 ? 1'd0 :
  1'd0;
assign pe_2_2_clk = clk;
assign pe_2_2_top =
  _guard6761 ? top_2_2_out :
  32'd0;
assign pe_2_2_left =
  _guard6774 ? left_2_2_out :
  32'd0;
assign pe_2_2_reset = reset;
assign pe_2_2_go = _guard6787;
assign pe_4_1_mul_ready =
  _guard6790 ? 1'd1 :
  _guard6793 ? 1'd0 :
  1'd0;
assign pe_4_1_clk = clk;
assign pe_4_1_top =
  _guard6806 ? top_4_1_out :
  32'd0;
assign pe_4_1_left =
  _guard6819 ? left_4_1_out :
  32'd0;
assign pe_4_1_reset = reset;
assign pe_4_1_go = _guard6832;
assign left_4_3_write_en = _guard6835;
assign left_4_3_clk = clk;
assign left_4_3_reset = reset;
assign left_4_3_in = left_4_2_out;
assign left_6_3_write_en = _guard6841;
assign left_6_3_clk = clk;
assign left_6_3_reset = reset;
assign left_6_3_in = left_6_2_out;
assign l2_add_left = 4'd1;
assign l2_add_right = l2_idx_out;
assign l5_idx_write_en = _guard6855;
assign l5_idx_clk = clk;
assign l5_idx_reset = reset;
assign l5_idx_in =
  _guard6856 ? 4'd0 :
  _guard6859 ? l5_add_out :
  'x;
assign l6_add_left = 4'd1;
assign l6_add_right = l6_idx_out;
assign cond_reg_write_en = _guard6868;
assign cond_reg_clk = clk;
assign cond_reg_reset = reset;
assign cond_reg_in =
  _guard6869 ? 1'd1 :
  _guard6870 ? lt_iter_limit_out :
  'x;
assign idx_between_depth_plus_12_depth_plus_13_reg_write_en = _guard6873;
assign idx_between_depth_plus_12_depth_plus_13_reg_clk = clk;
assign idx_between_depth_plus_12_depth_plus_13_reg_reset = reset;
assign idx_between_depth_plus_12_depth_plus_13_reg_in =
  _guard6874 ? idx_between_depth_plus_12_depth_plus_13_comb_out :
  _guard6875 ? 1'd0 :
  'x;
assign index_ge_depth_plus_8_left = idx_add_out;
assign index_ge_depth_plus_8_right = depth_plus_8_out;
assign index_lt_depth_plus_14_left = idx_add_out;
assign index_lt_depth_plus_14_right = depth_plus_14_out;
assign index_ge_depth_plus_13_left = idx_add_out;
assign index_ge_depth_plus_13_right = depth_plus_13_out;
assign index_lt_depth_plus_16_left = idx_add_out;
assign index_lt_depth_plus_16_right = depth_plus_16_out;
assign idx_between_3_depth_plus_3_comb_left = index_ge_3_out;
assign idx_between_3_depth_plus_3_comb_right = index_lt_depth_plus_3_out;
assign idx_between_13_depth_plus_13_comb_left = index_ge_13_out;
assign idx_between_13_depth_plus_13_comb_right = index_lt_depth_plus_13_out;
assign idx_between_depth_plus_15_depth_plus_16_reg_write_en = _guard6890;
assign idx_between_depth_plus_15_depth_plus_16_reg_clk = clk;
assign idx_between_depth_plus_15_depth_plus_16_reg_reset = reset;
assign idx_between_depth_plus_15_depth_plus_16_reg_in =
  _guard6891 ? idx_between_depth_plus_15_depth_plus_16_comb_out :
  _guard6892 ? 1'd0 :
  'x;
assign idx_between_5_depth_plus_5_reg_write_en = _guard6895;
assign idx_between_5_depth_plus_5_reg_clk = clk;
assign idx_between_5_depth_plus_5_reg_reset = reset;
assign idx_between_5_depth_plus_5_reg_in =
  _guard6896 ? idx_between_5_depth_plus_5_comb_out :
  _guard6897 ? 1'd0 :
  'x;
assign idx_between_14_min_depth_4_plus_14_comb_left = index_ge_14_out;
assign idx_between_14_min_depth_4_plus_14_comb_right = index_lt_min_depth_4_plus_14_out;
assign idx_between_9_depth_plus_9_comb_left = index_ge_9_out;
assign idx_between_9_depth_plus_9_comb_right = index_lt_depth_plus_9_out;
assign index_lt_depth_plus_1_left = idx_add_out;
assign index_lt_depth_plus_1_right = depth_plus_1_out;
assign idx_between_depth_plus_11_depth_plus_12_reg_write_en = _guard6906;
assign idx_between_depth_plus_11_depth_plus_12_reg_clk = clk;
assign idx_between_depth_plus_11_depth_plus_12_reg_reset = reset;
assign idx_between_depth_plus_11_depth_plus_12_reg_in =
  _guard6907 ? idx_between_depth_plus_11_depth_plus_12_comb_out :
  _guard6908 ? 1'd0 :
  'x;
assign cond_wire14_in =
  _guard6911 ? cond14_out :
  _guard6912 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond_wire21_in =
  _guard6915 ? cond21_out :
  _guard6916 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond38_write_en = _guard6917;
assign cond38_clk = clk;
assign cond38_reset = reset;
assign cond38_in =
  _guard6918 ? idx_between_depth_plus_12_depth_plus_13_reg_out :
  1'd0;
assign cond42_write_en = _guard6919;
assign cond42_clk = clk;
assign cond42_reset = reset;
assign cond42_in =
  _guard6920 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire51_in =
  _guard6921 ? idx_between_depth_plus_8_depth_plus_9_reg_out :
  _guard6924 ? cond51_out :
  1'd0;
assign cond59_write_en = _guard6925;
assign cond59_clk = clk;
assign cond59_reset = reset;
assign cond59_in =
  _guard6926 ? idx_between_depth_plus_10_depth_plus_11_reg_out :
  1'd0;
assign cond_wire78_in =
  _guard6929 ? cond78_out :
  _guard6930 ? idx_between_4_depth_plus_4_reg_out :
  1'd0;
assign cond_wire79_in =
  _guard6931 ? idx_between_8_depth_plus_8_reg_out :
  _guard6934 ? cond79_out :
  1'd0;
assign cond85_write_en = _guard6935;
assign cond85_clk = clk;
assign cond85_reset = reset;
assign cond85_in =
  _guard6936 ? idx_between_6_min_depth_4_plus_6_reg_out :
  1'd0;
assign cond_wire102_in =
  _guard6937 ? idx_between_10_depth_plus_10_reg_out :
  _guard6940 ? cond102_out :
  1'd0;
assign cond111_write_en = _guard6941;
assign cond111_clk = clk;
assign cond111_reset = reset;
assign cond111_in =
  _guard6942 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond_wire124_in =
  _guard6943 ? idx_between_12_depth_plus_12_reg_out :
  _guard6946 ? cond124_out :
  1'd0;
assign cond142_write_en = _guard6947;
assign cond142_clk = clk;
assign cond142_reset = reset;
assign cond142_in =
  _guard6948 ? idx_between_depth_plus_9_depth_plus_10_reg_out :
  1'd0;
assign cond157_write_en = _guard6949;
assign cond157_clk = clk;
assign cond157_reset = reset;
assign cond157_in =
  _guard6950 ? idx_between_13_depth_plus_13_reg_out :
  1'd0;
assign cond_wire166_in =
  _guard6953 ? cond166_out :
  _guard6954 ? idx_between_depth_plus_15_depth_plus_16_reg_out :
  1'd0;
assign cond_wire180_in =
  _guard6955 ? idx_between_8_min_depth_4_plus_8_reg_out :
  _guard6958 ? cond180_out :
  1'd0;
assign cond_wire183_in =
  _guard6961 ? cond183_out :
  _guard6962 ? idx_between_depth_plus_12_depth_plus_13_reg_out :
  1'd0;
assign cond_wire188_in =
  _guard6965 ? cond188_out :
  _guard6966 ? idx_between_10_min_depth_4_plus_10_reg_out :
  1'd0;
assign cond200_write_en = _guard6967;
assign cond200_clk = clk;
assign cond200_reset = reset;
assign cond200_in =
  _guard6968 ? idx_between_13_min_depth_4_plus_13_reg_out :
  1'd0;
assign cond_wire202_in =
  _guard6971 ? cond202_out :
  _guard6972 ? idx_between_17_depth_plus_17_reg_out :
  1'd0;
assign cond_wire211_in =
  _guard6973 ? idx_between_12_depth_plus_12_reg_out :
  _guard6976 ? cond211_out :
  1'd0;
assign cond_wire215_in =
  _guard6977 ? idx_between_13_depth_plus_13_reg_out :
  _guard6980 ? cond215_out :
  1'd0;
assign cond_wire226_in =
  _guard6981 ? idx_between_12_depth_plus_12_reg_out :
  _guard6984 ? cond226_out :
  1'd0;
assign cond_wire227_in =
  _guard6987 ? cond227_out :
  _guard6988 ? idx_between_16_depth_plus_16_reg_out :
  1'd0;
assign cond253_write_en = _guard6989;
assign cond253_clk = clk;
assign cond253_reset = reset;
assign cond253_in =
  _guard6990 ? idx_between_depth_plus_15_depth_plus_16_reg_out :
  1'd0;
assign cond254_write_en = _guard6991;
assign cond254_clk = clk;
assign cond254_reset = reset;
assign cond254_in =
  _guard6992 ? idx_between_12_min_depth_4_plus_12_reg_out :
  1'd0;
assign cond_wire254_in =
  _guard6993 ? idx_between_12_min_depth_4_plus_12_reg_out :
  _guard6996 ? cond254_out :
  1'd0;
assign while_wrapper_early_reset_static_par0_go_in = _guard7002;
assign while_wrapper_early_reset_static_par0_done_in = _guard7006;
// COMPONENT END: systolic_array_comp
endmodule
module main(
  input logic go,
  input logic clk,
  input logic reset,
  output logic done,
  output logic [3:0] t0_addr0,
  output logic [31:0] t0_write_data,
  output logic t0_write_en,
  output logic t0_clk,
  output logic t0_reset,
  input logic [31:0] t0_read_data,
  input logic t0_done,
  output logic [3:0] t1_addr0,
  output logic [31:0] t1_write_data,
  output logic t1_write_en,
  output logic t1_clk,
  output logic t1_reset,
  input logic [31:0] t1_read_data,
  input logic t1_done,
  output logic [3:0] t2_addr0,
  output logic [31:0] t2_write_data,
  output logic t2_write_en,
  output logic t2_clk,
  output logic t2_reset,
  input logic [31:0] t2_read_data,
  input logic t2_done,
  output logic [3:0] t3_addr0,
  output logic [31:0] t3_write_data,
  output logic t3_write_en,
  output logic t3_clk,
  output logic t3_reset,
  input logic [31:0] t3_read_data,
  input logic t3_done,
  output logic [3:0] t4_addr0,
  output logic [31:0] t4_write_data,
  output logic t4_write_en,
  output logic t4_clk,
  output logic t4_reset,
  input logic [31:0] t4_read_data,
  input logic t4_done,
  output logic [3:0] t5_addr0,
  output logic [31:0] t5_write_data,
  output logic t5_write_en,
  output logic t5_clk,
  output logic t5_reset,
  input logic [31:0] t5_read_data,
  input logic t5_done,
  output logic [3:0] t6_addr0,
  output logic [31:0] t6_write_data,
  output logic t6_write_en,
  output logic t6_clk,
  output logic t6_reset,
  input logic [31:0] t6_read_data,
  input logic t6_done,
  output logic [3:0] t7_addr0,
  output logic [31:0] t7_write_data,
  output logic t7_write_en,
  output logic t7_clk,
  output logic t7_reset,
  input logic [31:0] t7_read_data,
  input logic t7_done,
  output logic [3:0] l0_addr0,
  output logic [31:0] l0_write_data,
  output logic l0_write_en,
  output logic l0_clk,
  output logic l0_reset,
  input logic [31:0] l0_read_data,
  input logic l0_done,
  output logic [3:0] l1_addr0,
  output logic [31:0] l1_write_data,
  output logic l1_write_en,
  output logic l1_clk,
  output logic l1_reset,
  input logic [31:0] l1_read_data,
  input logic l1_done,
  output logic [3:0] l2_addr0,
  output logic [31:0] l2_write_data,
  output logic l2_write_en,
  output logic l2_clk,
  output logic l2_reset,
  input logic [31:0] l2_read_data,
  input logic l2_done,
  output logic [3:0] l3_addr0,
  output logic [31:0] l3_write_data,
  output logic l3_write_en,
  output logic l3_clk,
  output logic l3_reset,
  input logic [31:0] l3_read_data,
  input logic l3_done,
  output logic [3:0] l4_addr0,
  output logic [31:0] l4_write_data,
  output logic l4_write_en,
  output logic l4_clk,
  output logic l4_reset,
  input logic [31:0] l4_read_data,
  input logic l4_done,
  output logic [3:0] l5_addr0,
  output logic [31:0] l5_write_data,
  output logic l5_write_en,
  output logic l5_clk,
  output logic l5_reset,
  input logic [31:0] l5_read_data,
  input logic l5_done,
  output logic [3:0] l6_addr0,
  output logic [31:0] l6_write_data,
  output logic l6_write_en,
  output logic l6_clk,
  output logic l6_reset,
  input logic [31:0] l6_read_data,
  input logic l6_done,
  output logic [3:0] l7_addr0,
  output logic [31:0] l7_write_data,
  output logic l7_write_en,
  output logic l7_clk,
  output logic l7_reset,
  input logic [31:0] l7_read_data,
  input logic l7_done,
  output logic [31:0] out_mem_0_addr0,
  output logic [31:0] out_mem_0_write_data,
  output logic out_mem_0_write_en,
  output logic out_mem_0_clk,
  output logic out_mem_0_reset,
  input logic [31:0] out_mem_0_read_data,
  input logic out_mem_0_done,
  output logic [31:0] out_mem_1_addr0,
  output logic [31:0] out_mem_1_write_data,
  output logic out_mem_1_write_en,
  output logic out_mem_1_clk,
  output logic out_mem_1_reset,
  input logic [31:0] out_mem_1_read_data,
  input logic out_mem_1_done,
  output logic [31:0] out_mem_2_addr0,
  output logic [31:0] out_mem_2_write_data,
  output logic out_mem_2_write_en,
  output logic out_mem_2_clk,
  output logic out_mem_2_reset,
  input logic [31:0] out_mem_2_read_data,
  input logic out_mem_2_done,
  output logic [31:0] out_mem_3_addr0,
  output logic [31:0] out_mem_3_write_data,
  output logic out_mem_3_write_en,
  output logic out_mem_3_clk,
  output logic out_mem_3_reset,
  input logic [31:0] out_mem_3_read_data,
  input logic out_mem_3_done,
  output logic [31:0] out_mem_4_addr0,
  output logic [31:0] out_mem_4_write_data,
  output logic out_mem_4_write_en,
  output logic out_mem_4_clk,
  output logic out_mem_4_reset,
  input logic [31:0] out_mem_4_read_data,
  input logic out_mem_4_done,
  output logic [31:0] out_mem_5_addr0,
  output logic [31:0] out_mem_5_write_data,
  output logic out_mem_5_write_en,
  output logic out_mem_5_clk,
  output logic out_mem_5_reset,
  input logic [31:0] out_mem_5_read_data,
  input logic out_mem_5_done,
  output logic [31:0] out_mem_6_addr0,
  output logic [31:0] out_mem_6_write_data,
  output logic out_mem_6_write_en,
  output logic out_mem_6_clk,
  output logic out_mem_6_reset,
  input logic [31:0] out_mem_6_read_data,
  input logic out_mem_6_done,
  output logic [31:0] out_mem_7_addr0,
  output logic [31:0] out_mem_7_write_data,
  output logic out_mem_7_write_en,
  output logic out_mem_7_clk,
  output logic out_mem_7_reset,
  input logic [31:0] out_mem_7_read_data,
  input logic out_mem_7_done
);
// COMPONENT START: main
logic [31:0] systolic_array_depth;
logic [31:0] systolic_array_t0_read_data;
logic [31:0] systolic_array_t1_read_data;
logic [31:0] systolic_array_t2_read_data;
logic [31:0] systolic_array_t3_read_data;
logic [31:0] systolic_array_t4_read_data;
logic [31:0] systolic_array_t5_read_data;
logic [31:0] systolic_array_t6_read_data;
logic [31:0] systolic_array_t7_read_data;
logic [31:0] systolic_array_l0_read_data;
logic [31:0] systolic_array_l1_read_data;
logic [31:0] systolic_array_l2_read_data;
logic [31:0] systolic_array_l3_read_data;
logic [31:0] systolic_array_l4_read_data;
logic [31:0] systolic_array_l5_read_data;
logic [31:0] systolic_array_l6_read_data;
logic [31:0] systolic_array_l7_read_data;
logic [3:0] systolic_array_t0_addr0;
logic [3:0] systolic_array_t1_addr0;
logic [3:0] systolic_array_t2_addr0;
logic [3:0] systolic_array_t3_addr0;
logic [3:0] systolic_array_t4_addr0;
logic [3:0] systolic_array_t5_addr0;
logic [3:0] systolic_array_t6_addr0;
logic [3:0] systolic_array_t7_addr0;
logic [3:0] systolic_array_l0_addr0;
logic [3:0] systolic_array_l1_addr0;
logic [3:0] systolic_array_l2_addr0;
logic [3:0] systolic_array_l3_addr0;
logic [3:0] systolic_array_l4_addr0;
logic [3:0] systolic_array_l5_addr0;
logic [3:0] systolic_array_l6_addr0;
logic [3:0] systolic_array_l7_addr0;
logic [31:0] systolic_array_out_mem_0_addr0;
logic [31:0] systolic_array_out_mem_0_write_data;
logic systolic_array_out_mem_0_write_en;
logic [31:0] systolic_array_out_mem_1_addr0;
logic [31:0] systolic_array_out_mem_1_write_data;
logic systolic_array_out_mem_1_write_en;
logic [31:0] systolic_array_out_mem_2_addr0;
logic [31:0] systolic_array_out_mem_2_write_data;
logic systolic_array_out_mem_2_write_en;
logic [31:0] systolic_array_out_mem_3_addr0;
logic [31:0] systolic_array_out_mem_3_write_data;
logic systolic_array_out_mem_3_write_en;
logic [31:0] systolic_array_out_mem_4_addr0;
logic [31:0] systolic_array_out_mem_4_write_data;
logic systolic_array_out_mem_4_write_en;
logic [31:0] systolic_array_out_mem_5_addr0;
logic [31:0] systolic_array_out_mem_5_write_data;
logic systolic_array_out_mem_5_write_en;
logic [31:0] systolic_array_out_mem_6_addr0;
logic [31:0] systolic_array_out_mem_6_write_data;
logic systolic_array_out_mem_6_write_en;
logic [31:0] systolic_array_out_mem_7_addr0;
logic [31:0] systolic_array_out_mem_7_write_data;
logic systolic_array_out_mem_7_write_en;
logic systolic_array_go;
logic systolic_array_clk;
logic systolic_array_reset;
logic systolic_array_done;
logic invoke0_go_in;
logic invoke0_go_out;
logic invoke0_done_in;
logic invoke0_done_out;
systolic_array_comp systolic_array (
    .clk(systolic_array_clk),
    .depth(systolic_array_depth),
    .done(systolic_array_done),
    .go(systolic_array_go),
    .l0_addr0(systolic_array_l0_addr0),
    .l0_read_data(systolic_array_l0_read_data),
    .l1_addr0(systolic_array_l1_addr0),
    .l1_read_data(systolic_array_l1_read_data),
    .l2_addr0(systolic_array_l2_addr0),
    .l2_read_data(systolic_array_l2_read_data),
    .l3_addr0(systolic_array_l3_addr0),
    .l3_read_data(systolic_array_l3_read_data),
    .l4_addr0(systolic_array_l4_addr0),
    .l4_read_data(systolic_array_l4_read_data),
    .l5_addr0(systolic_array_l5_addr0),
    .l5_read_data(systolic_array_l5_read_data),
    .l6_addr0(systolic_array_l6_addr0),
    .l6_read_data(systolic_array_l6_read_data),
    .l7_addr0(systolic_array_l7_addr0),
    .l7_read_data(systolic_array_l7_read_data),
    .out_mem_0_addr0(systolic_array_out_mem_0_addr0),
    .out_mem_0_write_data(systolic_array_out_mem_0_write_data),
    .out_mem_0_write_en(systolic_array_out_mem_0_write_en),
    .out_mem_1_addr0(systolic_array_out_mem_1_addr0),
    .out_mem_1_write_data(systolic_array_out_mem_1_write_data),
    .out_mem_1_write_en(systolic_array_out_mem_1_write_en),
    .out_mem_2_addr0(systolic_array_out_mem_2_addr0),
    .out_mem_2_write_data(systolic_array_out_mem_2_write_data),
    .out_mem_2_write_en(systolic_array_out_mem_2_write_en),
    .out_mem_3_addr0(systolic_array_out_mem_3_addr0),
    .out_mem_3_write_data(systolic_array_out_mem_3_write_data),
    .out_mem_3_write_en(systolic_array_out_mem_3_write_en),
    .out_mem_4_addr0(systolic_array_out_mem_4_addr0),
    .out_mem_4_write_data(systolic_array_out_mem_4_write_data),
    .out_mem_4_write_en(systolic_array_out_mem_4_write_en),
    .out_mem_5_addr0(systolic_array_out_mem_5_addr0),
    .out_mem_5_write_data(systolic_array_out_mem_5_write_data),
    .out_mem_5_write_en(systolic_array_out_mem_5_write_en),
    .out_mem_6_addr0(systolic_array_out_mem_6_addr0),
    .out_mem_6_write_data(systolic_array_out_mem_6_write_data),
    .out_mem_6_write_en(systolic_array_out_mem_6_write_en),
    .out_mem_7_addr0(systolic_array_out_mem_7_addr0),
    .out_mem_7_write_data(systolic_array_out_mem_7_write_data),
    .out_mem_7_write_en(systolic_array_out_mem_7_write_en),
    .reset(systolic_array_reset),
    .t0_addr0(systolic_array_t0_addr0),
    .t0_read_data(systolic_array_t0_read_data),
    .t1_addr0(systolic_array_t1_addr0),
    .t1_read_data(systolic_array_t1_read_data),
    .t2_addr0(systolic_array_t2_addr0),
    .t2_read_data(systolic_array_t2_read_data),
    .t3_addr0(systolic_array_t3_addr0),
    .t3_read_data(systolic_array_t3_read_data),
    .t4_addr0(systolic_array_t4_addr0),
    .t4_read_data(systolic_array_t4_read_data),
    .t5_addr0(systolic_array_t5_addr0),
    .t5_read_data(systolic_array_t5_read_data),
    .t6_addr0(systolic_array_t6_addr0),
    .t6_read_data(systolic_array_t6_read_data),
    .t7_addr0(systolic_array_t7_addr0),
    .t7_read_data(systolic_array_t7_read_data)
);
std_wire # (
    .WIDTH(1)
) invoke0_go (
    .in(invoke0_go_in),
    .out(invoke0_go_out)
);
std_wire # (
    .WIDTH(1)
) invoke0_done (
    .in(invoke0_done_in),
    .out(invoke0_done_out)
);
wire _guard0 = 1;
wire _guard1 = invoke0_go_out;
wire _guard2 = invoke0_go_out;
wire _guard3 = invoke0_done_out;
wire _guard4 = invoke0_go_out;
wire _guard5 = invoke0_go_out;
wire _guard6 = invoke0_go_out;
wire _guard7 = invoke0_go_out;
wire _guard8 = invoke0_go_out;
wire _guard9 = invoke0_go_out;
wire _guard10 = invoke0_go_out;
wire _guard11 = invoke0_go_out;
wire _guard12 = invoke0_go_out;
wire _guard13 = invoke0_go_out;
wire _guard14 = invoke0_go_out;
wire _guard15 = invoke0_go_out;
wire _guard16 = invoke0_go_out;
wire _guard17 = invoke0_go_out;
wire _guard18 = invoke0_go_out;
wire _guard19 = invoke0_go_out;
wire _guard20 = invoke0_go_out;
wire _guard21 = invoke0_go_out;
wire _guard22 = invoke0_go_out;
wire _guard23 = invoke0_go_out;
wire _guard24 = invoke0_go_out;
wire _guard25 = invoke0_go_out;
wire _guard26 = invoke0_go_out;
wire _guard27 = invoke0_go_out;
wire _guard28 = invoke0_go_out;
wire _guard29 = invoke0_go_out;
wire _guard30 = invoke0_go_out;
wire _guard31 = invoke0_go_out;
wire _guard32 = invoke0_go_out;
wire _guard33 = invoke0_go_out;
wire _guard34 = invoke0_go_out;
wire _guard35 = invoke0_go_out;
wire _guard36 = invoke0_go_out;
wire _guard37 = invoke0_go_out;
wire _guard38 = invoke0_go_out;
wire _guard39 = invoke0_go_out;
wire _guard40 = invoke0_go_out;
wire _guard41 = invoke0_go_out;
wire _guard42 = invoke0_go_out;
wire _guard43 = invoke0_go_out;
wire _guard44 = invoke0_go_out;
wire _guard45 = invoke0_go_out;
wire _guard46 = invoke0_go_out;
wire _guard47 = invoke0_go_out;
wire _guard48 = invoke0_go_out;
wire _guard49 = invoke0_go_out;
wire _guard50 = invoke0_go_out;
wire _guard51 = invoke0_go_out;
wire _guard52 = invoke0_go_out;
wire _guard53 = invoke0_go_out;
wire _guard54 = invoke0_go_out;
wire _guard55 = invoke0_go_out;
wire _guard56 = invoke0_go_out;
wire _guard57 = invoke0_go_out;
wire _guard58 = invoke0_go_out;
wire _guard59 = invoke0_go_out;
assign t2_addr0 =
  _guard1 ? systolic_array_t2_addr0 :
  4'd0;
assign out_mem_4_write_data =
  _guard2 ? systolic_array_out_mem_4_write_data :
  32'd0;
assign done = _guard3;
assign t3_reset = reset;
assign l5_addr0 =
  _guard4 ? systolic_array_l5_addr0 :
  4'd0;
assign t0_reset = reset;
assign t6_reset = reset;
assign l5_clk = clk;
assign out_mem_2_reset = reset;
assign l0_addr0 =
  _guard5 ? systolic_array_l0_addr0 :
  4'd0;
assign out_mem_1_addr0 =
  _guard6 ? systolic_array_out_mem_1_addr0 :
  32'd0;
assign out_mem_5_addr0 =
  _guard7 ? systolic_array_out_mem_5_addr0 :
  32'd0;
assign out_mem_5_write_data =
  _guard8 ? systolic_array_out_mem_5_write_data :
  32'd0;
assign t2_clk = clk;
assign l3_clk = clk;
assign out_mem_1_clk = clk;
assign out_mem_3_reset = reset;
assign l6_addr0 =
  _guard9 ? systolic_array_l6_addr0 :
  4'd0;
assign out_mem_0_write_data =
  _guard10 ? systolic_array_out_mem_0_write_data :
  32'd0;
assign out_mem_5_clk = clk;
assign out_mem_6_addr0 =
  _guard11 ? systolic_array_out_mem_6_addr0 :
  32'd0;
assign t5_reset = reset;
assign l7_reset = reset;
assign out_mem_3_write_data =
  _guard12 ? systolic_array_out_mem_3_write_data :
  32'd0;
assign t0_clk = clk;
assign l5_reset = reset;
assign out_mem_1_reset = reset;
assign t5_addr0 =
  _guard13 ? systolic_array_t5_addr0 :
  4'd0;
assign l1_addr0 =
  _guard14 ? systolic_array_l1_addr0 :
  4'd0;
assign out_mem_5_write_en =
  _guard15 ? systolic_array_out_mem_5_write_en :
  1'd0;
assign out_mem_7_addr0 =
  _guard16 ? systolic_array_out_mem_7_addr0 :
  32'd0;
assign t4_reset = reset;
assign t5_clk = clk;
assign t6_clk = clk;
assign l0_reset = reset;
assign l7_clk = clk;
assign out_mem_5_reset = reset;
assign t4_clk = clk;
assign t4_addr0 =
  _guard17 ? systolic_array_t4_addr0 :
  4'd0;
assign t6_addr0 =
  _guard18 ? systolic_array_t6_addr0 :
  4'd0;
assign out_mem_7_write_en =
  _guard19 ? systolic_array_out_mem_7_write_en :
  1'd0;
assign out_mem_0_clk = clk;
assign out_mem_7_clk = clk;
assign out_mem_7_reset = reset;
assign out_mem_4_addr0 =
  _guard20 ? systolic_array_out_mem_4_addr0 :
  32'd0;
assign t1_reset = reset;
assign l6_clk = clk;
assign out_mem_3_clk = clk;
assign out_mem_4_clk = clk;
assign out_mem_4_reset = reset;
assign out_mem_6_reset = reset;
assign l3_addr0 =
  _guard21 ? systolic_array_l3_addr0 :
  4'd0;
assign out_mem_2_write_data =
  _guard22 ? systolic_array_out_mem_2_write_data :
  32'd0;
assign t7_clk = clk;
assign l4_reset = reset;
assign l4_addr0 =
  _guard23 ? systolic_array_l4_addr0 :
  4'd0;
assign l7_addr0 =
  _guard24 ? systolic_array_l7_addr0 :
  4'd0;
assign out_mem_1_write_data =
  _guard25 ? systolic_array_out_mem_1_write_data :
  32'd0;
assign out_mem_1_write_en =
  _guard26 ? systolic_array_out_mem_1_write_en :
  1'd0;
assign out_mem_4_write_en =
  _guard27 ? systolic_array_out_mem_4_write_en :
  1'd0;
assign out_mem_0_reset = reset;
assign out_mem_6_clk = clk;
assign t0_addr0 =
  _guard28 ? systolic_array_t0_addr0 :
  4'd0;
assign t1_addr0 =
  _guard29 ? systolic_array_t1_addr0 :
  4'd0;
assign out_mem_0_write_en =
  _guard30 ? systolic_array_out_mem_0_write_en :
  1'd0;
assign out_mem_2_write_en =
  _guard31 ? systolic_array_out_mem_2_write_en :
  1'd0;
assign t1_clk = clk;
assign l1_reset = reset;
assign l2_clk = clk;
assign l2_reset = reset;
assign out_mem_2_clk = clk;
assign out_mem_3_write_en =
  _guard32 ? systolic_array_out_mem_3_write_en :
  1'd0;
assign out_mem_6_write_data =
  _guard33 ? systolic_array_out_mem_6_write_data :
  32'd0;
assign out_mem_6_write_en =
  _guard34 ? systolic_array_out_mem_6_write_en :
  1'd0;
assign out_mem_7_write_data =
  _guard35 ? systolic_array_out_mem_7_write_data :
  32'd0;
assign t3_clk = clk;
assign t7_reset = reset;
assign l2_addr0 =
  _guard36 ? systolic_array_l2_addr0 :
  4'd0;
assign out_mem_0_addr0 =
  _guard37 ? systolic_array_out_mem_0_addr0 :
  32'd0;
assign out_mem_3_addr0 =
  _guard38 ? systolic_array_out_mem_3_addr0 :
  32'd0;
assign l0_clk = clk;
assign l1_clk = clk;
assign l3_reset = reset;
assign l4_clk = clk;
assign l6_reset = reset;
assign t3_addr0 =
  _guard39 ? systolic_array_t3_addr0 :
  4'd0;
assign t7_addr0 =
  _guard40 ? systolic_array_t7_addr0 :
  4'd0;
assign out_mem_2_addr0 =
  _guard41 ? systolic_array_out_mem_2_addr0 :
  32'd0;
assign t2_reset = reset;
assign invoke0_go_in = go;
assign invoke0_done_in = systolic_array_done;
assign systolic_array_l1_read_data =
  _guard42 ? l1_read_data :
  32'd0;
assign systolic_array_l2_read_data =
  _guard43 ? l2_read_data :
  32'd0;
assign systolic_array_l3_read_data =
  _guard44 ? l3_read_data :
  32'd0;
assign systolic_array_l4_read_data =
  _guard45 ? l4_read_data :
  32'd0;
assign systolic_array_depth =
  _guard46 ? 32'd8 :
  32'd0;
assign systolic_array_t4_read_data =
  _guard47 ? t4_read_data :
  32'd0;
assign systolic_array_l5_read_data =
  _guard48 ? l5_read_data :
  32'd0;
assign systolic_array_l7_read_data =
  _guard49 ? l7_read_data :
  32'd0;
assign systolic_array_clk = clk;
assign systolic_array_t5_read_data =
  _guard50 ? t5_read_data :
  32'd0;
assign systolic_array_t3_read_data =
  _guard51 ? t3_read_data :
  32'd0;
assign systolic_array_l0_read_data =
  _guard52 ? l0_read_data :
  32'd0;
assign systolic_array_l6_read_data =
  _guard53 ? l6_read_data :
  32'd0;
assign systolic_array_reset = reset;
assign systolic_array_go = _guard54;
assign systolic_array_t1_read_data =
  _guard55 ? t1_read_data :
  32'd0;
assign systolic_array_t6_read_data =
  _guard56 ? t6_read_data :
  32'd0;
assign systolic_array_t7_read_data =
  _guard57 ? t7_read_data :
  32'd0;
assign systolic_array_t0_read_data =
  _guard58 ? t0_read_data :
  32'd0;
assign systolic_array_t2_read_data =
  _guard59 ? t2_read_data :
  32'd0;
// COMPONENT END: main
endmodule

