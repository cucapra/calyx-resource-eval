
/// This is mostly used for testing the static guarantees currently.
/// A realistic implementation would probably take four cycles.
module pipelined_mult (
    input wire clk,
    input wire reset,
    // inputs
    input wire [31:0] left,
    input wire [31:0] right,
    // The input has been committed
    output wire [31:0] out
);

logic [31:0] lt, rt, buff0, buff1, buff2, tmp_prod;

assign out = buff2;
assign tmp_prod = lt * rt;

always_ff @(posedge clk) begin
    if (reset) begin
        lt <= 0;
        rt <= 0;
        buff0 <= 0;
        buff1 <= 0;
        buff2 <= 0;
    end else begin
        lt <= left;
        rt <= right;
        buff0 <= tmp_prod;
        buff1 <= buff0;
        buff2 <= buff1;
    end
end

endmodule

module bb_pipelined_mult(
	               input wire [31:0] left,
	               input wire [31:0] right,
	               output wire [31:0] out,
	               input wire clk
	               );
`ifdef __ICARUS__
   reg [31:0] reg0;
   reg [31:0] reg1;
   reg [31:0] reg2;
   reg [31:0] reg3;
   always @( posedge clk ) begin
      reg0 <= left * right;
      reg1 <= reg0;
      reg2 <= reg1;
      reg3 <= reg2;
   end
   assign out = reg3;
`elsif VERILATOR
   reg [31:0] reg0;
   reg [31:0] reg1;
   reg [31:0] reg2;
   reg [31:0] reg3;
   always @( posedge clk ) begin
      reg0 <= left * right;
      reg1 <= reg0;
      reg2 <= reg1;
      reg3 <= reg2;
   end
   assign out = reg3;
`else
   // mul_uint32 is a black box module generated by Xilinx's IP Core generator.
   // Generation commands are in the synth.tcl file.
   mul_uint32 mul_uint32 (
                   .A(left),
                   .B(right),
                   .P(out),
                   .CLK(clk)
                   );
`endif
endmodule
/* verilator lint_off MULTITOP */
/// =================== Unsigned, Fixed Point =========================
module std_fp_add #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  assign out = left + right;
endmodule

module std_fp_sub #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module std_fp_mult_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16,
    parameter SIGNED = 0
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    input  logic             go,
    input  logic             clk,
    input  logic             reset,
    output logic [WIDTH-1:0] out,
    output logic             done
);
  logic [WIDTH-1:0]          rtmp;
  logic [WIDTH-1:0]          ltmp;
  logic [(WIDTH << 1) - 1:0] out_tmp;
  // Buffer used to walk through the 3 cycles of the pipeline.
  logic done_buf[1:0];

  assign done = done_buf[1];

  assign out = out_tmp[(WIDTH << 1) - INT_WIDTH - 1 : WIDTH - INT_WIDTH];

  // If the done buffer is completely empty and go is high then execution
  // just started.
  logic start;
  assign start = go;

  // Start sending the done signal.
  always_ff @(posedge clk) begin
    if (start)
      done_buf[0] <= 1;
    else
      done_buf[0] <= 0;
  end

  // Push the done signal through the pipeline.
  always_ff @(posedge clk) begin
    if (go) begin
      done_buf[1] <= done_buf[0];
    end else begin
      done_buf[1] <= 0;
    end
  end

  // Register the inputs
  always_ff @(posedge clk) begin
    if (reset) begin
      rtmp <= 0;
      ltmp <= 0;
    end else if (go) begin
      if (SIGNED) begin
        rtmp <= $signed(right);
        ltmp <= $signed(left);
      end else begin
        rtmp <= right;
        ltmp <= left;
      end
    end else begin
      rtmp <= 0;
      ltmp <= 0;
    end

  end

  // Compute the output and save it into out_tmp
  always_ff @(posedge clk) begin
    if (reset) begin
      out_tmp <= 0;
    end else if (go) begin
      if (SIGNED) begin
        // In the first cycle, this performs an invalid computation because
        // ltmp and rtmp only get their actual values in cycle 1
        out_tmp <= $signed(
          { {WIDTH{ltmp[WIDTH-1]}}, ltmp} *
          { {WIDTH{rtmp[WIDTH-1]}}, rtmp}
        );
      end else begin
        out_tmp <= ltmp * rtmp;
      end
    end else begin
      out_tmp <= out_tmp;
    end
  end
endmodule

/* verilator lint_off WIDTH */
module std_fp_div_pipe #(
  parameter WIDTH = 32,
  parameter INT_WIDTH = 16,
  parameter FRAC_WIDTH = 16
) (
    input  logic             go,
    input  logic             clk,
    input  logic             reset,
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out_remainder,
    output logic [WIDTH-1:0] out_quotient,
    output logic             done
);
    localparam ITERATIONS = WIDTH + FRAC_WIDTH;

    logic [WIDTH-1:0] quotient, quotient_next;
    logic [WIDTH:0] acc, acc_next;
    logic [$clog2(ITERATIONS)-1:0] idx;
    logic start, running, finished, dividend_is_zero;

    assign start = go && !running;
    assign dividend_is_zero = start && left == 0;
    assign finished = idx == ITERATIONS - 1 && running;

    always_ff @(posedge clk) begin
      if (reset || finished || dividend_is_zero)
        running <= 0;
      else if (start)
        running <= 1;
      else
        running <= running;
    end

    always_comb begin
      if (acc >= {1'b0, right}) begin
        acc_next = acc - right;
        {acc_next, quotient_next} = {acc_next[WIDTH-1:0], quotient, 1'b1};
      end else begin
        {acc_next, quotient_next} = {acc, quotient} << 1;
      end
    end

    // `done` signaling
    always_ff @(posedge clk) begin
      if (dividend_is_zero || finished)
        done <= 1;
      else
        done <= 0;
    end

    always_ff @(posedge clk) begin
      if (running)
        idx <= idx + 1;
      else
        idx <= 0;
    end

    always_ff @(posedge clk) begin
      if (reset) begin
        out_quotient <= 0;
        out_remainder <= 0;
      end else if (start) begin
        out_quotient <= 0;
        out_remainder <= left;
      end else if (go == 0) begin
        out_quotient <= out_quotient;
        out_remainder <= out_remainder;
      end else if (dividend_is_zero) begin
        out_quotient <= 0;
        out_remainder <= 0;
      end else if (finished) begin
        out_quotient <= quotient_next;
        out_remainder <= out_remainder;
      end else begin
        out_quotient <= out_quotient;
        if (right <= out_remainder)
          out_remainder <= out_remainder - right;
        else
          out_remainder <= out_remainder;
      end
    end

    always_ff @(posedge clk) begin
      if (reset) begin
        acc <= 0;
        quotient <= 0;
      end else if (start) begin
        {acc, quotient} <= {{WIDTH{1'b0}}, left, 1'b0};
      end else begin
        acc <= acc_next;
        quotient <= quotient_next;
      end
    end
endmodule

module std_fp_gt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic             out
);
  assign out = left > right;
endmodule

/// =================== Signed, Fixed Point =========================
module std_fp_sadd #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left + right);
endmodule

module std_fp_ssub #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);

  assign out = $signed(left - right);
endmodule

module std_fp_smult_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  [WIDTH-1:0]              left,
    input  [WIDTH-1:0]              right,
    input  logic                    reset,
    input  logic                    go,
    input  logic                    clk,
    output logic [WIDTH-1:0]        out,
    output logic                    done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(INT_WIDTH),
    .FRAC_WIDTH(FRAC_WIDTH),
    .SIGNED(1)
  ) comp (
    .clk(clk),
    .done(done),
    .reset(reset),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

module std_fp_sdiv_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input                     clk,
    input                     go,
    input                     reset,
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out_quotient,
    output signed [WIDTH-1:0] out_remainder,
    output logic              done
);

  logic signed [WIDTH-1:0] left_abs, right_abs, comp_out_q, comp_out_r, right_save, out_rem_intermediate;

  // Registers to figure out how to transform outputs.
  logic different_signs, left_sign, right_sign;

  // Latch the value of control registers so that their available after
  // go signal becomes low.
  always_ff @(posedge clk) begin
    if (go) begin
      right_save <= right_abs;
      left_sign <= left[WIDTH-1];
      right_sign <= right[WIDTH-1];
    end else begin
      left_sign <= left_sign;
      right_save <= right_save;
      right_sign <= right_sign;
    end
  end

  assign right_abs = right[WIDTH-1] ? -right : right;
  assign left_abs = left[WIDTH-1] ? -left : left;

  assign different_signs = left_sign ^ right_sign;
  assign out_quotient = different_signs ? -comp_out_q : comp_out_q;

  // Remainder is computed as:
  //  t0 = |left| % |right|
  //  t1 = if left * right < 0 and t0 != 0 then |right| - t0 else t0
  //  rem = if right < 0 then -t1 else t1
  assign out_rem_intermediate = different_signs & |comp_out_r ? $signed(right_save - comp_out_r) : comp_out_r;
  assign out_remainder = right_sign ? -out_rem_intermediate : out_rem_intermediate;

  std_fp_div_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(INT_WIDTH),
    .FRAC_WIDTH(FRAC_WIDTH)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left_abs),
    .right(right_abs),
    .out_quotient(comp_out_q),
    .out_remainder(comp_out_r)
  );
endmodule

module std_fp_sgt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic signed [WIDTH-1:0] left,
    input  logic signed [WIDTH-1:0] right,
    output logic signed             out
);
  assign out = $signed(left > right);
endmodule

module std_fp_slt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
   input logic signed [WIDTH-1:0] left,
   input logic signed [WIDTH-1:0] right,
   output logic signed            out
);
  assign out = $signed(left < right);
endmodule

/// =================== Unsigned, Bitnum =========================
module std_mult_pipe #(
    parameter WIDTH = 32
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    input  logic             reset,
    input  logic             go,
    input  logic             clk,
    output logic [WIDTH-1:0] out,
    output logic             done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(WIDTH),
    .FRAC_WIDTH(0),
    .SIGNED(0)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

module std_div_pipe #(
    parameter WIDTH = 32
) (
    input                    reset,
    input                    clk,
    input                    go,
    input        [WIDTH-1:0] left,
    input        [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out_remainder,
    output logic [WIDTH-1:0] out_quotient,
    output logic             done
);

  logic [WIDTH-1:0] dividend;
  logic [(WIDTH-1)*2:0] divisor;
  logic [WIDTH-1:0] quotient;
  logic [WIDTH-1:0] quotient_msk;
  logic start, running, finished, dividend_is_zero;

  assign start = go && !running;
  assign finished = quotient_msk == 0 && running;
  assign dividend_is_zero = start && left == 0;

  always_ff @(posedge clk) begin
    // Early return if the divisor is zero.
    if (finished || dividend_is_zero)
      done <= 1;
    else
      done <= 0;
  end

  always_ff @(posedge clk) begin
    if (reset || finished || dividend_is_zero)
      running <= 0;
    else if (start)
      running <= 1;
    else
      running <= running;
  end

  // Outputs
  always_ff @(posedge clk) begin
    if (dividend_is_zero || start) begin
      out_quotient <= 0;
      out_remainder <= 0;
    end else if (finished) begin
      out_quotient <= quotient;
      out_remainder <= dividend;
    end else begin
      // Otherwise, explicitly latch the values.
      out_quotient <= out_quotient;
      out_remainder <= out_remainder;
    end
  end

  // Calculate the quotient mask.
  always_ff @(posedge clk) begin
    if (start)
      quotient_msk <= 1 << WIDTH - 1;
    else if (running)
      quotient_msk <= quotient_msk >> 1;
    else
      quotient_msk <= quotient_msk;
  end

  // Calculate the quotient.
  always_ff @(posedge clk) begin
    if (start)
      quotient <= 0;
    else if (divisor <= dividend)
      quotient <= quotient | quotient_msk;
    else
      quotient <= quotient;
  end

  // Calculate the dividend.
  always_ff @(posedge clk) begin
    if (start)
      dividend <= left;
    else if (divisor <= dividend)
      dividend <= dividend - divisor;
    else
      dividend <= dividend;
  end

  always_ff @(posedge clk) begin
    if (start) begin
      divisor <= right << WIDTH - 1;
    end else if (finished) begin
      divisor <= 0;
    end else begin
      divisor <= divisor >> 1;
    end
  end

  // Simulation self test against unsynthesizable implementation.
  `ifdef VERILATOR
    logic [WIDTH-1:0] l, r;
    always_ff @(posedge clk) begin
      if (go) begin
        l <= left;
        r <= right;
      end else begin
        l <= l;
        r <= r;
      end
    end

    always @(posedge clk) begin
      if (done && $unsigned(out_remainder) != $unsigned(l % r))
        $error(
          "\nstd_div_pipe (Remainder): Computed and golden outputs do not match!\n",
          "left: %0d", $unsigned(l),
          "  right: %0d\n", $unsigned(r),
          "expected: %0d", $unsigned(l % r),
          "  computed: %0d", $unsigned(out_remainder)
        );

      if (done && $unsigned(out_quotient) != $unsigned(l / r))
        $error(
          "\nstd_div_pipe (Quotient): Computed and golden outputs do not match!\n",
          "left: %0d", $unsigned(l),
          "  right: %0d\n", $unsigned(r),
          "expected: %0d", $unsigned(l / r),
          "  computed: %0d", $unsigned(out_quotient)
        );
    end
  `endif
endmodule

/// =================== Signed, Bitnum =========================
module std_sadd #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left + right);
endmodule

module std_ssub #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left - right);
endmodule

module std_smult_pipe #(
    parameter WIDTH = 32
) (
    input  logic                    reset,
    input  logic                    go,
    input  logic                    clk,
    input  signed       [WIDTH-1:0] left,
    input  signed       [WIDTH-1:0] right,
    output logic signed [WIDTH-1:0] out,
    output logic                    done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(WIDTH),
    .FRAC_WIDTH(0),
    .SIGNED(1)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

/* verilator lint_off WIDTH */
module std_sdiv_pipe #(
    parameter WIDTH = 32
) (
    input                           reset,
    input                           clk,
    input                           go,
    input  logic signed [WIDTH-1:0] left,
    input  logic signed [WIDTH-1:0] right,
    output logic signed [WIDTH-1:0] out_quotient,
    output logic signed [WIDTH-1:0] out_remainder,
    output logic                    done
);

  logic signed [WIDTH-1:0] left_abs, right_abs, comp_out_q, comp_out_r, right_save, out_rem_intermediate;

  // Registers to figure out how to transform outputs.
  logic different_signs, left_sign, right_sign;

  // Latch the value of control registers so that their available after
  // go signal becomes low.
  always_ff @(posedge clk) begin
    if (go) begin
      right_save <= right_abs;
      left_sign <= left[WIDTH-1];
      right_sign <= right[WIDTH-1];
    end else begin
      left_sign <= left_sign;
      right_save <= right_save;
      right_sign <= right_sign;
    end
  end

  assign right_abs = right[WIDTH-1] ? -right : right;
  assign left_abs = left[WIDTH-1] ? -left : left;

  assign different_signs = left_sign ^ right_sign;
  assign out_quotient = different_signs ? -comp_out_q : comp_out_q;

  // Remainder is computed as:
  //  t0 = |left| % |right|
  //  t1 = if left * right < 0 and t0 != 0 then |right| - t0 else t0
  //  rem = if right < 0 then -t1 else t1
  assign out_rem_intermediate = different_signs & |comp_out_r ? $signed(right_save - comp_out_r) : comp_out_r;
  assign out_remainder = right_sign ? -out_rem_intermediate : out_rem_intermediate;

  std_div_pipe #(
    .WIDTH(WIDTH)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left_abs),
    .right(right_abs),
    .out_quotient(comp_out_q),
    .out_remainder(comp_out_r)
  );

  // Simulation self test against unsynthesizable implementation.
  `ifdef VERILATOR
    logic signed [WIDTH-1:0] l, r;
    always_ff @(posedge clk) begin
      if (go) begin
        l <= left;
        r <= right;
      end else begin
        l <= l;
        r <= r;
      end
    end

    always @(posedge clk) begin
      if (done && out_quotient != $signed(l / r))
        $error(
          "\nstd_sdiv_pipe (Quotient): Computed and golden outputs do not match!\n",
          "left: %0d", l,
          "  right: %0d\n", r,
          "expected: %0d", $signed(l / r),
          "  computed: %0d", $signed(out_quotient),
        );
      if (done && out_remainder != $signed(((l % r) + r) % r))
        $error(
          "\nstd_sdiv_pipe (Remainder): Computed and golden outputs do not match!\n",
          "left: %0d", l,
          "  right: %0d\n", r,
          "expected: %0d", $signed(((l % r) + r) % r),
          "  computed: %0d", $signed(out_remainder),
        );
    end
  `endif
endmodule

module std_sgt #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left > right);
endmodule

module std_slt #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left < right);
endmodule

module std_seq #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left == right);
endmodule

module std_sneq #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left != right);
endmodule

module std_sge #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left >= right);
endmodule

module std_sle #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left <= right);
endmodule

module std_slsh #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = left <<< right;
endmodule

module std_srsh #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = left >>> right;
endmodule

/**
 * Core primitives for Calyx.
 * Implements core primitives used by the compiler.
 *
 * Conventions:
 * - All parameter names must be SNAKE_CASE and all caps.
 * - Port names must be snake_case, no caps.
 */
`default_nettype none

module std_slice #(
    parameter IN_WIDTH  = 32,
    parameter OUT_WIDTH = 32
) (
   input wire                   logic [ IN_WIDTH-1:0] in,
   output logic [OUT_WIDTH-1:0] out
);
  assign out = in[OUT_WIDTH-1:0];

  `ifdef VERILATOR
    always_comb begin
      if (IN_WIDTH < OUT_WIDTH)
        $error(
          "std_slice: Input width less than output width\n",
          "IN_WIDTH: %0d", IN_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_pad #(
    parameter IN_WIDTH  = 32,
    parameter OUT_WIDTH = 32
) (
   input wire logic [IN_WIDTH-1:0]  in,
   output logic     [OUT_WIDTH-1:0] out
);
  localparam EXTEND = OUT_WIDTH - IN_WIDTH;
  assign out = { {EXTEND {1'b0}}, in};

  `ifdef VERILATOR
    always_comb begin
      if (IN_WIDTH > OUT_WIDTH)
        $error(
          "std_pad: Output width less than input width\n",
          "IN_WIDTH: %0d", IN_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_cat #(
  parameter LEFT_WIDTH  = 32,
  parameter RIGHT_WIDTH = 32,
  parameter OUT_WIDTH = 64
) (
  input wire logic [LEFT_WIDTH-1:0] left,
  input wire logic [RIGHT_WIDTH-1:0] right,
  output logic [OUT_WIDTH-1:0] out
);
  assign out = {left, right};

  `ifdef VERILATOR
    always_comb begin
      if (LEFT_WIDTH + RIGHT_WIDTH != OUT_WIDTH)
        $error(
          "std_cat: Output width must equal sum of input widths\n",
          "LEFT_WIDTH: %0d", LEFT_WIDTH,
          "RIGHT_WIDTH: %0d", RIGHT_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_not #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] in,
   output logic [WIDTH-1:0] out
);
  assign out = ~in;
endmodule

module std_and #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left & right;
endmodule

module std_or #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left | right;
endmodule

module std_xor #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left ^ right;
endmodule

module std_sub #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module std_gt #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left > right;
endmodule

module std_lt #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left < right;
endmodule

module std_eq #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left == right;
endmodule

module std_neq #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left != right;
endmodule

module std_ge #(
    parameter WIDTH = 32
) (
    input wire   logic [WIDTH-1:0] left,
    input wire   logic [WIDTH-1:0] right,
    output logic out
);
  assign out = left >= right;
endmodule

module std_le #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left <= right;
endmodule

module std_lsh #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left << right;
endmodule

module std_rsh #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left >> right;
endmodule

/// this primitive is intended to be used
/// for lowering purposes (not in source programs)
module std_mux #(
    parameter WIDTH = 32
) (
   input wire               logic cond,
   input wire               logic [WIDTH-1:0] tru,
   input wire               logic [WIDTH-1:0] fal,
   output logic [WIDTH-1:0] out
);
  assign out = cond ? tru : fal;
endmodule

module std_mem_d1 #(
    parameter WIDTH = 32,
    parameter SIZE = 16,
    parameter IDX_SIZE = 4
) (
   input wire                logic [IDX_SIZE-1:0] addr0,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  logic [WIDTH-1:0] mem[SIZE-1:0];

  /* verilator lint_off WIDTH */
  assign read_data = mem[addr0];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= SIZE)
        $error(
          "std_mem_d1: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "SIZE: %0d", SIZE
        );
    end
  `endif
endmodule

module std_mem_d2 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0];

  assign read_data = mem[addr0][addr1];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d2: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d2: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
    end
  `endif
endmodule

module std_mem_d3 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D2_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4,
    parameter D2_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [D2_IDX_SIZE-1:0] addr2,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0][D2_SIZE-1:0];

  assign read_data = mem[addr0][addr1][addr2];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1][addr2] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
      if (addr2 >= D2_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr2: %0d\n", addr2,
          "D2_SIZE: %0d", D2_SIZE
        );
    end
  `endif
endmodule

module std_mem_d4 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D2_SIZE = 16,
    parameter D3_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4,
    parameter D2_IDX_SIZE = 4,
    parameter D3_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [D2_IDX_SIZE-1:0] addr2,
   input wire                logic [D3_IDX_SIZE-1:0] addr3,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0][D2_SIZE-1:0][D3_SIZE-1:0];

  assign read_data = mem[addr0][addr1][addr2][addr3];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1][addr2][addr3] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
      if (addr2 >= D2_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr2: %0d\n", addr2,
          "D2_SIZE: %0d", D2_SIZE
        );
      if (addr3 >= D3_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr3: %0d\n", addr3,
          "D3_SIZE: %0d", D3_SIZE
        );
    end
  `endif
endmodule

`default_nettype wire

module undef #(
    parameter WIDTH = 32
) (
   output logic [WIDTH-1:0] out
);
assign out = 'x;
endmodule

module std_const #(
    parameter WIDTH = 32,
    parameter VALUE = 32
) (
   output logic [WIDTH-1:0] out
);
assign out = VALUE;
endmodule

module std_wire #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] in,
   output logic [WIDTH-1:0] out
);
assign out = in;
endmodule

module std_add #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] left,
   input logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
assign out = left + right;
endmodule

module std_reg #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] in,
   input logic write_en,
   input logic clk,
   input logic reset,
   output logic [WIDTH-1:0] out,
   output logic done
);
always_ff @(posedge clk) begin
    if (reset) begin
       out <= 0;
       done <= 0;
    end else if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module mac_pe(
  input logic [31:0] top,
  input logic [31:0] left,
  input logic mul_ready,
  output logic [31:0] out,
  input logic go,
  input logic clk,
  input logic reset,
  output logic done
);
// COMPONENT START: mac_pe
logic [31:0] acc_in;
logic acc_write_en;
logic acc_clk;
logic acc_reset;
logic [31:0] acc_out;
logic acc_done;
logic [31:0] add_left;
logic [31:0] add_right;
logic [31:0] add_out;
logic mul_clk;
logic [31:0] mul_left;
logic [31:0] mul_right;
logic [31:0] mul_out;
logic fsm_in;
logic fsm_write_en;
logic fsm_clk;
logic fsm_reset;
logic fsm_out;
logic fsm_done;
logic ud_out;
logic adder_left;
logic adder_right;
logic adder_out;
logic signal_reg_in;
logic signal_reg_write_en;
logic signal_reg_clk;
logic signal_reg_reset;
logic signal_reg_out;
logic signal_reg_done;
logic early_reset_static_par_go_in;
logic early_reset_static_par_go_out;
logic early_reset_static_par_done_in;
logic early_reset_static_par_done_out;
logic wrapper_early_reset_static_par_go_in;
logic wrapper_early_reset_static_par_go_out;
logic wrapper_early_reset_static_par_done_in;
logic wrapper_early_reset_static_par_done_out;
std_reg # (
    .WIDTH(32)
) acc (
    .clk(acc_clk),
    .done(acc_done),
    .in(acc_in),
    .out(acc_out),
    .reset(acc_reset),
    .write_en(acc_write_en)
);
std_add # (
    .WIDTH(32)
) add (
    .left(add_left),
    .out(add_out),
    .right(add_right)
);
bb_pipelined_mult mul (
    .clk(mul_clk),
    .left(mul_left),
    .out(mul_out),
    .right(mul_right)
);
std_reg # (
    .WIDTH(1)
) fsm (
    .clk(fsm_clk),
    .done(fsm_done),
    .in(fsm_in),
    .out(fsm_out),
    .reset(fsm_reset),
    .write_en(fsm_write_en)
);
undef # (
    .WIDTH(1)
) ud (
    .out(ud_out)
);
std_add # (
    .WIDTH(1)
) adder (
    .left(adder_left),
    .out(adder_out),
    .right(adder_right)
);
std_reg # (
    .WIDTH(1)
) signal_reg (
    .clk(signal_reg_clk),
    .done(signal_reg_done),
    .in(signal_reg_in),
    .out(signal_reg_out),
    .reset(signal_reg_reset),
    .write_en(signal_reg_write_en)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_go (
    .in(early_reset_static_par_go_in),
    .out(early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_done (
    .in(early_reset_static_par_done_in),
    .out(early_reset_static_par_done_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_go (
    .in(wrapper_early_reset_static_par_go_in),
    .out(wrapper_early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_done (
    .in(wrapper_early_reset_static_par_done_in),
    .out(wrapper_early_reset_static_par_done_out)
);
wire _guard0 = 1;
wire _guard1 = early_reset_static_par_go_out;
wire _guard2 = early_reset_static_par_go_out;
wire _guard3 = wrapper_early_reset_static_par_done_out;
wire _guard4 = early_reset_static_par_go_out;
wire _guard5 = fsm_out != 1'd0;
wire _guard6 = early_reset_static_par_go_out;
wire _guard7 = _guard5 & _guard6;
wire _guard8 = fsm_out == 1'd0;
wire _guard9 = early_reset_static_par_go_out;
wire _guard10 = _guard8 & _guard9;
wire _guard11 = early_reset_static_par_go_out;
wire _guard12 = early_reset_static_par_go_out;
wire _guard13 = fsm_out == 1'd0;
wire _guard14 = signal_reg_out;
wire _guard15 = _guard13 & _guard14;
wire _guard16 = fsm_out == 1'd0;
wire _guard17 = signal_reg_out;
wire _guard18 = _guard16 & _guard17;
wire _guard19 = fsm_out == 1'd0;
wire _guard20 = signal_reg_out;
wire _guard21 = ~_guard20;
wire _guard22 = _guard19 & _guard21;
wire _guard23 = wrapper_early_reset_static_par_go_out;
wire _guard24 = _guard22 & _guard23;
wire _guard25 = _guard18 | _guard24;
wire _guard26 = fsm_out == 1'd0;
wire _guard27 = signal_reg_out;
wire _guard28 = ~_guard27;
wire _guard29 = _guard26 & _guard28;
wire _guard30 = wrapper_early_reset_static_par_go_out;
wire _guard31 = _guard29 & _guard30;
wire _guard32 = fsm_out == 1'd0;
wire _guard33 = signal_reg_out;
wire _guard34 = _guard32 & _guard33;
wire _guard35 = early_reset_static_par_go_out;
wire _guard36 = early_reset_static_par_go_out;
wire _guard37 = early_reset_static_par_go_out;
wire _guard38 = early_reset_static_par_go_out;
wire _guard39 = wrapper_early_reset_static_par_go_out;
assign acc_write_en =
  _guard1 ? mul_ready :
  1'd0;
assign acc_clk = clk;
assign acc_reset = reset;
assign acc_in = add_out;
assign done = _guard3;
assign out = acc_out;
assign fsm_write_en = _guard4;
assign fsm_clk = clk;
assign fsm_reset = reset;
assign fsm_in =
  _guard7 ? adder_out :
  _guard10 ? 1'd0 :
  1'd0;
assign adder_left =
  _guard11 ? fsm_out :
  1'd0;
assign adder_right = _guard12;
assign wrapper_early_reset_static_par_go_in = go;
assign wrapper_early_reset_static_par_done_in = _guard15;
assign early_reset_static_par_done_in = ud_out;
assign signal_reg_write_en = _guard25;
assign signal_reg_clk = clk;
assign signal_reg_reset = reset;
assign signal_reg_in =
  _guard31 ? 1'd1 :
  _guard34 ? 1'd0 :
  1'd0;
assign add_left = acc_out;
assign add_right = mul_out;
assign mul_clk = clk;
assign mul_left =
  _guard37 ? top :
  32'd0;
assign mul_right =
  _guard38 ? left :
  32'd0;
assign early_reset_static_par_go_in = _guard39;
// COMPONENT END: mac_pe
endmodule
module systolic_array_comp(
  input logic [31:0] depth,
  input logic [31:0] t0_read_data,
  input logic [31:0] t1_read_data,
  input logic [31:0] t2_read_data,
  input logic [31:0] t3_read_data,
  input logic [31:0] l0_read_data,
  input logic [31:0] l1_read_data,
  input logic [31:0] l2_read_data,
  input logic [31:0] l3_read_data,
  output logic [2:0] t0_addr0,
  output logic [2:0] t1_addr0,
  output logic [2:0] t2_addr0,
  output logic [2:0] t3_addr0,
  output logic [2:0] l0_addr0,
  output logic [2:0] l1_addr0,
  output logic [2:0] l2_addr0,
  output logic [2:0] l3_addr0,
  output logic [31:0] out_mem_0_addr0,
  output logic [31:0] out_mem_0_write_data,
  output logic out_mem_0_write_en,
  output logic [31:0] out_mem_1_addr0,
  output logic [31:0] out_mem_1_write_data,
  output logic out_mem_1_write_en,
  output logic [31:0] out_mem_2_addr0,
  output logic [31:0] out_mem_2_write_data,
  output logic out_mem_2_write_en,
  output logic [31:0] out_mem_3_addr0,
  output logic [31:0] out_mem_3_write_data,
  output logic out_mem_3_write_en,
  input logic go,
  input logic clk,
  input logic reset,
  output logic done
);
// COMPONENT START: systolic_array_comp
logic [31:0] min_depth_4_in;
logic min_depth_4_write_en;
logic min_depth_4_clk;
logic min_depth_4_reset;
logic [31:0] min_depth_4_out;
logic min_depth_4_done;
logic [31:0] iter_limit_in;
logic iter_limit_write_en;
logic iter_limit_clk;
logic iter_limit_reset;
logic [31:0] iter_limit_out;
logic iter_limit_done;
logic [31:0] depth_plus_8_left;
logic [31:0] depth_plus_8_right;
logic [31:0] depth_plus_8_out;
logic [31:0] depth_plus_9_left;
logic [31:0] depth_plus_9_right;
logic [31:0] depth_plus_9_out;
logic [31:0] min_depth_4_plus_2_left;
logic [31:0] min_depth_4_plus_2_right;
logic [31:0] min_depth_4_plus_2_out;
logic [31:0] depth_plus_2_left;
logic [31:0] depth_plus_2_right;
logic [31:0] depth_plus_2_out;
logic [31:0] depth_plus_11_left;
logic [31:0] depth_plus_11_right;
logic [31:0] depth_plus_11_out;
logic [31:0] min_depth_4_plus_7_left;
logic [31:0] min_depth_4_plus_7_right;
logic [31:0] min_depth_4_plus_7_out;
logic [31:0] depth_plus_7_left;
logic [31:0] depth_plus_7_right;
logic [31:0] depth_plus_7_out;
logic [31:0] depth_plus_3_left;
logic [31:0] depth_plus_3_right;
logic [31:0] depth_plus_3_out;
logic [31:0] min_depth_4_plus_3_left;
logic [31:0] min_depth_4_plus_3_right;
logic [31:0] min_depth_4_plus_3_out;
logic [31:0] depth_plus_5_left;
logic [31:0] depth_plus_5_right;
logic [31:0] depth_plus_5_out;
logic [31:0] depth_plus_6_left;
logic [31:0] depth_plus_6_right;
logic [31:0] depth_plus_6_out;
logic [31:0] depth_plus_10_left;
logic [31:0] depth_plus_10_right;
logic [31:0] depth_plus_10_out;
logic [31:0] depth_plus_4_left;
logic [31:0] depth_plus_4_right;
logic [31:0] depth_plus_4_out;
logic [31:0] min_depth_4_plus_4_left;
logic [31:0] min_depth_4_plus_4_right;
logic [31:0] min_depth_4_plus_4_out;
logic [31:0] min_depth_4_plus_5_left;
logic [31:0] min_depth_4_plus_5_right;
logic [31:0] min_depth_4_plus_5_out;
logic [31:0] depth_plus_0_left;
logic [31:0] depth_plus_0_right;
logic [31:0] depth_plus_0_out;
logic [31:0] depth_plus_1_left;
logic [31:0] depth_plus_1_right;
logic [31:0] depth_plus_1_out;
logic [31:0] min_depth_4_plus_1_left;
logic [31:0] min_depth_4_plus_1_right;
logic [31:0] min_depth_4_plus_1_out;
logic [31:0] depth_plus_12_left;
logic [31:0] depth_plus_12_right;
logic [31:0] depth_plus_12_out;
logic [31:0] min_depth_4_plus_6_left;
logic [31:0] min_depth_4_plus_6_right;
logic [31:0] min_depth_4_plus_6_out;
logic [31:0] pe_0_0_top;
logic [31:0] pe_0_0_left;
logic pe_0_0_mul_ready;
logic [31:0] pe_0_0_out;
logic pe_0_0_go;
logic pe_0_0_clk;
logic pe_0_0_reset;
logic pe_0_0_done;
logic [31:0] top_0_0_in;
logic top_0_0_write_en;
logic top_0_0_clk;
logic top_0_0_reset;
logic [31:0] top_0_0_out;
logic top_0_0_done;
logic [31:0] left_0_0_in;
logic left_0_0_write_en;
logic left_0_0_clk;
logic left_0_0_reset;
logic [31:0] left_0_0_out;
logic left_0_0_done;
logic [31:0] pe_0_1_top;
logic [31:0] pe_0_1_left;
logic pe_0_1_mul_ready;
logic [31:0] pe_0_1_out;
logic pe_0_1_go;
logic pe_0_1_clk;
logic pe_0_1_reset;
logic pe_0_1_done;
logic [31:0] top_0_1_in;
logic top_0_1_write_en;
logic top_0_1_clk;
logic top_0_1_reset;
logic [31:0] top_0_1_out;
logic top_0_1_done;
logic [31:0] left_0_1_in;
logic left_0_1_write_en;
logic left_0_1_clk;
logic left_0_1_reset;
logic [31:0] left_0_1_out;
logic left_0_1_done;
logic [31:0] pe_0_2_top;
logic [31:0] pe_0_2_left;
logic pe_0_2_mul_ready;
logic [31:0] pe_0_2_out;
logic pe_0_2_go;
logic pe_0_2_clk;
logic pe_0_2_reset;
logic pe_0_2_done;
logic [31:0] top_0_2_in;
logic top_0_2_write_en;
logic top_0_2_clk;
logic top_0_2_reset;
logic [31:0] top_0_2_out;
logic top_0_2_done;
logic [31:0] left_0_2_in;
logic left_0_2_write_en;
logic left_0_2_clk;
logic left_0_2_reset;
logic [31:0] left_0_2_out;
logic left_0_2_done;
logic [31:0] pe_0_3_top;
logic [31:0] pe_0_3_left;
logic pe_0_3_mul_ready;
logic [31:0] pe_0_3_out;
logic pe_0_3_go;
logic pe_0_3_clk;
logic pe_0_3_reset;
logic pe_0_3_done;
logic [31:0] top_0_3_in;
logic top_0_3_write_en;
logic top_0_3_clk;
logic top_0_3_reset;
logic [31:0] top_0_3_out;
logic top_0_3_done;
logic [31:0] left_0_3_in;
logic left_0_3_write_en;
logic left_0_3_clk;
logic left_0_3_reset;
logic [31:0] left_0_3_out;
logic left_0_3_done;
logic [31:0] pe_1_0_top;
logic [31:0] pe_1_0_left;
logic pe_1_0_mul_ready;
logic [31:0] pe_1_0_out;
logic pe_1_0_go;
logic pe_1_0_clk;
logic pe_1_0_reset;
logic pe_1_0_done;
logic [31:0] top_1_0_in;
logic top_1_0_write_en;
logic top_1_0_clk;
logic top_1_0_reset;
logic [31:0] top_1_0_out;
logic top_1_0_done;
logic [31:0] left_1_0_in;
logic left_1_0_write_en;
logic left_1_0_clk;
logic left_1_0_reset;
logic [31:0] left_1_0_out;
logic left_1_0_done;
logic [31:0] pe_1_1_top;
logic [31:0] pe_1_1_left;
logic pe_1_1_mul_ready;
logic [31:0] pe_1_1_out;
logic pe_1_1_go;
logic pe_1_1_clk;
logic pe_1_1_reset;
logic pe_1_1_done;
logic [31:0] top_1_1_in;
logic top_1_1_write_en;
logic top_1_1_clk;
logic top_1_1_reset;
logic [31:0] top_1_1_out;
logic top_1_1_done;
logic [31:0] left_1_1_in;
logic left_1_1_write_en;
logic left_1_1_clk;
logic left_1_1_reset;
logic [31:0] left_1_1_out;
logic left_1_1_done;
logic [31:0] pe_1_2_top;
logic [31:0] pe_1_2_left;
logic pe_1_2_mul_ready;
logic [31:0] pe_1_2_out;
logic pe_1_2_go;
logic pe_1_2_clk;
logic pe_1_2_reset;
logic pe_1_2_done;
logic [31:0] top_1_2_in;
logic top_1_2_write_en;
logic top_1_2_clk;
logic top_1_2_reset;
logic [31:0] top_1_2_out;
logic top_1_2_done;
logic [31:0] left_1_2_in;
logic left_1_2_write_en;
logic left_1_2_clk;
logic left_1_2_reset;
logic [31:0] left_1_2_out;
logic left_1_2_done;
logic [31:0] pe_1_3_top;
logic [31:0] pe_1_3_left;
logic pe_1_3_mul_ready;
logic [31:0] pe_1_3_out;
logic pe_1_3_go;
logic pe_1_3_clk;
logic pe_1_3_reset;
logic pe_1_3_done;
logic [31:0] top_1_3_in;
logic top_1_3_write_en;
logic top_1_3_clk;
logic top_1_3_reset;
logic [31:0] top_1_3_out;
logic top_1_3_done;
logic [31:0] left_1_3_in;
logic left_1_3_write_en;
logic left_1_3_clk;
logic left_1_3_reset;
logic [31:0] left_1_3_out;
logic left_1_3_done;
logic [31:0] pe_2_0_top;
logic [31:0] pe_2_0_left;
logic pe_2_0_mul_ready;
logic [31:0] pe_2_0_out;
logic pe_2_0_go;
logic pe_2_0_clk;
logic pe_2_0_reset;
logic pe_2_0_done;
logic [31:0] top_2_0_in;
logic top_2_0_write_en;
logic top_2_0_clk;
logic top_2_0_reset;
logic [31:0] top_2_0_out;
logic top_2_0_done;
logic [31:0] left_2_0_in;
logic left_2_0_write_en;
logic left_2_0_clk;
logic left_2_0_reset;
logic [31:0] left_2_0_out;
logic left_2_0_done;
logic [31:0] pe_2_1_top;
logic [31:0] pe_2_1_left;
logic pe_2_1_mul_ready;
logic [31:0] pe_2_1_out;
logic pe_2_1_go;
logic pe_2_1_clk;
logic pe_2_1_reset;
logic pe_2_1_done;
logic [31:0] top_2_1_in;
logic top_2_1_write_en;
logic top_2_1_clk;
logic top_2_1_reset;
logic [31:0] top_2_1_out;
logic top_2_1_done;
logic [31:0] left_2_1_in;
logic left_2_1_write_en;
logic left_2_1_clk;
logic left_2_1_reset;
logic [31:0] left_2_1_out;
logic left_2_1_done;
logic [31:0] pe_2_2_top;
logic [31:0] pe_2_2_left;
logic pe_2_2_mul_ready;
logic [31:0] pe_2_2_out;
logic pe_2_2_go;
logic pe_2_2_clk;
logic pe_2_2_reset;
logic pe_2_2_done;
logic [31:0] top_2_2_in;
logic top_2_2_write_en;
logic top_2_2_clk;
logic top_2_2_reset;
logic [31:0] top_2_2_out;
logic top_2_2_done;
logic [31:0] left_2_2_in;
logic left_2_2_write_en;
logic left_2_2_clk;
logic left_2_2_reset;
logic [31:0] left_2_2_out;
logic left_2_2_done;
logic [31:0] pe_2_3_top;
logic [31:0] pe_2_3_left;
logic pe_2_3_mul_ready;
logic [31:0] pe_2_3_out;
logic pe_2_3_go;
logic pe_2_3_clk;
logic pe_2_3_reset;
logic pe_2_3_done;
logic [31:0] top_2_3_in;
logic top_2_3_write_en;
logic top_2_3_clk;
logic top_2_3_reset;
logic [31:0] top_2_3_out;
logic top_2_3_done;
logic [31:0] left_2_3_in;
logic left_2_3_write_en;
logic left_2_3_clk;
logic left_2_3_reset;
logic [31:0] left_2_3_out;
logic left_2_3_done;
logic [31:0] pe_3_0_top;
logic [31:0] pe_3_0_left;
logic pe_3_0_mul_ready;
logic [31:0] pe_3_0_out;
logic pe_3_0_go;
logic pe_3_0_clk;
logic pe_3_0_reset;
logic pe_3_0_done;
logic [31:0] top_3_0_in;
logic top_3_0_write_en;
logic top_3_0_clk;
logic top_3_0_reset;
logic [31:0] top_3_0_out;
logic top_3_0_done;
logic [31:0] left_3_0_in;
logic left_3_0_write_en;
logic left_3_0_clk;
logic left_3_0_reset;
logic [31:0] left_3_0_out;
logic left_3_0_done;
logic [31:0] pe_3_1_top;
logic [31:0] pe_3_1_left;
logic pe_3_1_mul_ready;
logic [31:0] pe_3_1_out;
logic pe_3_1_go;
logic pe_3_1_clk;
logic pe_3_1_reset;
logic pe_3_1_done;
logic [31:0] top_3_1_in;
logic top_3_1_write_en;
logic top_3_1_clk;
logic top_3_1_reset;
logic [31:0] top_3_1_out;
logic top_3_1_done;
logic [31:0] left_3_1_in;
logic left_3_1_write_en;
logic left_3_1_clk;
logic left_3_1_reset;
logic [31:0] left_3_1_out;
logic left_3_1_done;
logic [31:0] pe_3_2_top;
logic [31:0] pe_3_2_left;
logic pe_3_2_mul_ready;
logic [31:0] pe_3_2_out;
logic pe_3_2_go;
logic pe_3_2_clk;
logic pe_3_2_reset;
logic pe_3_2_done;
logic [31:0] top_3_2_in;
logic top_3_2_write_en;
logic top_3_2_clk;
logic top_3_2_reset;
logic [31:0] top_3_2_out;
logic top_3_2_done;
logic [31:0] left_3_2_in;
logic left_3_2_write_en;
logic left_3_2_clk;
logic left_3_2_reset;
logic [31:0] left_3_2_out;
logic left_3_2_done;
logic [31:0] pe_3_3_top;
logic [31:0] pe_3_3_left;
logic pe_3_3_mul_ready;
logic [31:0] pe_3_3_out;
logic pe_3_3_go;
logic pe_3_3_clk;
logic pe_3_3_reset;
logic pe_3_3_done;
logic [31:0] top_3_3_in;
logic top_3_3_write_en;
logic top_3_3_clk;
logic top_3_3_reset;
logic [31:0] top_3_3_out;
logic top_3_3_done;
logic [31:0] left_3_3_in;
logic left_3_3_write_en;
logic left_3_3_clk;
logic left_3_3_reset;
logic [31:0] left_3_3_out;
logic left_3_3_done;
logic [2:0] t0_idx_in;
logic t0_idx_write_en;
logic t0_idx_clk;
logic t0_idx_reset;
logic [2:0] t0_idx_out;
logic t0_idx_done;
logic [2:0] t0_add_left;
logic [2:0] t0_add_right;
logic [2:0] t0_add_out;
logic [2:0] t1_idx_in;
logic t1_idx_write_en;
logic t1_idx_clk;
logic t1_idx_reset;
logic [2:0] t1_idx_out;
logic t1_idx_done;
logic [2:0] t1_add_left;
logic [2:0] t1_add_right;
logic [2:0] t1_add_out;
logic [2:0] t2_idx_in;
logic t2_idx_write_en;
logic t2_idx_clk;
logic t2_idx_reset;
logic [2:0] t2_idx_out;
logic t2_idx_done;
logic [2:0] t2_add_left;
logic [2:0] t2_add_right;
logic [2:0] t2_add_out;
logic [2:0] t3_idx_in;
logic t3_idx_write_en;
logic t3_idx_clk;
logic t3_idx_reset;
logic [2:0] t3_idx_out;
logic t3_idx_done;
logic [2:0] t3_add_left;
logic [2:0] t3_add_right;
logic [2:0] t3_add_out;
logic [2:0] l0_idx_in;
logic l0_idx_write_en;
logic l0_idx_clk;
logic l0_idx_reset;
logic [2:0] l0_idx_out;
logic l0_idx_done;
logic [2:0] l0_add_left;
logic [2:0] l0_add_right;
logic [2:0] l0_add_out;
logic [2:0] l1_idx_in;
logic l1_idx_write_en;
logic l1_idx_clk;
logic l1_idx_reset;
logic [2:0] l1_idx_out;
logic l1_idx_done;
logic [2:0] l1_add_left;
logic [2:0] l1_add_right;
logic [2:0] l1_add_out;
logic [2:0] l2_idx_in;
logic l2_idx_write_en;
logic l2_idx_clk;
logic l2_idx_reset;
logic [2:0] l2_idx_out;
logic l2_idx_done;
logic [2:0] l2_add_left;
logic [2:0] l2_add_right;
logic [2:0] l2_add_out;
logic [2:0] l3_idx_in;
logic l3_idx_write_en;
logic l3_idx_clk;
logic l3_idx_reset;
logic [2:0] l3_idx_out;
logic l3_idx_done;
logic [2:0] l3_add_left;
logic [2:0] l3_add_right;
logic [2:0] l3_add_out;
logic [31:0] idx_in;
logic idx_write_en;
logic idx_clk;
logic idx_reset;
logic [31:0] idx_out;
logic idx_done;
logic [31:0] idx_add_left;
logic [31:0] idx_add_right;
logic [31:0] idx_add_out;
logic [31:0] lt_iter_limit_left;
logic [31:0] lt_iter_limit_right;
logic lt_iter_limit_out;
logic cond_reg_in;
logic cond_reg_write_en;
logic cond_reg_clk;
logic cond_reg_reset;
logic cond_reg_out;
logic cond_reg_done;
logic idx_between_depth_plus_8_depth_plus_9_reg_in;
logic idx_between_depth_plus_8_depth_plus_9_reg_write_en;
logic idx_between_depth_plus_8_depth_plus_9_reg_clk;
logic idx_between_depth_plus_8_depth_plus_9_reg_reset;
logic idx_between_depth_plus_8_depth_plus_9_reg_out;
logic idx_between_depth_plus_8_depth_plus_9_reg_done;
logic [31:0] index_lt_depth_plus_9_left;
logic [31:0] index_lt_depth_plus_9_right;
logic index_lt_depth_plus_9_out;
logic [31:0] index_ge_depth_plus_8_left;
logic [31:0] index_ge_depth_plus_8_right;
logic index_ge_depth_plus_8_out;
logic idx_between_depth_plus_8_depth_plus_9_comb_left;
logic idx_between_depth_plus_8_depth_plus_9_comb_right;
logic idx_between_depth_plus_8_depth_plus_9_comb_out;
logic idx_between_2_min_depth_4_plus_2_reg_in;
logic idx_between_2_min_depth_4_plus_2_reg_write_en;
logic idx_between_2_min_depth_4_plus_2_reg_clk;
logic idx_between_2_min_depth_4_plus_2_reg_reset;
logic idx_between_2_min_depth_4_plus_2_reg_out;
logic idx_between_2_min_depth_4_plus_2_reg_done;
logic [31:0] index_lt_min_depth_4_plus_2_left;
logic [31:0] index_lt_min_depth_4_plus_2_right;
logic index_lt_min_depth_4_plus_2_out;
logic [31:0] index_ge_2_left;
logic [31:0] index_ge_2_right;
logic index_ge_2_out;
logic idx_between_2_min_depth_4_plus_2_comb_left;
logic idx_between_2_min_depth_4_plus_2_comb_right;
logic idx_between_2_min_depth_4_plus_2_comb_out;
logic idx_between_2_depth_plus_2_reg_in;
logic idx_between_2_depth_plus_2_reg_write_en;
logic idx_between_2_depth_plus_2_reg_clk;
logic idx_between_2_depth_plus_2_reg_reset;
logic idx_between_2_depth_plus_2_reg_out;
logic idx_between_2_depth_plus_2_reg_done;
logic [31:0] index_lt_depth_plus_2_left;
logic [31:0] index_lt_depth_plus_2_right;
logic index_lt_depth_plus_2_out;
logic idx_between_2_depth_plus_2_comb_left;
logic idx_between_2_depth_plus_2_comb_right;
logic idx_between_2_depth_plus_2_comb_out;
logic idx_between_11_depth_plus_11_reg_in;
logic idx_between_11_depth_plus_11_reg_write_en;
logic idx_between_11_depth_plus_11_reg_clk;
logic idx_between_11_depth_plus_11_reg_reset;
logic idx_between_11_depth_plus_11_reg_out;
logic idx_between_11_depth_plus_11_reg_done;
logic [31:0] index_lt_depth_plus_11_left;
logic [31:0] index_lt_depth_plus_11_right;
logic index_lt_depth_plus_11_out;
logic [31:0] index_ge_11_left;
logic [31:0] index_ge_11_right;
logic index_ge_11_out;
logic idx_between_11_depth_plus_11_comb_left;
logic idx_between_11_depth_plus_11_comb_right;
logic idx_between_11_depth_plus_11_comb_out;
logic idx_between_7_min_depth_4_plus_7_reg_in;
logic idx_between_7_min_depth_4_plus_7_reg_write_en;
logic idx_between_7_min_depth_4_plus_7_reg_clk;
logic idx_between_7_min_depth_4_plus_7_reg_reset;
logic idx_between_7_min_depth_4_plus_7_reg_out;
logic idx_between_7_min_depth_4_plus_7_reg_done;
logic [31:0] index_lt_min_depth_4_plus_7_left;
logic [31:0] index_lt_min_depth_4_plus_7_right;
logic index_lt_min_depth_4_plus_7_out;
logic [31:0] index_ge_7_left;
logic [31:0] index_ge_7_right;
logic index_ge_7_out;
logic idx_between_7_min_depth_4_plus_7_comb_left;
logic idx_between_7_min_depth_4_plus_7_comb_right;
logic idx_between_7_min_depth_4_plus_7_comb_out;
logic idx_between_7_depth_plus_7_reg_in;
logic idx_between_7_depth_plus_7_reg_write_en;
logic idx_between_7_depth_plus_7_reg_clk;
logic idx_between_7_depth_plus_7_reg_reset;
logic idx_between_7_depth_plus_7_reg_out;
logic idx_between_7_depth_plus_7_reg_done;
logic [31:0] index_lt_depth_plus_7_left;
logic [31:0] index_lt_depth_plus_7_right;
logic index_lt_depth_plus_7_out;
logic idx_between_7_depth_plus_7_comb_left;
logic idx_between_7_depth_plus_7_comb_right;
logic idx_between_7_depth_plus_7_comb_out;
logic idx_between_3_depth_plus_3_reg_in;
logic idx_between_3_depth_plus_3_reg_write_en;
logic idx_between_3_depth_plus_3_reg_clk;
logic idx_between_3_depth_plus_3_reg_reset;
logic idx_between_3_depth_plus_3_reg_out;
logic idx_between_3_depth_plus_3_reg_done;
logic [31:0] index_lt_depth_plus_3_left;
logic [31:0] index_lt_depth_plus_3_right;
logic index_lt_depth_plus_3_out;
logic [31:0] index_ge_3_left;
logic [31:0] index_ge_3_right;
logic index_ge_3_out;
logic idx_between_3_depth_plus_3_comb_left;
logic idx_between_3_depth_plus_3_comb_right;
logic idx_between_3_depth_plus_3_comb_out;
logic idx_between_3_min_depth_4_plus_3_reg_in;
logic idx_between_3_min_depth_4_plus_3_reg_write_en;
logic idx_between_3_min_depth_4_plus_3_reg_clk;
logic idx_between_3_min_depth_4_plus_3_reg_reset;
logic idx_between_3_min_depth_4_plus_3_reg_out;
logic idx_between_3_min_depth_4_plus_3_reg_done;
logic [31:0] index_lt_min_depth_4_plus_3_left;
logic [31:0] index_lt_min_depth_4_plus_3_right;
logic index_lt_min_depth_4_plus_3_out;
logic idx_between_3_min_depth_4_plus_3_comb_left;
logic idx_between_3_min_depth_4_plus_3_comb_right;
logic idx_between_3_min_depth_4_plus_3_comb_out;
logic idx_between_depth_plus_5_depth_plus_6_reg_in;
logic idx_between_depth_plus_5_depth_plus_6_reg_write_en;
logic idx_between_depth_plus_5_depth_plus_6_reg_clk;
logic idx_between_depth_plus_5_depth_plus_6_reg_reset;
logic idx_between_depth_plus_5_depth_plus_6_reg_out;
logic idx_between_depth_plus_5_depth_plus_6_reg_done;
logic [31:0] index_lt_depth_plus_6_left;
logic [31:0] index_lt_depth_plus_6_right;
logic index_lt_depth_plus_6_out;
logic [31:0] index_ge_depth_plus_5_left;
logic [31:0] index_ge_depth_plus_5_right;
logic index_ge_depth_plus_5_out;
logic idx_between_depth_plus_5_depth_plus_6_comb_left;
logic idx_between_depth_plus_5_depth_plus_6_comb_right;
logic idx_between_depth_plus_5_depth_plus_6_comb_out;
logic idx_between_depth_plus_9_depth_plus_10_reg_in;
logic idx_between_depth_plus_9_depth_plus_10_reg_write_en;
logic idx_between_depth_plus_9_depth_plus_10_reg_clk;
logic idx_between_depth_plus_9_depth_plus_10_reg_reset;
logic idx_between_depth_plus_9_depth_plus_10_reg_out;
logic idx_between_depth_plus_9_depth_plus_10_reg_done;
logic [31:0] index_lt_depth_plus_10_left;
logic [31:0] index_lt_depth_plus_10_right;
logic index_lt_depth_plus_10_out;
logic [31:0] index_ge_depth_plus_9_left;
logic [31:0] index_ge_depth_plus_9_right;
logic index_ge_depth_plus_9_out;
logic idx_between_depth_plus_9_depth_plus_10_comb_left;
logic idx_between_depth_plus_9_depth_plus_10_comb_right;
logic idx_between_depth_plus_9_depth_plus_10_comb_out;
logic idx_between_8_depth_plus_8_reg_in;
logic idx_between_8_depth_plus_8_reg_write_en;
logic idx_between_8_depth_plus_8_reg_clk;
logic idx_between_8_depth_plus_8_reg_reset;
logic idx_between_8_depth_plus_8_reg_out;
logic idx_between_8_depth_plus_8_reg_done;
logic [31:0] index_lt_depth_plus_8_left;
logic [31:0] index_lt_depth_plus_8_right;
logic index_lt_depth_plus_8_out;
logic [31:0] index_ge_8_left;
logic [31:0] index_ge_8_right;
logic index_ge_8_out;
logic idx_between_8_depth_plus_8_comb_left;
logic idx_between_8_depth_plus_8_comb_right;
logic idx_between_8_depth_plus_8_comb_out;
logic idx_between_depth_plus_10_depth_plus_11_reg_in;
logic idx_between_depth_plus_10_depth_plus_11_reg_write_en;
logic idx_between_depth_plus_10_depth_plus_11_reg_clk;
logic idx_between_depth_plus_10_depth_plus_11_reg_reset;
logic idx_between_depth_plus_10_depth_plus_11_reg_out;
logic idx_between_depth_plus_10_depth_plus_11_reg_done;
logic [31:0] index_ge_depth_plus_10_left;
logic [31:0] index_ge_depth_plus_10_right;
logic index_ge_depth_plus_10_out;
logic idx_between_depth_plus_10_depth_plus_11_comb_left;
logic idx_between_depth_plus_10_depth_plus_11_comb_right;
logic idx_between_depth_plus_10_depth_plus_11_comb_out;
logic idx_between_6_depth_plus_6_reg_in;
logic idx_between_6_depth_plus_6_reg_write_en;
logic idx_between_6_depth_plus_6_reg_clk;
logic idx_between_6_depth_plus_6_reg_reset;
logic idx_between_6_depth_plus_6_reg_out;
logic idx_between_6_depth_plus_6_reg_done;
logic [31:0] index_ge_6_left;
logic [31:0] index_ge_6_right;
logic index_ge_6_out;
logic idx_between_6_depth_plus_6_comb_left;
logic idx_between_6_depth_plus_6_comb_right;
logic idx_between_6_depth_plus_6_comb_out;
logic idx_between_depth_plus_6_depth_plus_7_reg_in;
logic idx_between_depth_plus_6_depth_plus_7_reg_write_en;
logic idx_between_depth_plus_6_depth_plus_7_reg_clk;
logic idx_between_depth_plus_6_depth_plus_7_reg_reset;
logic idx_between_depth_plus_6_depth_plus_7_reg_out;
logic idx_between_depth_plus_6_depth_plus_7_reg_done;
logic [31:0] index_ge_depth_plus_6_left;
logic [31:0] index_ge_depth_plus_6_right;
logic index_ge_depth_plus_6_out;
logic idx_between_depth_plus_6_depth_plus_7_comb_left;
logic idx_between_depth_plus_6_depth_plus_7_comb_right;
logic idx_between_depth_plus_6_depth_plus_7_comb_out;
logic idx_between_4_depth_plus_4_reg_in;
logic idx_between_4_depth_plus_4_reg_write_en;
logic idx_between_4_depth_plus_4_reg_clk;
logic idx_between_4_depth_plus_4_reg_reset;
logic idx_between_4_depth_plus_4_reg_out;
logic idx_between_4_depth_plus_4_reg_done;
logic [31:0] index_lt_depth_plus_4_left;
logic [31:0] index_lt_depth_plus_4_right;
logic index_lt_depth_plus_4_out;
logic [31:0] index_ge_4_left;
logic [31:0] index_ge_4_right;
logic index_ge_4_out;
logic idx_between_4_depth_plus_4_comb_left;
logic idx_between_4_depth_plus_4_comb_right;
logic idx_between_4_depth_plus_4_comb_out;
logic idx_between_4_min_depth_4_plus_4_reg_in;
logic idx_between_4_min_depth_4_plus_4_reg_write_en;
logic idx_between_4_min_depth_4_plus_4_reg_clk;
logic idx_between_4_min_depth_4_plus_4_reg_reset;
logic idx_between_4_min_depth_4_plus_4_reg_out;
logic idx_between_4_min_depth_4_plus_4_reg_done;
logic [31:0] index_lt_min_depth_4_plus_4_left;
logic [31:0] index_lt_min_depth_4_plus_4_right;
logic index_lt_min_depth_4_plus_4_out;
logic idx_between_4_min_depth_4_plus_4_comb_left;
logic idx_between_4_min_depth_4_plus_4_comb_right;
logic idx_between_4_min_depth_4_plus_4_comb_out;
logic idx_between_5_depth_plus_5_reg_in;
logic idx_between_5_depth_plus_5_reg_write_en;
logic idx_between_5_depth_plus_5_reg_clk;
logic idx_between_5_depth_plus_5_reg_reset;
logic idx_between_5_depth_plus_5_reg_out;
logic idx_between_5_depth_plus_5_reg_done;
logic [31:0] index_lt_depth_plus_5_left;
logic [31:0] index_lt_depth_plus_5_right;
logic index_lt_depth_plus_5_out;
logic [31:0] index_ge_5_left;
logic [31:0] index_ge_5_right;
logic index_ge_5_out;
logic idx_between_5_depth_plus_5_comb_left;
logic idx_between_5_depth_plus_5_comb_right;
logic idx_between_5_depth_plus_5_comb_out;
logic idx_between_5_min_depth_4_plus_5_reg_in;
logic idx_between_5_min_depth_4_plus_5_reg_write_en;
logic idx_between_5_min_depth_4_plus_5_reg_clk;
logic idx_between_5_min_depth_4_plus_5_reg_reset;
logic idx_between_5_min_depth_4_plus_5_reg_out;
logic idx_between_5_min_depth_4_plus_5_reg_done;
logic [31:0] index_lt_min_depth_4_plus_5_left;
logic [31:0] index_lt_min_depth_4_plus_5_right;
logic index_lt_min_depth_4_plus_5_out;
logic idx_between_5_min_depth_4_plus_5_comb_left;
logic idx_between_5_min_depth_4_plus_5_comb_right;
logic idx_between_5_min_depth_4_plus_5_comb_out;
logic idx_between_0_depth_plus_0_reg_in;
logic idx_between_0_depth_plus_0_reg_write_en;
logic idx_between_0_depth_plus_0_reg_clk;
logic idx_between_0_depth_plus_0_reg_reset;
logic idx_between_0_depth_plus_0_reg_out;
logic idx_between_0_depth_plus_0_reg_done;
logic [31:0] index_lt_depth_plus_0_left;
logic [31:0] index_lt_depth_plus_0_right;
logic index_lt_depth_plus_0_out;
logic idx_between_9_depth_plus_9_reg_in;
logic idx_between_9_depth_plus_9_reg_write_en;
logic idx_between_9_depth_plus_9_reg_clk;
logic idx_between_9_depth_plus_9_reg_reset;
logic idx_between_9_depth_plus_9_reg_out;
logic idx_between_9_depth_plus_9_reg_done;
logic [31:0] index_ge_9_left;
logic [31:0] index_ge_9_right;
logic index_ge_9_out;
logic idx_between_9_depth_plus_9_comb_left;
logic idx_between_9_depth_plus_9_comb_right;
logic idx_between_9_depth_plus_9_comb_out;
logic idx_between_1_depth_plus_1_reg_in;
logic idx_between_1_depth_plus_1_reg_write_en;
logic idx_between_1_depth_plus_1_reg_clk;
logic idx_between_1_depth_plus_1_reg_reset;
logic idx_between_1_depth_plus_1_reg_out;
logic idx_between_1_depth_plus_1_reg_done;
logic [31:0] index_lt_depth_plus_1_left;
logic [31:0] index_lt_depth_plus_1_right;
logic index_lt_depth_plus_1_out;
logic [31:0] index_ge_1_left;
logic [31:0] index_ge_1_right;
logic index_ge_1_out;
logic idx_between_1_depth_plus_1_comb_left;
logic idx_between_1_depth_plus_1_comb_right;
logic idx_between_1_depth_plus_1_comb_out;
logic idx_between_1_min_depth_4_plus_1_reg_in;
logic idx_between_1_min_depth_4_plus_1_reg_write_en;
logic idx_between_1_min_depth_4_plus_1_reg_clk;
logic idx_between_1_min_depth_4_plus_1_reg_reset;
logic idx_between_1_min_depth_4_plus_1_reg_out;
logic idx_between_1_min_depth_4_plus_1_reg_done;
logic [31:0] index_lt_min_depth_4_plus_1_left;
logic [31:0] index_lt_min_depth_4_plus_1_right;
logic index_lt_min_depth_4_plus_1_out;
logic idx_between_1_min_depth_4_plus_1_comb_left;
logic idx_between_1_min_depth_4_plus_1_comb_right;
logic idx_between_1_min_depth_4_plus_1_comb_out;
logic idx_between_depth_plus_11_depth_plus_12_reg_in;
logic idx_between_depth_plus_11_depth_plus_12_reg_write_en;
logic idx_between_depth_plus_11_depth_plus_12_reg_clk;
logic idx_between_depth_plus_11_depth_plus_12_reg_reset;
logic idx_between_depth_plus_11_depth_plus_12_reg_out;
logic idx_between_depth_plus_11_depth_plus_12_reg_done;
logic [31:0] index_lt_depth_plus_12_left;
logic [31:0] index_lt_depth_plus_12_right;
logic index_lt_depth_plus_12_out;
logic [31:0] index_ge_depth_plus_11_left;
logic [31:0] index_ge_depth_plus_11_right;
logic index_ge_depth_plus_11_out;
logic idx_between_depth_plus_11_depth_plus_12_comb_left;
logic idx_between_depth_plus_11_depth_plus_12_comb_right;
logic idx_between_depth_plus_11_depth_plus_12_comb_out;
logic idx_between_10_depth_plus_10_reg_in;
logic idx_between_10_depth_plus_10_reg_write_en;
logic idx_between_10_depth_plus_10_reg_clk;
logic idx_between_10_depth_plus_10_reg_reset;
logic idx_between_10_depth_plus_10_reg_out;
logic idx_between_10_depth_plus_10_reg_done;
logic [31:0] index_ge_10_left;
logic [31:0] index_ge_10_right;
logic index_ge_10_out;
logic idx_between_10_depth_plus_10_comb_left;
logic idx_between_10_depth_plus_10_comb_right;
logic idx_between_10_depth_plus_10_comb_out;
logic idx_between_6_min_depth_4_plus_6_reg_in;
logic idx_between_6_min_depth_4_plus_6_reg_write_en;
logic idx_between_6_min_depth_4_plus_6_reg_clk;
logic idx_between_6_min_depth_4_plus_6_reg_reset;
logic idx_between_6_min_depth_4_plus_6_reg_out;
logic idx_between_6_min_depth_4_plus_6_reg_done;
logic [31:0] index_lt_min_depth_4_plus_6_left;
logic [31:0] index_lt_min_depth_4_plus_6_right;
logic index_lt_min_depth_4_plus_6_out;
logic idx_between_6_min_depth_4_plus_6_comb_left;
logic idx_between_6_min_depth_4_plus_6_comb_right;
logic idx_between_6_min_depth_4_plus_6_comb_out;
logic idx_between_depth_plus_7_depth_plus_8_reg_in;
logic idx_between_depth_plus_7_depth_plus_8_reg_write_en;
logic idx_between_depth_plus_7_depth_plus_8_reg_clk;
logic idx_between_depth_plus_7_depth_plus_8_reg_reset;
logic idx_between_depth_plus_7_depth_plus_8_reg_out;
logic idx_between_depth_plus_7_depth_plus_8_reg_done;
logic [31:0] index_ge_depth_plus_7_left;
logic [31:0] index_ge_depth_plus_7_right;
logic index_ge_depth_plus_7_out;
logic idx_between_depth_plus_7_depth_plus_8_comb_left;
logic idx_between_depth_plus_7_depth_plus_8_comb_right;
logic idx_between_depth_plus_7_depth_plus_8_comb_out;
logic cond_in;
logic cond_write_en;
logic cond_clk;
logic cond_reset;
logic cond_out;
logic cond_done;
logic cond_wire_in;
logic cond_wire_out;
logic cond0_in;
logic cond0_write_en;
logic cond0_clk;
logic cond0_reset;
logic cond0_out;
logic cond0_done;
logic cond_wire0_in;
logic cond_wire0_out;
logic cond1_in;
logic cond1_write_en;
logic cond1_clk;
logic cond1_reset;
logic cond1_out;
logic cond1_done;
logic cond_wire1_in;
logic cond_wire1_out;
logic cond2_in;
logic cond2_write_en;
logic cond2_clk;
logic cond2_reset;
logic cond2_out;
logic cond2_done;
logic cond_wire2_in;
logic cond_wire2_out;
logic cond3_in;
logic cond3_write_en;
logic cond3_clk;
logic cond3_reset;
logic cond3_out;
logic cond3_done;
logic cond_wire3_in;
logic cond_wire3_out;
logic cond4_in;
logic cond4_write_en;
logic cond4_clk;
logic cond4_reset;
logic cond4_out;
logic cond4_done;
logic cond_wire4_in;
logic cond_wire4_out;
logic cond5_in;
logic cond5_write_en;
logic cond5_clk;
logic cond5_reset;
logic cond5_out;
logic cond5_done;
logic cond_wire5_in;
logic cond_wire5_out;
logic cond6_in;
logic cond6_write_en;
logic cond6_clk;
logic cond6_reset;
logic cond6_out;
logic cond6_done;
logic cond_wire6_in;
logic cond_wire6_out;
logic cond7_in;
logic cond7_write_en;
logic cond7_clk;
logic cond7_reset;
logic cond7_out;
logic cond7_done;
logic cond_wire7_in;
logic cond_wire7_out;
logic cond8_in;
logic cond8_write_en;
logic cond8_clk;
logic cond8_reset;
logic cond8_out;
logic cond8_done;
logic cond_wire8_in;
logic cond_wire8_out;
logic cond9_in;
logic cond9_write_en;
logic cond9_clk;
logic cond9_reset;
logic cond9_out;
logic cond9_done;
logic cond_wire9_in;
logic cond_wire9_out;
logic cond10_in;
logic cond10_write_en;
logic cond10_clk;
logic cond10_reset;
logic cond10_out;
logic cond10_done;
logic cond_wire10_in;
logic cond_wire10_out;
logic cond11_in;
logic cond11_write_en;
logic cond11_clk;
logic cond11_reset;
logic cond11_out;
logic cond11_done;
logic cond_wire11_in;
logic cond_wire11_out;
logic cond12_in;
logic cond12_write_en;
logic cond12_clk;
logic cond12_reset;
logic cond12_out;
logic cond12_done;
logic cond_wire12_in;
logic cond_wire12_out;
logic cond13_in;
logic cond13_write_en;
logic cond13_clk;
logic cond13_reset;
logic cond13_out;
logic cond13_done;
logic cond_wire13_in;
logic cond_wire13_out;
logic cond14_in;
logic cond14_write_en;
logic cond14_clk;
logic cond14_reset;
logic cond14_out;
logic cond14_done;
logic cond_wire14_in;
logic cond_wire14_out;
logic cond15_in;
logic cond15_write_en;
logic cond15_clk;
logic cond15_reset;
logic cond15_out;
logic cond15_done;
logic cond_wire15_in;
logic cond_wire15_out;
logic cond16_in;
logic cond16_write_en;
logic cond16_clk;
logic cond16_reset;
logic cond16_out;
logic cond16_done;
logic cond_wire16_in;
logic cond_wire16_out;
logic cond17_in;
logic cond17_write_en;
logic cond17_clk;
logic cond17_reset;
logic cond17_out;
logic cond17_done;
logic cond_wire17_in;
logic cond_wire17_out;
logic cond18_in;
logic cond18_write_en;
logic cond18_clk;
logic cond18_reset;
logic cond18_out;
logic cond18_done;
logic cond_wire18_in;
logic cond_wire18_out;
logic cond19_in;
logic cond19_write_en;
logic cond19_clk;
logic cond19_reset;
logic cond19_out;
logic cond19_done;
logic cond_wire19_in;
logic cond_wire19_out;
logic cond20_in;
logic cond20_write_en;
logic cond20_clk;
logic cond20_reset;
logic cond20_out;
logic cond20_done;
logic cond_wire20_in;
logic cond_wire20_out;
logic cond21_in;
logic cond21_write_en;
logic cond21_clk;
logic cond21_reset;
logic cond21_out;
logic cond21_done;
logic cond_wire21_in;
logic cond_wire21_out;
logic cond22_in;
logic cond22_write_en;
logic cond22_clk;
logic cond22_reset;
logic cond22_out;
logic cond22_done;
logic cond_wire22_in;
logic cond_wire22_out;
logic cond23_in;
logic cond23_write_en;
logic cond23_clk;
logic cond23_reset;
logic cond23_out;
logic cond23_done;
logic cond_wire23_in;
logic cond_wire23_out;
logic cond24_in;
logic cond24_write_en;
logic cond24_clk;
logic cond24_reset;
logic cond24_out;
logic cond24_done;
logic cond_wire24_in;
logic cond_wire24_out;
logic cond25_in;
logic cond25_write_en;
logic cond25_clk;
logic cond25_reset;
logic cond25_out;
logic cond25_done;
logic cond_wire25_in;
logic cond_wire25_out;
logic cond26_in;
logic cond26_write_en;
logic cond26_clk;
logic cond26_reset;
logic cond26_out;
logic cond26_done;
logic cond_wire26_in;
logic cond_wire26_out;
logic cond27_in;
logic cond27_write_en;
logic cond27_clk;
logic cond27_reset;
logic cond27_out;
logic cond27_done;
logic cond_wire27_in;
logic cond_wire27_out;
logic cond28_in;
logic cond28_write_en;
logic cond28_clk;
logic cond28_reset;
logic cond28_out;
logic cond28_done;
logic cond_wire28_in;
logic cond_wire28_out;
logic cond29_in;
logic cond29_write_en;
logic cond29_clk;
logic cond29_reset;
logic cond29_out;
logic cond29_done;
logic cond_wire29_in;
logic cond_wire29_out;
logic cond30_in;
logic cond30_write_en;
logic cond30_clk;
logic cond30_reset;
logic cond30_out;
logic cond30_done;
logic cond_wire30_in;
logic cond_wire30_out;
logic cond31_in;
logic cond31_write_en;
logic cond31_clk;
logic cond31_reset;
logic cond31_out;
logic cond31_done;
logic cond_wire31_in;
logic cond_wire31_out;
logic cond32_in;
logic cond32_write_en;
logic cond32_clk;
logic cond32_reset;
logic cond32_out;
logic cond32_done;
logic cond_wire32_in;
logic cond_wire32_out;
logic cond33_in;
logic cond33_write_en;
logic cond33_clk;
logic cond33_reset;
logic cond33_out;
logic cond33_done;
logic cond_wire33_in;
logic cond_wire33_out;
logic cond34_in;
logic cond34_write_en;
logic cond34_clk;
logic cond34_reset;
logic cond34_out;
logic cond34_done;
logic cond_wire34_in;
logic cond_wire34_out;
logic cond35_in;
logic cond35_write_en;
logic cond35_clk;
logic cond35_reset;
logic cond35_out;
logic cond35_done;
logic cond_wire35_in;
logic cond_wire35_out;
logic cond36_in;
logic cond36_write_en;
logic cond36_clk;
logic cond36_reset;
logic cond36_out;
logic cond36_done;
logic cond_wire36_in;
logic cond_wire36_out;
logic cond37_in;
logic cond37_write_en;
logic cond37_clk;
logic cond37_reset;
logic cond37_out;
logic cond37_done;
logic cond_wire37_in;
logic cond_wire37_out;
logic cond38_in;
logic cond38_write_en;
logic cond38_clk;
logic cond38_reset;
logic cond38_out;
logic cond38_done;
logic cond_wire38_in;
logic cond_wire38_out;
logic cond39_in;
logic cond39_write_en;
logic cond39_clk;
logic cond39_reset;
logic cond39_out;
logic cond39_done;
logic cond_wire39_in;
logic cond_wire39_out;
logic cond40_in;
logic cond40_write_en;
logic cond40_clk;
logic cond40_reset;
logic cond40_out;
logic cond40_done;
logic cond_wire40_in;
logic cond_wire40_out;
logic cond41_in;
logic cond41_write_en;
logic cond41_clk;
logic cond41_reset;
logic cond41_out;
logic cond41_done;
logic cond_wire41_in;
logic cond_wire41_out;
logic cond42_in;
logic cond42_write_en;
logic cond42_clk;
logic cond42_reset;
logic cond42_out;
logic cond42_done;
logic cond_wire42_in;
logic cond_wire42_out;
logic cond43_in;
logic cond43_write_en;
logic cond43_clk;
logic cond43_reset;
logic cond43_out;
logic cond43_done;
logic cond_wire43_in;
logic cond_wire43_out;
logic cond44_in;
logic cond44_write_en;
logic cond44_clk;
logic cond44_reset;
logic cond44_out;
logic cond44_done;
logic cond_wire44_in;
logic cond_wire44_out;
logic cond45_in;
logic cond45_write_en;
logic cond45_clk;
logic cond45_reset;
logic cond45_out;
logic cond45_done;
logic cond_wire45_in;
logic cond_wire45_out;
logic cond46_in;
logic cond46_write_en;
logic cond46_clk;
logic cond46_reset;
logic cond46_out;
logic cond46_done;
logic cond_wire46_in;
logic cond_wire46_out;
logic cond47_in;
logic cond47_write_en;
logic cond47_clk;
logic cond47_reset;
logic cond47_out;
logic cond47_done;
logic cond_wire47_in;
logic cond_wire47_out;
logic cond48_in;
logic cond48_write_en;
logic cond48_clk;
logic cond48_reset;
logic cond48_out;
logic cond48_done;
logic cond_wire48_in;
logic cond_wire48_out;
logic cond49_in;
logic cond49_write_en;
logic cond49_clk;
logic cond49_reset;
logic cond49_out;
logic cond49_done;
logic cond_wire49_in;
logic cond_wire49_out;
logic cond50_in;
logic cond50_write_en;
logic cond50_clk;
logic cond50_reset;
logic cond50_out;
logic cond50_done;
logic cond_wire50_in;
logic cond_wire50_out;
logic cond51_in;
logic cond51_write_en;
logic cond51_clk;
logic cond51_reset;
logic cond51_out;
logic cond51_done;
logic cond_wire51_in;
logic cond_wire51_out;
logic cond52_in;
logic cond52_write_en;
logic cond52_clk;
logic cond52_reset;
logic cond52_out;
logic cond52_done;
logic cond_wire52_in;
logic cond_wire52_out;
logic cond53_in;
logic cond53_write_en;
logic cond53_clk;
logic cond53_reset;
logic cond53_out;
logic cond53_done;
logic cond_wire53_in;
logic cond_wire53_out;
logic cond54_in;
logic cond54_write_en;
logic cond54_clk;
logic cond54_reset;
logic cond54_out;
logic cond54_done;
logic cond_wire54_in;
logic cond_wire54_out;
logic cond55_in;
logic cond55_write_en;
logic cond55_clk;
logic cond55_reset;
logic cond55_out;
logic cond55_done;
logic cond_wire55_in;
logic cond_wire55_out;
logic cond56_in;
logic cond56_write_en;
logic cond56_clk;
logic cond56_reset;
logic cond56_out;
logic cond56_done;
logic cond_wire56_in;
logic cond_wire56_out;
logic cond57_in;
logic cond57_write_en;
logic cond57_clk;
logic cond57_reset;
logic cond57_out;
logic cond57_done;
logic cond_wire57_in;
logic cond_wire57_out;
logic cond58_in;
logic cond58_write_en;
logic cond58_clk;
logic cond58_reset;
logic cond58_out;
logic cond58_done;
logic cond_wire58_in;
logic cond_wire58_out;
logic cond59_in;
logic cond59_write_en;
logic cond59_clk;
logic cond59_reset;
logic cond59_out;
logic cond59_done;
logic cond_wire59_in;
logic cond_wire59_out;
logic cond60_in;
logic cond60_write_en;
logic cond60_clk;
logic cond60_reset;
logic cond60_out;
logic cond60_done;
logic cond_wire60_in;
logic cond_wire60_out;
logic cond61_in;
logic cond61_write_en;
logic cond61_clk;
logic cond61_reset;
logic cond61_out;
logic cond61_done;
logic cond_wire61_in;
logic cond_wire61_out;
logic cond62_in;
logic cond62_write_en;
logic cond62_clk;
logic cond62_reset;
logic cond62_out;
logic cond62_done;
logic cond_wire62_in;
logic cond_wire62_out;
logic cond63_in;
logic cond63_write_en;
logic cond63_clk;
logic cond63_reset;
logic cond63_out;
logic cond63_done;
logic cond_wire63_in;
logic cond_wire63_out;
logic cond64_in;
logic cond64_write_en;
logic cond64_clk;
logic cond64_reset;
logic cond64_out;
logic cond64_done;
logic cond_wire64_in;
logic cond_wire64_out;
logic cond65_in;
logic cond65_write_en;
logic cond65_clk;
logic cond65_reset;
logic cond65_out;
logic cond65_done;
logic cond_wire65_in;
logic cond_wire65_out;
logic cond66_in;
logic cond66_write_en;
logic cond66_clk;
logic cond66_reset;
logic cond66_out;
logic cond66_done;
logic cond_wire66_in;
logic cond_wire66_out;
logic cond67_in;
logic cond67_write_en;
logic cond67_clk;
logic cond67_reset;
logic cond67_out;
logic cond67_done;
logic cond_wire67_in;
logic cond_wire67_out;
logic cond68_in;
logic cond68_write_en;
logic cond68_clk;
logic cond68_reset;
logic cond68_out;
logic cond68_done;
logic cond_wire68_in;
logic cond_wire68_out;
logic fsm_in;
logic fsm_write_en;
logic fsm_clk;
logic fsm_reset;
logic fsm_out;
logic fsm_done;
logic ud_out;
logic adder_left;
logic adder_right;
logic adder_out;
logic ud0_out;
logic adder0_left;
logic adder0_right;
logic adder0_out;
logic signal_reg_in;
logic signal_reg_write_en;
logic signal_reg_clk;
logic signal_reg_reset;
logic signal_reg_out;
logic signal_reg_done;
logic [1:0] fsm0_in;
logic fsm0_write_en;
logic fsm0_clk;
logic fsm0_reset;
logic [1:0] fsm0_out;
logic fsm0_done;
logic early_reset_static_par_go_in;
logic early_reset_static_par_go_out;
logic early_reset_static_par_done_in;
logic early_reset_static_par_done_out;
logic early_reset_static_par0_go_in;
logic early_reset_static_par0_go_out;
logic early_reset_static_par0_done_in;
logic early_reset_static_par0_done_out;
logic wrapper_early_reset_static_par_go_in;
logic wrapper_early_reset_static_par_go_out;
logic wrapper_early_reset_static_par_done_in;
logic wrapper_early_reset_static_par_done_out;
logic while_wrapper_early_reset_static_par0_go_in;
logic while_wrapper_early_reset_static_par0_go_out;
logic while_wrapper_early_reset_static_par0_done_in;
logic while_wrapper_early_reset_static_par0_done_out;
logic tdcc_go_in;
logic tdcc_go_out;
logic tdcc_done_in;
logic tdcc_done_out;
std_reg # (
    .WIDTH(32)
) min_depth_4 (
    .clk(min_depth_4_clk),
    .done(min_depth_4_done),
    .in(min_depth_4_in),
    .out(min_depth_4_out),
    .reset(min_depth_4_reset),
    .write_en(min_depth_4_write_en)
);
std_reg # (
    .WIDTH(32)
) iter_limit (
    .clk(iter_limit_clk),
    .done(iter_limit_done),
    .in(iter_limit_in),
    .out(iter_limit_out),
    .reset(iter_limit_reset),
    .write_en(iter_limit_write_en)
);
std_add # (
    .WIDTH(32)
) depth_plus_8 (
    .left(depth_plus_8_left),
    .out(depth_plus_8_out),
    .right(depth_plus_8_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_9 (
    .left(depth_plus_9_left),
    .out(depth_plus_9_out),
    .right(depth_plus_9_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_2 (
    .left(min_depth_4_plus_2_left),
    .out(min_depth_4_plus_2_out),
    .right(min_depth_4_plus_2_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_2 (
    .left(depth_plus_2_left),
    .out(depth_plus_2_out),
    .right(depth_plus_2_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_11 (
    .left(depth_plus_11_left),
    .out(depth_plus_11_out),
    .right(depth_plus_11_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_7 (
    .left(min_depth_4_plus_7_left),
    .out(min_depth_4_plus_7_out),
    .right(min_depth_4_plus_7_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_7 (
    .left(depth_plus_7_left),
    .out(depth_plus_7_out),
    .right(depth_plus_7_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_3 (
    .left(depth_plus_3_left),
    .out(depth_plus_3_out),
    .right(depth_plus_3_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_3 (
    .left(min_depth_4_plus_3_left),
    .out(min_depth_4_plus_3_out),
    .right(min_depth_4_plus_3_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_5 (
    .left(depth_plus_5_left),
    .out(depth_plus_5_out),
    .right(depth_plus_5_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_6 (
    .left(depth_plus_6_left),
    .out(depth_plus_6_out),
    .right(depth_plus_6_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_10 (
    .left(depth_plus_10_left),
    .out(depth_plus_10_out),
    .right(depth_plus_10_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_4 (
    .left(depth_plus_4_left),
    .out(depth_plus_4_out),
    .right(depth_plus_4_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_4 (
    .left(min_depth_4_plus_4_left),
    .out(min_depth_4_plus_4_out),
    .right(min_depth_4_plus_4_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_5 (
    .left(min_depth_4_plus_5_left),
    .out(min_depth_4_plus_5_out),
    .right(min_depth_4_plus_5_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_0 (
    .left(depth_plus_0_left),
    .out(depth_plus_0_out),
    .right(depth_plus_0_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_1 (
    .left(depth_plus_1_left),
    .out(depth_plus_1_out),
    .right(depth_plus_1_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_1 (
    .left(min_depth_4_plus_1_left),
    .out(min_depth_4_plus_1_out),
    .right(min_depth_4_plus_1_right)
);
std_add # (
    .WIDTH(32)
) depth_plus_12 (
    .left(depth_plus_12_left),
    .out(depth_plus_12_out),
    .right(depth_plus_12_right)
);
std_add # (
    .WIDTH(32)
) min_depth_4_plus_6 (
    .left(min_depth_4_plus_6_left),
    .out(min_depth_4_plus_6_out),
    .right(min_depth_4_plus_6_right)
);
mac_pe pe_0_0 (
    .clk(pe_0_0_clk),
    .done(pe_0_0_done),
    .go(pe_0_0_go),
    .left(pe_0_0_left),
    .mul_ready(pe_0_0_mul_ready),
    .out(pe_0_0_out),
    .reset(pe_0_0_reset),
    .top(pe_0_0_top)
);
std_reg # (
    .WIDTH(32)
) top_0_0 (
    .clk(top_0_0_clk),
    .done(top_0_0_done),
    .in(top_0_0_in),
    .out(top_0_0_out),
    .reset(top_0_0_reset),
    .write_en(top_0_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_0 (
    .clk(left_0_0_clk),
    .done(left_0_0_done),
    .in(left_0_0_in),
    .out(left_0_0_out),
    .reset(left_0_0_reset),
    .write_en(left_0_0_write_en)
);
mac_pe pe_0_1 (
    .clk(pe_0_1_clk),
    .done(pe_0_1_done),
    .go(pe_0_1_go),
    .left(pe_0_1_left),
    .mul_ready(pe_0_1_mul_ready),
    .out(pe_0_1_out),
    .reset(pe_0_1_reset),
    .top(pe_0_1_top)
);
std_reg # (
    .WIDTH(32)
) top_0_1 (
    .clk(top_0_1_clk),
    .done(top_0_1_done),
    .in(top_0_1_in),
    .out(top_0_1_out),
    .reset(top_0_1_reset),
    .write_en(top_0_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_1 (
    .clk(left_0_1_clk),
    .done(left_0_1_done),
    .in(left_0_1_in),
    .out(left_0_1_out),
    .reset(left_0_1_reset),
    .write_en(left_0_1_write_en)
);
mac_pe pe_0_2 (
    .clk(pe_0_2_clk),
    .done(pe_0_2_done),
    .go(pe_0_2_go),
    .left(pe_0_2_left),
    .mul_ready(pe_0_2_mul_ready),
    .out(pe_0_2_out),
    .reset(pe_0_2_reset),
    .top(pe_0_2_top)
);
std_reg # (
    .WIDTH(32)
) top_0_2 (
    .clk(top_0_2_clk),
    .done(top_0_2_done),
    .in(top_0_2_in),
    .out(top_0_2_out),
    .reset(top_0_2_reset),
    .write_en(top_0_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_2 (
    .clk(left_0_2_clk),
    .done(left_0_2_done),
    .in(left_0_2_in),
    .out(left_0_2_out),
    .reset(left_0_2_reset),
    .write_en(left_0_2_write_en)
);
mac_pe pe_0_3 (
    .clk(pe_0_3_clk),
    .done(pe_0_3_done),
    .go(pe_0_3_go),
    .left(pe_0_3_left),
    .mul_ready(pe_0_3_mul_ready),
    .out(pe_0_3_out),
    .reset(pe_0_3_reset),
    .top(pe_0_3_top)
);
std_reg # (
    .WIDTH(32)
) top_0_3 (
    .clk(top_0_3_clk),
    .done(top_0_3_done),
    .in(top_0_3_in),
    .out(top_0_3_out),
    .reset(top_0_3_reset),
    .write_en(top_0_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_3 (
    .clk(left_0_3_clk),
    .done(left_0_3_done),
    .in(left_0_3_in),
    .out(left_0_3_out),
    .reset(left_0_3_reset),
    .write_en(left_0_3_write_en)
);
mac_pe pe_1_0 (
    .clk(pe_1_0_clk),
    .done(pe_1_0_done),
    .go(pe_1_0_go),
    .left(pe_1_0_left),
    .mul_ready(pe_1_0_mul_ready),
    .out(pe_1_0_out),
    .reset(pe_1_0_reset),
    .top(pe_1_0_top)
);
std_reg # (
    .WIDTH(32)
) top_1_0 (
    .clk(top_1_0_clk),
    .done(top_1_0_done),
    .in(top_1_0_in),
    .out(top_1_0_out),
    .reset(top_1_0_reset),
    .write_en(top_1_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_0 (
    .clk(left_1_0_clk),
    .done(left_1_0_done),
    .in(left_1_0_in),
    .out(left_1_0_out),
    .reset(left_1_0_reset),
    .write_en(left_1_0_write_en)
);
mac_pe pe_1_1 (
    .clk(pe_1_1_clk),
    .done(pe_1_1_done),
    .go(pe_1_1_go),
    .left(pe_1_1_left),
    .mul_ready(pe_1_1_mul_ready),
    .out(pe_1_1_out),
    .reset(pe_1_1_reset),
    .top(pe_1_1_top)
);
std_reg # (
    .WIDTH(32)
) top_1_1 (
    .clk(top_1_1_clk),
    .done(top_1_1_done),
    .in(top_1_1_in),
    .out(top_1_1_out),
    .reset(top_1_1_reset),
    .write_en(top_1_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_1 (
    .clk(left_1_1_clk),
    .done(left_1_1_done),
    .in(left_1_1_in),
    .out(left_1_1_out),
    .reset(left_1_1_reset),
    .write_en(left_1_1_write_en)
);
mac_pe pe_1_2 (
    .clk(pe_1_2_clk),
    .done(pe_1_2_done),
    .go(pe_1_2_go),
    .left(pe_1_2_left),
    .mul_ready(pe_1_2_mul_ready),
    .out(pe_1_2_out),
    .reset(pe_1_2_reset),
    .top(pe_1_2_top)
);
std_reg # (
    .WIDTH(32)
) top_1_2 (
    .clk(top_1_2_clk),
    .done(top_1_2_done),
    .in(top_1_2_in),
    .out(top_1_2_out),
    .reset(top_1_2_reset),
    .write_en(top_1_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_2 (
    .clk(left_1_2_clk),
    .done(left_1_2_done),
    .in(left_1_2_in),
    .out(left_1_2_out),
    .reset(left_1_2_reset),
    .write_en(left_1_2_write_en)
);
mac_pe pe_1_3 (
    .clk(pe_1_3_clk),
    .done(pe_1_3_done),
    .go(pe_1_3_go),
    .left(pe_1_3_left),
    .mul_ready(pe_1_3_mul_ready),
    .out(pe_1_3_out),
    .reset(pe_1_3_reset),
    .top(pe_1_3_top)
);
std_reg # (
    .WIDTH(32)
) top_1_3 (
    .clk(top_1_3_clk),
    .done(top_1_3_done),
    .in(top_1_3_in),
    .out(top_1_3_out),
    .reset(top_1_3_reset),
    .write_en(top_1_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_3 (
    .clk(left_1_3_clk),
    .done(left_1_3_done),
    .in(left_1_3_in),
    .out(left_1_3_out),
    .reset(left_1_3_reset),
    .write_en(left_1_3_write_en)
);
mac_pe pe_2_0 (
    .clk(pe_2_0_clk),
    .done(pe_2_0_done),
    .go(pe_2_0_go),
    .left(pe_2_0_left),
    .mul_ready(pe_2_0_mul_ready),
    .out(pe_2_0_out),
    .reset(pe_2_0_reset),
    .top(pe_2_0_top)
);
std_reg # (
    .WIDTH(32)
) top_2_0 (
    .clk(top_2_0_clk),
    .done(top_2_0_done),
    .in(top_2_0_in),
    .out(top_2_0_out),
    .reset(top_2_0_reset),
    .write_en(top_2_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_0 (
    .clk(left_2_0_clk),
    .done(left_2_0_done),
    .in(left_2_0_in),
    .out(left_2_0_out),
    .reset(left_2_0_reset),
    .write_en(left_2_0_write_en)
);
mac_pe pe_2_1 (
    .clk(pe_2_1_clk),
    .done(pe_2_1_done),
    .go(pe_2_1_go),
    .left(pe_2_1_left),
    .mul_ready(pe_2_1_mul_ready),
    .out(pe_2_1_out),
    .reset(pe_2_1_reset),
    .top(pe_2_1_top)
);
std_reg # (
    .WIDTH(32)
) top_2_1 (
    .clk(top_2_1_clk),
    .done(top_2_1_done),
    .in(top_2_1_in),
    .out(top_2_1_out),
    .reset(top_2_1_reset),
    .write_en(top_2_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_1 (
    .clk(left_2_1_clk),
    .done(left_2_1_done),
    .in(left_2_1_in),
    .out(left_2_1_out),
    .reset(left_2_1_reset),
    .write_en(left_2_1_write_en)
);
mac_pe pe_2_2 (
    .clk(pe_2_2_clk),
    .done(pe_2_2_done),
    .go(pe_2_2_go),
    .left(pe_2_2_left),
    .mul_ready(pe_2_2_mul_ready),
    .out(pe_2_2_out),
    .reset(pe_2_2_reset),
    .top(pe_2_2_top)
);
std_reg # (
    .WIDTH(32)
) top_2_2 (
    .clk(top_2_2_clk),
    .done(top_2_2_done),
    .in(top_2_2_in),
    .out(top_2_2_out),
    .reset(top_2_2_reset),
    .write_en(top_2_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_2 (
    .clk(left_2_2_clk),
    .done(left_2_2_done),
    .in(left_2_2_in),
    .out(left_2_2_out),
    .reset(left_2_2_reset),
    .write_en(left_2_2_write_en)
);
mac_pe pe_2_3 (
    .clk(pe_2_3_clk),
    .done(pe_2_3_done),
    .go(pe_2_3_go),
    .left(pe_2_3_left),
    .mul_ready(pe_2_3_mul_ready),
    .out(pe_2_3_out),
    .reset(pe_2_3_reset),
    .top(pe_2_3_top)
);
std_reg # (
    .WIDTH(32)
) top_2_3 (
    .clk(top_2_3_clk),
    .done(top_2_3_done),
    .in(top_2_3_in),
    .out(top_2_3_out),
    .reset(top_2_3_reset),
    .write_en(top_2_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_3 (
    .clk(left_2_3_clk),
    .done(left_2_3_done),
    .in(left_2_3_in),
    .out(left_2_3_out),
    .reset(left_2_3_reset),
    .write_en(left_2_3_write_en)
);
mac_pe pe_3_0 (
    .clk(pe_3_0_clk),
    .done(pe_3_0_done),
    .go(pe_3_0_go),
    .left(pe_3_0_left),
    .mul_ready(pe_3_0_mul_ready),
    .out(pe_3_0_out),
    .reset(pe_3_0_reset),
    .top(pe_3_0_top)
);
std_reg # (
    .WIDTH(32)
) top_3_0 (
    .clk(top_3_0_clk),
    .done(top_3_0_done),
    .in(top_3_0_in),
    .out(top_3_0_out),
    .reset(top_3_0_reset),
    .write_en(top_3_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_0 (
    .clk(left_3_0_clk),
    .done(left_3_0_done),
    .in(left_3_0_in),
    .out(left_3_0_out),
    .reset(left_3_0_reset),
    .write_en(left_3_0_write_en)
);
mac_pe pe_3_1 (
    .clk(pe_3_1_clk),
    .done(pe_3_1_done),
    .go(pe_3_1_go),
    .left(pe_3_1_left),
    .mul_ready(pe_3_1_mul_ready),
    .out(pe_3_1_out),
    .reset(pe_3_1_reset),
    .top(pe_3_1_top)
);
std_reg # (
    .WIDTH(32)
) top_3_1 (
    .clk(top_3_1_clk),
    .done(top_3_1_done),
    .in(top_3_1_in),
    .out(top_3_1_out),
    .reset(top_3_1_reset),
    .write_en(top_3_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_1 (
    .clk(left_3_1_clk),
    .done(left_3_1_done),
    .in(left_3_1_in),
    .out(left_3_1_out),
    .reset(left_3_1_reset),
    .write_en(left_3_1_write_en)
);
mac_pe pe_3_2 (
    .clk(pe_3_2_clk),
    .done(pe_3_2_done),
    .go(pe_3_2_go),
    .left(pe_3_2_left),
    .mul_ready(pe_3_2_mul_ready),
    .out(pe_3_2_out),
    .reset(pe_3_2_reset),
    .top(pe_3_2_top)
);
std_reg # (
    .WIDTH(32)
) top_3_2 (
    .clk(top_3_2_clk),
    .done(top_3_2_done),
    .in(top_3_2_in),
    .out(top_3_2_out),
    .reset(top_3_2_reset),
    .write_en(top_3_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_2 (
    .clk(left_3_2_clk),
    .done(left_3_2_done),
    .in(left_3_2_in),
    .out(left_3_2_out),
    .reset(left_3_2_reset),
    .write_en(left_3_2_write_en)
);
mac_pe pe_3_3 (
    .clk(pe_3_3_clk),
    .done(pe_3_3_done),
    .go(pe_3_3_go),
    .left(pe_3_3_left),
    .mul_ready(pe_3_3_mul_ready),
    .out(pe_3_3_out),
    .reset(pe_3_3_reset),
    .top(pe_3_3_top)
);
std_reg # (
    .WIDTH(32)
) top_3_3 (
    .clk(top_3_3_clk),
    .done(top_3_3_done),
    .in(top_3_3_in),
    .out(top_3_3_out),
    .reset(top_3_3_reset),
    .write_en(top_3_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_3 (
    .clk(left_3_3_clk),
    .done(left_3_3_done),
    .in(left_3_3_in),
    .out(left_3_3_out),
    .reset(left_3_3_reset),
    .write_en(left_3_3_write_en)
);
std_reg # (
    .WIDTH(3)
) t0_idx (
    .clk(t0_idx_clk),
    .done(t0_idx_done),
    .in(t0_idx_in),
    .out(t0_idx_out),
    .reset(t0_idx_reset),
    .write_en(t0_idx_write_en)
);
std_add # (
    .WIDTH(3)
) t0_add (
    .left(t0_add_left),
    .out(t0_add_out),
    .right(t0_add_right)
);
std_reg # (
    .WIDTH(3)
) t1_idx (
    .clk(t1_idx_clk),
    .done(t1_idx_done),
    .in(t1_idx_in),
    .out(t1_idx_out),
    .reset(t1_idx_reset),
    .write_en(t1_idx_write_en)
);
std_add # (
    .WIDTH(3)
) t1_add (
    .left(t1_add_left),
    .out(t1_add_out),
    .right(t1_add_right)
);
std_reg # (
    .WIDTH(3)
) t2_idx (
    .clk(t2_idx_clk),
    .done(t2_idx_done),
    .in(t2_idx_in),
    .out(t2_idx_out),
    .reset(t2_idx_reset),
    .write_en(t2_idx_write_en)
);
std_add # (
    .WIDTH(3)
) t2_add (
    .left(t2_add_left),
    .out(t2_add_out),
    .right(t2_add_right)
);
std_reg # (
    .WIDTH(3)
) t3_idx (
    .clk(t3_idx_clk),
    .done(t3_idx_done),
    .in(t3_idx_in),
    .out(t3_idx_out),
    .reset(t3_idx_reset),
    .write_en(t3_idx_write_en)
);
std_add # (
    .WIDTH(3)
) t3_add (
    .left(t3_add_left),
    .out(t3_add_out),
    .right(t3_add_right)
);
std_reg # (
    .WIDTH(3)
) l0_idx (
    .clk(l0_idx_clk),
    .done(l0_idx_done),
    .in(l0_idx_in),
    .out(l0_idx_out),
    .reset(l0_idx_reset),
    .write_en(l0_idx_write_en)
);
std_add # (
    .WIDTH(3)
) l0_add (
    .left(l0_add_left),
    .out(l0_add_out),
    .right(l0_add_right)
);
std_reg # (
    .WIDTH(3)
) l1_idx (
    .clk(l1_idx_clk),
    .done(l1_idx_done),
    .in(l1_idx_in),
    .out(l1_idx_out),
    .reset(l1_idx_reset),
    .write_en(l1_idx_write_en)
);
std_add # (
    .WIDTH(3)
) l1_add (
    .left(l1_add_left),
    .out(l1_add_out),
    .right(l1_add_right)
);
std_reg # (
    .WIDTH(3)
) l2_idx (
    .clk(l2_idx_clk),
    .done(l2_idx_done),
    .in(l2_idx_in),
    .out(l2_idx_out),
    .reset(l2_idx_reset),
    .write_en(l2_idx_write_en)
);
std_add # (
    .WIDTH(3)
) l2_add (
    .left(l2_add_left),
    .out(l2_add_out),
    .right(l2_add_right)
);
std_reg # (
    .WIDTH(3)
) l3_idx (
    .clk(l3_idx_clk),
    .done(l3_idx_done),
    .in(l3_idx_in),
    .out(l3_idx_out),
    .reset(l3_idx_reset),
    .write_en(l3_idx_write_en)
);
std_add # (
    .WIDTH(3)
) l3_add (
    .left(l3_add_left),
    .out(l3_add_out),
    .right(l3_add_right)
);
std_reg # (
    .WIDTH(32)
) idx (
    .clk(idx_clk),
    .done(idx_done),
    .in(idx_in),
    .out(idx_out),
    .reset(idx_reset),
    .write_en(idx_write_en)
);
std_add # (
    .WIDTH(32)
) idx_add (
    .left(idx_add_left),
    .out(idx_add_out),
    .right(idx_add_right)
);
std_lt # (
    .WIDTH(32)
) lt_iter_limit (
    .left(lt_iter_limit_left),
    .out(lt_iter_limit_out),
    .right(lt_iter_limit_right)
);
std_reg # (
    .WIDTH(1)
) cond_reg (
    .clk(cond_reg_clk),
    .done(cond_reg_done),
    .in(cond_reg_in),
    .out(cond_reg_out),
    .reset(cond_reg_reset),
    .write_en(cond_reg_write_en)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_8_depth_plus_9_reg (
    .clk(idx_between_depth_plus_8_depth_plus_9_reg_clk),
    .done(idx_between_depth_plus_8_depth_plus_9_reg_done),
    .in(idx_between_depth_plus_8_depth_plus_9_reg_in),
    .out(idx_between_depth_plus_8_depth_plus_9_reg_out),
    .reset(idx_between_depth_plus_8_depth_plus_9_reg_reset),
    .write_en(idx_between_depth_plus_8_depth_plus_9_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_9 (
    .left(index_lt_depth_plus_9_left),
    .out(index_lt_depth_plus_9_out),
    .right(index_lt_depth_plus_9_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_8 (
    .left(index_ge_depth_plus_8_left),
    .out(index_ge_depth_plus_8_out),
    .right(index_ge_depth_plus_8_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_8_depth_plus_9_comb (
    .left(idx_between_depth_plus_8_depth_plus_9_comb_left),
    .out(idx_between_depth_plus_8_depth_plus_9_comb_out),
    .right(idx_between_depth_plus_8_depth_plus_9_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_2_min_depth_4_plus_2_reg (
    .clk(idx_between_2_min_depth_4_plus_2_reg_clk),
    .done(idx_between_2_min_depth_4_plus_2_reg_done),
    .in(idx_between_2_min_depth_4_plus_2_reg_in),
    .out(idx_between_2_min_depth_4_plus_2_reg_out),
    .reset(idx_between_2_min_depth_4_plus_2_reg_reset),
    .write_en(idx_between_2_min_depth_4_plus_2_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_2 (
    .left(index_lt_min_depth_4_plus_2_left),
    .out(index_lt_min_depth_4_plus_2_out),
    .right(index_lt_min_depth_4_plus_2_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_2 (
    .left(index_ge_2_left),
    .out(index_ge_2_out),
    .right(index_ge_2_right)
);
std_and # (
    .WIDTH(1)
) idx_between_2_min_depth_4_plus_2_comb (
    .left(idx_between_2_min_depth_4_plus_2_comb_left),
    .out(idx_between_2_min_depth_4_plus_2_comb_out),
    .right(idx_between_2_min_depth_4_plus_2_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_2_depth_plus_2_reg (
    .clk(idx_between_2_depth_plus_2_reg_clk),
    .done(idx_between_2_depth_plus_2_reg_done),
    .in(idx_between_2_depth_plus_2_reg_in),
    .out(idx_between_2_depth_plus_2_reg_out),
    .reset(idx_between_2_depth_plus_2_reg_reset),
    .write_en(idx_between_2_depth_plus_2_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_2 (
    .left(index_lt_depth_plus_2_left),
    .out(index_lt_depth_plus_2_out),
    .right(index_lt_depth_plus_2_right)
);
std_and # (
    .WIDTH(1)
) idx_between_2_depth_plus_2_comb (
    .left(idx_between_2_depth_plus_2_comb_left),
    .out(idx_between_2_depth_plus_2_comb_out),
    .right(idx_between_2_depth_plus_2_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_11_depth_plus_11_reg (
    .clk(idx_between_11_depth_plus_11_reg_clk),
    .done(idx_between_11_depth_plus_11_reg_done),
    .in(idx_between_11_depth_plus_11_reg_in),
    .out(idx_between_11_depth_plus_11_reg_out),
    .reset(idx_between_11_depth_plus_11_reg_reset),
    .write_en(idx_between_11_depth_plus_11_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_11 (
    .left(index_lt_depth_plus_11_left),
    .out(index_lt_depth_plus_11_out),
    .right(index_lt_depth_plus_11_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_11 (
    .left(index_ge_11_left),
    .out(index_ge_11_out),
    .right(index_ge_11_right)
);
std_and # (
    .WIDTH(1)
) idx_between_11_depth_plus_11_comb (
    .left(idx_between_11_depth_plus_11_comb_left),
    .out(idx_between_11_depth_plus_11_comb_out),
    .right(idx_between_11_depth_plus_11_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_7_min_depth_4_plus_7_reg (
    .clk(idx_between_7_min_depth_4_plus_7_reg_clk),
    .done(idx_between_7_min_depth_4_plus_7_reg_done),
    .in(idx_between_7_min_depth_4_plus_7_reg_in),
    .out(idx_between_7_min_depth_4_plus_7_reg_out),
    .reset(idx_between_7_min_depth_4_plus_7_reg_reset),
    .write_en(idx_between_7_min_depth_4_plus_7_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_7 (
    .left(index_lt_min_depth_4_plus_7_left),
    .out(index_lt_min_depth_4_plus_7_out),
    .right(index_lt_min_depth_4_plus_7_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_7 (
    .left(index_ge_7_left),
    .out(index_ge_7_out),
    .right(index_ge_7_right)
);
std_and # (
    .WIDTH(1)
) idx_between_7_min_depth_4_plus_7_comb (
    .left(idx_between_7_min_depth_4_plus_7_comb_left),
    .out(idx_between_7_min_depth_4_plus_7_comb_out),
    .right(idx_between_7_min_depth_4_plus_7_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_7_depth_plus_7_reg (
    .clk(idx_between_7_depth_plus_7_reg_clk),
    .done(idx_between_7_depth_plus_7_reg_done),
    .in(idx_between_7_depth_plus_7_reg_in),
    .out(idx_between_7_depth_plus_7_reg_out),
    .reset(idx_between_7_depth_plus_7_reg_reset),
    .write_en(idx_between_7_depth_plus_7_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_7 (
    .left(index_lt_depth_plus_7_left),
    .out(index_lt_depth_plus_7_out),
    .right(index_lt_depth_plus_7_right)
);
std_and # (
    .WIDTH(1)
) idx_between_7_depth_plus_7_comb (
    .left(idx_between_7_depth_plus_7_comb_left),
    .out(idx_between_7_depth_plus_7_comb_out),
    .right(idx_between_7_depth_plus_7_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_3_depth_plus_3_reg (
    .clk(idx_between_3_depth_plus_3_reg_clk),
    .done(idx_between_3_depth_plus_3_reg_done),
    .in(idx_between_3_depth_plus_3_reg_in),
    .out(idx_between_3_depth_plus_3_reg_out),
    .reset(idx_between_3_depth_plus_3_reg_reset),
    .write_en(idx_between_3_depth_plus_3_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_3 (
    .left(index_lt_depth_plus_3_left),
    .out(index_lt_depth_plus_3_out),
    .right(index_lt_depth_plus_3_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_3 (
    .left(index_ge_3_left),
    .out(index_ge_3_out),
    .right(index_ge_3_right)
);
std_and # (
    .WIDTH(1)
) idx_between_3_depth_plus_3_comb (
    .left(idx_between_3_depth_plus_3_comb_left),
    .out(idx_between_3_depth_plus_3_comb_out),
    .right(idx_between_3_depth_plus_3_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_3_min_depth_4_plus_3_reg (
    .clk(idx_between_3_min_depth_4_plus_3_reg_clk),
    .done(idx_between_3_min_depth_4_plus_3_reg_done),
    .in(idx_between_3_min_depth_4_plus_3_reg_in),
    .out(idx_between_3_min_depth_4_plus_3_reg_out),
    .reset(idx_between_3_min_depth_4_plus_3_reg_reset),
    .write_en(idx_between_3_min_depth_4_plus_3_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_3 (
    .left(index_lt_min_depth_4_plus_3_left),
    .out(index_lt_min_depth_4_plus_3_out),
    .right(index_lt_min_depth_4_plus_3_right)
);
std_and # (
    .WIDTH(1)
) idx_between_3_min_depth_4_plus_3_comb (
    .left(idx_between_3_min_depth_4_plus_3_comb_left),
    .out(idx_between_3_min_depth_4_plus_3_comb_out),
    .right(idx_between_3_min_depth_4_plus_3_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_5_depth_plus_6_reg (
    .clk(idx_between_depth_plus_5_depth_plus_6_reg_clk),
    .done(idx_between_depth_plus_5_depth_plus_6_reg_done),
    .in(idx_between_depth_plus_5_depth_plus_6_reg_in),
    .out(idx_between_depth_plus_5_depth_plus_6_reg_out),
    .reset(idx_between_depth_plus_5_depth_plus_6_reg_reset),
    .write_en(idx_between_depth_plus_5_depth_plus_6_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_6 (
    .left(index_lt_depth_plus_6_left),
    .out(index_lt_depth_plus_6_out),
    .right(index_lt_depth_plus_6_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_5 (
    .left(index_ge_depth_plus_5_left),
    .out(index_ge_depth_plus_5_out),
    .right(index_ge_depth_plus_5_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_5_depth_plus_6_comb (
    .left(idx_between_depth_plus_5_depth_plus_6_comb_left),
    .out(idx_between_depth_plus_5_depth_plus_6_comb_out),
    .right(idx_between_depth_plus_5_depth_plus_6_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_9_depth_plus_10_reg (
    .clk(idx_between_depth_plus_9_depth_plus_10_reg_clk),
    .done(idx_between_depth_plus_9_depth_plus_10_reg_done),
    .in(idx_between_depth_plus_9_depth_plus_10_reg_in),
    .out(idx_between_depth_plus_9_depth_plus_10_reg_out),
    .reset(idx_between_depth_plus_9_depth_plus_10_reg_reset),
    .write_en(idx_between_depth_plus_9_depth_plus_10_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_10 (
    .left(index_lt_depth_plus_10_left),
    .out(index_lt_depth_plus_10_out),
    .right(index_lt_depth_plus_10_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_9 (
    .left(index_ge_depth_plus_9_left),
    .out(index_ge_depth_plus_9_out),
    .right(index_ge_depth_plus_9_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_9_depth_plus_10_comb (
    .left(idx_between_depth_plus_9_depth_plus_10_comb_left),
    .out(idx_between_depth_plus_9_depth_plus_10_comb_out),
    .right(idx_between_depth_plus_9_depth_plus_10_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_8_depth_plus_8_reg (
    .clk(idx_between_8_depth_plus_8_reg_clk),
    .done(idx_between_8_depth_plus_8_reg_done),
    .in(idx_between_8_depth_plus_8_reg_in),
    .out(idx_between_8_depth_plus_8_reg_out),
    .reset(idx_between_8_depth_plus_8_reg_reset),
    .write_en(idx_between_8_depth_plus_8_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_8 (
    .left(index_lt_depth_plus_8_left),
    .out(index_lt_depth_plus_8_out),
    .right(index_lt_depth_plus_8_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_8 (
    .left(index_ge_8_left),
    .out(index_ge_8_out),
    .right(index_ge_8_right)
);
std_and # (
    .WIDTH(1)
) idx_between_8_depth_plus_8_comb (
    .left(idx_between_8_depth_plus_8_comb_left),
    .out(idx_between_8_depth_plus_8_comb_out),
    .right(idx_between_8_depth_plus_8_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_10_depth_plus_11_reg (
    .clk(idx_between_depth_plus_10_depth_plus_11_reg_clk),
    .done(idx_between_depth_plus_10_depth_plus_11_reg_done),
    .in(idx_between_depth_plus_10_depth_plus_11_reg_in),
    .out(idx_between_depth_plus_10_depth_plus_11_reg_out),
    .reset(idx_between_depth_plus_10_depth_plus_11_reg_reset),
    .write_en(idx_between_depth_plus_10_depth_plus_11_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_10 (
    .left(index_ge_depth_plus_10_left),
    .out(index_ge_depth_plus_10_out),
    .right(index_ge_depth_plus_10_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_10_depth_plus_11_comb (
    .left(idx_between_depth_plus_10_depth_plus_11_comb_left),
    .out(idx_between_depth_plus_10_depth_plus_11_comb_out),
    .right(idx_between_depth_plus_10_depth_plus_11_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_6_depth_plus_6_reg (
    .clk(idx_between_6_depth_plus_6_reg_clk),
    .done(idx_between_6_depth_plus_6_reg_done),
    .in(idx_between_6_depth_plus_6_reg_in),
    .out(idx_between_6_depth_plus_6_reg_out),
    .reset(idx_between_6_depth_plus_6_reg_reset),
    .write_en(idx_between_6_depth_plus_6_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_6 (
    .left(index_ge_6_left),
    .out(index_ge_6_out),
    .right(index_ge_6_right)
);
std_and # (
    .WIDTH(1)
) idx_between_6_depth_plus_6_comb (
    .left(idx_between_6_depth_plus_6_comb_left),
    .out(idx_between_6_depth_plus_6_comb_out),
    .right(idx_between_6_depth_plus_6_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_6_depth_plus_7_reg (
    .clk(idx_between_depth_plus_6_depth_plus_7_reg_clk),
    .done(idx_between_depth_plus_6_depth_plus_7_reg_done),
    .in(idx_between_depth_plus_6_depth_plus_7_reg_in),
    .out(idx_between_depth_plus_6_depth_plus_7_reg_out),
    .reset(idx_between_depth_plus_6_depth_plus_7_reg_reset),
    .write_en(idx_between_depth_plus_6_depth_plus_7_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_6 (
    .left(index_ge_depth_plus_6_left),
    .out(index_ge_depth_plus_6_out),
    .right(index_ge_depth_plus_6_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_6_depth_plus_7_comb (
    .left(idx_between_depth_plus_6_depth_plus_7_comb_left),
    .out(idx_between_depth_plus_6_depth_plus_7_comb_out),
    .right(idx_between_depth_plus_6_depth_plus_7_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_4_depth_plus_4_reg (
    .clk(idx_between_4_depth_plus_4_reg_clk),
    .done(idx_between_4_depth_plus_4_reg_done),
    .in(idx_between_4_depth_plus_4_reg_in),
    .out(idx_between_4_depth_plus_4_reg_out),
    .reset(idx_between_4_depth_plus_4_reg_reset),
    .write_en(idx_between_4_depth_plus_4_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_4 (
    .left(index_lt_depth_plus_4_left),
    .out(index_lt_depth_plus_4_out),
    .right(index_lt_depth_plus_4_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_4 (
    .left(index_ge_4_left),
    .out(index_ge_4_out),
    .right(index_ge_4_right)
);
std_and # (
    .WIDTH(1)
) idx_between_4_depth_plus_4_comb (
    .left(idx_between_4_depth_plus_4_comb_left),
    .out(idx_between_4_depth_plus_4_comb_out),
    .right(idx_between_4_depth_plus_4_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_4_min_depth_4_plus_4_reg (
    .clk(idx_between_4_min_depth_4_plus_4_reg_clk),
    .done(idx_between_4_min_depth_4_plus_4_reg_done),
    .in(idx_between_4_min_depth_4_plus_4_reg_in),
    .out(idx_between_4_min_depth_4_plus_4_reg_out),
    .reset(idx_between_4_min_depth_4_plus_4_reg_reset),
    .write_en(idx_between_4_min_depth_4_plus_4_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_4 (
    .left(index_lt_min_depth_4_plus_4_left),
    .out(index_lt_min_depth_4_plus_4_out),
    .right(index_lt_min_depth_4_plus_4_right)
);
std_and # (
    .WIDTH(1)
) idx_between_4_min_depth_4_plus_4_comb (
    .left(idx_between_4_min_depth_4_plus_4_comb_left),
    .out(idx_between_4_min_depth_4_plus_4_comb_out),
    .right(idx_between_4_min_depth_4_plus_4_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_5_depth_plus_5_reg (
    .clk(idx_between_5_depth_plus_5_reg_clk),
    .done(idx_between_5_depth_plus_5_reg_done),
    .in(idx_between_5_depth_plus_5_reg_in),
    .out(idx_between_5_depth_plus_5_reg_out),
    .reset(idx_between_5_depth_plus_5_reg_reset),
    .write_en(idx_between_5_depth_plus_5_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_5 (
    .left(index_lt_depth_plus_5_left),
    .out(index_lt_depth_plus_5_out),
    .right(index_lt_depth_plus_5_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_5 (
    .left(index_ge_5_left),
    .out(index_ge_5_out),
    .right(index_ge_5_right)
);
std_and # (
    .WIDTH(1)
) idx_between_5_depth_plus_5_comb (
    .left(idx_between_5_depth_plus_5_comb_left),
    .out(idx_between_5_depth_plus_5_comb_out),
    .right(idx_between_5_depth_plus_5_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_5_min_depth_4_plus_5_reg (
    .clk(idx_between_5_min_depth_4_plus_5_reg_clk),
    .done(idx_between_5_min_depth_4_plus_5_reg_done),
    .in(idx_between_5_min_depth_4_plus_5_reg_in),
    .out(idx_between_5_min_depth_4_plus_5_reg_out),
    .reset(idx_between_5_min_depth_4_plus_5_reg_reset),
    .write_en(idx_between_5_min_depth_4_plus_5_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_5 (
    .left(index_lt_min_depth_4_plus_5_left),
    .out(index_lt_min_depth_4_plus_5_out),
    .right(index_lt_min_depth_4_plus_5_right)
);
std_and # (
    .WIDTH(1)
) idx_between_5_min_depth_4_plus_5_comb (
    .left(idx_between_5_min_depth_4_plus_5_comb_left),
    .out(idx_between_5_min_depth_4_plus_5_comb_out),
    .right(idx_between_5_min_depth_4_plus_5_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_0_depth_plus_0_reg (
    .clk(idx_between_0_depth_plus_0_reg_clk),
    .done(idx_between_0_depth_plus_0_reg_done),
    .in(idx_between_0_depth_plus_0_reg_in),
    .out(idx_between_0_depth_plus_0_reg_out),
    .reset(idx_between_0_depth_plus_0_reg_reset),
    .write_en(idx_between_0_depth_plus_0_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_0 (
    .left(index_lt_depth_plus_0_left),
    .out(index_lt_depth_plus_0_out),
    .right(index_lt_depth_plus_0_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_9_depth_plus_9_reg (
    .clk(idx_between_9_depth_plus_9_reg_clk),
    .done(idx_between_9_depth_plus_9_reg_done),
    .in(idx_between_9_depth_plus_9_reg_in),
    .out(idx_between_9_depth_plus_9_reg_out),
    .reset(idx_between_9_depth_plus_9_reg_reset),
    .write_en(idx_between_9_depth_plus_9_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_9 (
    .left(index_ge_9_left),
    .out(index_ge_9_out),
    .right(index_ge_9_right)
);
std_and # (
    .WIDTH(1)
) idx_between_9_depth_plus_9_comb (
    .left(idx_between_9_depth_plus_9_comb_left),
    .out(idx_between_9_depth_plus_9_comb_out),
    .right(idx_between_9_depth_plus_9_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_1_depth_plus_1_reg (
    .clk(idx_between_1_depth_plus_1_reg_clk),
    .done(idx_between_1_depth_plus_1_reg_done),
    .in(idx_between_1_depth_plus_1_reg_in),
    .out(idx_between_1_depth_plus_1_reg_out),
    .reset(idx_between_1_depth_plus_1_reg_reset),
    .write_en(idx_between_1_depth_plus_1_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_1 (
    .left(index_lt_depth_plus_1_left),
    .out(index_lt_depth_plus_1_out),
    .right(index_lt_depth_plus_1_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_1 (
    .left(index_ge_1_left),
    .out(index_ge_1_out),
    .right(index_ge_1_right)
);
std_and # (
    .WIDTH(1)
) idx_between_1_depth_plus_1_comb (
    .left(idx_between_1_depth_plus_1_comb_left),
    .out(idx_between_1_depth_plus_1_comb_out),
    .right(idx_between_1_depth_plus_1_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_1_min_depth_4_plus_1_reg (
    .clk(idx_between_1_min_depth_4_plus_1_reg_clk),
    .done(idx_between_1_min_depth_4_plus_1_reg_done),
    .in(idx_between_1_min_depth_4_plus_1_reg_in),
    .out(idx_between_1_min_depth_4_plus_1_reg_out),
    .reset(idx_between_1_min_depth_4_plus_1_reg_reset),
    .write_en(idx_between_1_min_depth_4_plus_1_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_1 (
    .left(index_lt_min_depth_4_plus_1_left),
    .out(index_lt_min_depth_4_plus_1_out),
    .right(index_lt_min_depth_4_plus_1_right)
);
std_and # (
    .WIDTH(1)
) idx_between_1_min_depth_4_plus_1_comb (
    .left(idx_between_1_min_depth_4_plus_1_comb_left),
    .out(idx_between_1_min_depth_4_plus_1_comb_out),
    .right(idx_between_1_min_depth_4_plus_1_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_11_depth_plus_12_reg (
    .clk(idx_between_depth_plus_11_depth_plus_12_reg_clk),
    .done(idx_between_depth_plus_11_depth_plus_12_reg_done),
    .in(idx_between_depth_plus_11_depth_plus_12_reg_in),
    .out(idx_between_depth_plus_11_depth_plus_12_reg_out),
    .reset(idx_between_depth_plus_11_depth_plus_12_reg_reset),
    .write_en(idx_between_depth_plus_11_depth_plus_12_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_depth_plus_12 (
    .left(index_lt_depth_plus_12_left),
    .out(index_lt_depth_plus_12_out),
    .right(index_lt_depth_plus_12_right)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_11 (
    .left(index_ge_depth_plus_11_left),
    .out(index_ge_depth_plus_11_out),
    .right(index_ge_depth_plus_11_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_11_depth_plus_12_comb (
    .left(idx_between_depth_plus_11_depth_plus_12_comb_left),
    .out(idx_between_depth_plus_11_depth_plus_12_comb_out),
    .right(idx_between_depth_plus_11_depth_plus_12_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_10_depth_plus_10_reg (
    .clk(idx_between_10_depth_plus_10_reg_clk),
    .done(idx_between_10_depth_plus_10_reg_done),
    .in(idx_between_10_depth_plus_10_reg_in),
    .out(idx_between_10_depth_plus_10_reg_out),
    .reset(idx_between_10_depth_plus_10_reg_reset),
    .write_en(idx_between_10_depth_plus_10_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_10 (
    .left(index_ge_10_left),
    .out(index_ge_10_out),
    .right(index_ge_10_right)
);
std_and # (
    .WIDTH(1)
) idx_between_10_depth_plus_10_comb (
    .left(idx_between_10_depth_plus_10_comb_left),
    .out(idx_between_10_depth_plus_10_comb_out),
    .right(idx_between_10_depth_plus_10_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_6_min_depth_4_plus_6_reg (
    .clk(idx_between_6_min_depth_4_plus_6_reg_clk),
    .done(idx_between_6_min_depth_4_plus_6_reg_done),
    .in(idx_between_6_min_depth_4_plus_6_reg_in),
    .out(idx_between_6_min_depth_4_plus_6_reg_out),
    .reset(idx_between_6_min_depth_4_plus_6_reg_reset),
    .write_en(idx_between_6_min_depth_4_plus_6_reg_write_en)
);
std_lt # (
    .WIDTH(32)
) index_lt_min_depth_4_plus_6 (
    .left(index_lt_min_depth_4_plus_6_left),
    .out(index_lt_min_depth_4_plus_6_out),
    .right(index_lt_min_depth_4_plus_6_right)
);
std_and # (
    .WIDTH(1)
) idx_between_6_min_depth_4_plus_6_comb (
    .left(idx_between_6_min_depth_4_plus_6_comb_left),
    .out(idx_between_6_min_depth_4_plus_6_comb_out),
    .right(idx_between_6_min_depth_4_plus_6_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_depth_plus_7_depth_plus_8_reg (
    .clk(idx_between_depth_plus_7_depth_plus_8_reg_clk),
    .done(idx_between_depth_plus_7_depth_plus_8_reg_done),
    .in(idx_between_depth_plus_7_depth_plus_8_reg_in),
    .out(idx_between_depth_plus_7_depth_plus_8_reg_out),
    .reset(idx_between_depth_plus_7_depth_plus_8_reg_reset),
    .write_en(idx_between_depth_plus_7_depth_plus_8_reg_write_en)
);
std_ge # (
    .WIDTH(32)
) index_ge_depth_plus_7 (
    .left(index_ge_depth_plus_7_left),
    .out(index_ge_depth_plus_7_out),
    .right(index_ge_depth_plus_7_right)
);
std_and # (
    .WIDTH(1)
) idx_between_depth_plus_7_depth_plus_8_comb (
    .left(idx_between_depth_plus_7_depth_plus_8_comb_left),
    .out(idx_between_depth_plus_7_depth_plus_8_comb_out),
    .right(idx_between_depth_plus_7_depth_plus_8_comb_right)
);
std_reg # (
    .WIDTH(1)
) cond (
    .clk(cond_clk),
    .done(cond_done),
    .in(cond_in),
    .out(cond_out),
    .reset(cond_reset),
    .write_en(cond_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire (
    .in(cond_wire_in),
    .out(cond_wire_out)
);
std_reg # (
    .WIDTH(1)
) cond0 (
    .clk(cond0_clk),
    .done(cond0_done),
    .in(cond0_in),
    .out(cond0_out),
    .reset(cond0_reset),
    .write_en(cond0_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire0 (
    .in(cond_wire0_in),
    .out(cond_wire0_out)
);
std_reg # (
    .WIDTH(1)
) cond1 (
    .clk(cond1_clk),
    .done(cond1_done),
    .in(cond1_in),
    .out(cond1_out),
    .reset(cond1_reset),
    .write_en(cond1_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1 (
    .in(cond_wire1_in),
    .out(cond_wire1_out)
);
std_reg # (
    .WIDTH(1)
) cond2 (
    .clk(cond2_clk),
    .done(cond2_done),
    .in(cond2_in),
    .out(cond2_out),
    .reset(cond2_reset),
    .write_en(cond2_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire2 (
    .in(cond_wire2_in),
    .out(cond_wire2_out)
);
std_reg # (
    .WIDTH(1)
) cond3 (
    .clk(cond3_clk),
    .done(cond3_done),
    .in(cond3_in),
    .out(cond3_out),
    .reset(cond3_reset),
    .write_en(cond3_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire3 (
    .in(cond_wire3_in),
    .out(cond_wire3_out)
);
std_reg # (
    .WIDTH(1)
) cond4 (
    .clk(cond4_clk),
    .done(cond4_done),
    .in(cond4_in),
    .out(cond4_out),
    .reset(cond4_reset),
    .write_en(cond4_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire4 (
    .in(cond_wire4_in),
    .out(cond_wire4_out)
);
std_reg # (
    .WIDTH(1)
) cond5 (
    .clk(cond5_clk),
    .done(cond5_done),
    .in(cond5_in),
    .out(cond5_out),
    .reset(cond5_reset),
    .write_en(cond5_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire5 (
    .in(cond_wire5_in),
    .out(cond_wire5_out)
);
std_reg # (
    .WIDTH(1)
) cond6 (
    .clk(cond6_clk),
    .done(cond6_done),
    .in(cond6_in),
    .out(cond6_out),
    .reset(cond6_reset),
    .write_en(cond6_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire6 (
    .in(cond_wire6_in),
    .out(cond_wire6_out)
);
std_reg # (
    .WIDTH(1)
) cond7 (
    .clk(cond7_clk),
    .done(cond7_done),
    .in(cond7_in),
    .out(cond7_out),
    .reset(cond7_reset),
    .write_en(cond7_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire7 (
    .in(cond_wire7_in),
    .out(cond_wire7_out)
);
std_reg # (
    .WIDTH(1)
) cond8 (
    .clk(cond8_clk),
    .done(cond8_done),
    .in(cond8_in),
    .out(cond8_out),
    .reset(cond8_reset),
    .write_en(cond8_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire8 (
    .in(cond_wire8_in),
    .out(cond_wire8_out)
);
std_reg # (
    .WIDTH(1)
) cond9 (
    .clk(cond9_clk),
    .done(cond9_done),
    .in(cond9_in),
    .out(cond9_out),
    .reset(cond9_reset),
    .write_en(cond9_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire9 (
    .in(cond_wire9_in),
    .out(cond_wire9_out)
);
std_reg # (
    .WIDTH(1)
) cond10 (
    .clk(cond10_clk),
    .done(cond10_done),
    .in(cond10_in),
    .out(cond10_out),
    .reset(cond10_reset),
    .write_en(cond10_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire10 (
    .in(cond_wire10_in),
    .out(cond_wire10_out)
);
std_reg # (
    .WIDTH(1)
) cond11 (
    .clk(cond11_clk),
    .done(cond11_done),
    .in(cond11_in),
    .out(cond11_out),
    .reset(cond11_reset),
    .write_en(cond11_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire11 (
    .in(cond_wire11_in),
    .out(cond_wire11_out)
);
std_reg # (
    .WIDTH(1)
) cond12 (
    .clk(cond12_clk),
    .done(cond12_done),
    .in(cond12_in),
    .out(cond12_out),
    .reset(cond12_reset),
    .write_en(cond12_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire12 (
    .in(cond_wire12_in),
    .out(cond_wire12_out)
);
std_reg # (
    .WIDTH(1)
) cond13 (
    .clk(cond13_clk),
    .done(cond13_done),
    .in(cond13_in),
    .out(cond13_out),
    .reset(cond13_reset),
    .write_en(cond13_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire13 (
    .in(cond_wire13_in),
    .out(cond_wire13_out)
);
std_reg # (
    .WIDTH(1)
) cond14 (
    .clk(cond14_clk),
    .done(cond14_done),
    .in(cond14_in),
    .out(cond14_out),
    .reset(cond14_reset),
    .write_en(cond14_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire14 (
    .in(cond_wire14_in),
    .out(cond_wire14_out)
);
std_reg # (
    .WIDTH(1)
) cond15 (
    .clk(cond15_clk),
    .done(cond15_done),
    .in(cond15_in),
    .out(cond15_out),
    .reset(cond15_reset),
    .write_en(cond15_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire15 (
    .in(cond_wire15_in),
    .out(cond_wire15_out)
);
std_reg # (
    .WIDTH(1)
) cond16 (
    .clk(cond16_clk),
    .done(cond16_done),
    .in(cond16_in),
    .out(cond16_out),
    .reset(cond16_reset),
    .write_en(cond16_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire16 (
    .in(cond_wire16_in),
    .out(cond_wire16_out)
);
std_reg # (
    .WIDTH(1)
) cond17 (
    .clk(cond17_clk),
    .done(cond17_done),
    .in(cond17_in),
    .out(cond17_out),
    .reset(cond17_reset),
    .write_en(cond17_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire17 (
    .in(cond_wire17_in),
    .out(cond_wire17_out)
);
std_reg # (
    .WIDTH(1)
) cond18 (
    .clk(cond18_clk),
    .done(cond18_done),
    .in(cond18_in),
    .out(cond18_out),
    .reset(cond18_reset),
    .write_en(cond18_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire18 (
    .in(cond_wire18_in),
    .out(cond_wire18_out)
);
std_reg # (
    .WIDTH(1)
) cond19 (
    .clk(cond19_clk),
    .done(cond19_done),
    .in(cond19_in),
    .out(cond19_out),
    .reset(cond19_reset),
    .write_en(cond19_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire19 (
    .in(cond_wire19_in),
    .out(cond_wire19_out)
);
std_reg # (
    .WIDTH(1)
) cond20 (
    .clk(cond20_clk),
    .done(cond20_done),
    .in(cond20_in),
    .out(cond20_out),
    .reset(cond20_reset),
    .write_en(cond20_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire20 (
    .in(cond_wire20_in),
    .out(cond_wire20_out)
);
std_reg # (
    .WIDTH(1)
) cond21 (
    .clk(cond21_clk),
    .done(cond21_done),
    .in(cond21_in),
    .out(cond21_out),
    .reset(cond21_reset),
    .write_en(cond21_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire21 (
    .in(cond_wire21_in),
    .out(cond_wire21_out)
);
std_reg # (
    .WIDTH(1)
) cond22 (
    .clk(cond22_clk),
    .done(cond22_done),
    .in(cond22_in),
    .out(cond22_out),
    .reset(cond22_reset),
    .write_en(cond22_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire22 (
    .in(cond_wire22_in),
    .out(cond_wire22_out)
);
std_reg # (
    .WIDTH(1)
) cond23 (
    .clk(cond23_clk),
    .done(cond23_done),
    .in(cond23_in),
    .out(cond23_out),
    .reset(cond23_reset),
    .write_en(cond23_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire23 (
    .in(cond_wire23_in),
    .out(cond_wire23_out)
);
std_reg # (
    .WIDTH(1)
) cond24 (
    .clk(cond24_clk),
    .done(cond24_done),
    .in(cond24_in),
    .out(cond24_out),
    .reset(cond24_reset),
    .write_en(cond24_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire24 (
    .in(cond_wire24_in),
    .out(cond_wire24_out)
);
std_reg # (
    .WIDTH(1)
) cond25 (
    .clk(cond25_clk),
    .done(cond25_done),
    .in(cond25_in),
    .out(cond25_out),
    .reset(cond25_reset),
    .write_en(cond25_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire25 (
    .in(cond_wire25_in),
    .out(cond_wire25_out)
);
std_reg # (
    .WIDTH(1)
) cond26 (
    .clk(cond26_clk),
    .done(cond26_done),
    .in(cond26_in),
    .out(cond26_out),
    .reset(cond26_reset),
    .write_en(cond26_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire26 (
    .in(cond_wire26_in),
    .out(cond_wire26_out)
);
std_reg # (
    .WIDTH(1)
) cond27 (
    .clk(cond27_clk),
    .done(cond27_done),
    .in(cond27_in),
    .out(cond27_out),
    .reset(cond27_reset),
    .write_en(cond27_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire27 (
    .in(cond_wire27_in),
    .out(cond_wire27_out)
);
std_reg # (
    .WIDTH(1)
) cond28 (
    .clk(cond28_clk),
    .done(cond28_done),
    .in(cond28_in),
    .out(cond28_out),
    .reset(cond28_reset),
    .write_en(cond28_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire28 (
    .in(cond_wire28_in),
    .out(cond_wire28_out)
);
std_reg # (
    .WIDTH(1)
) cond29 (
    .clk(cond29_clk),
    .done(cond29_done),
    .in(cond29_in),
    .out(cond29_out),
    .reset(cond29_reset),
    .write_en(cond29_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire29 (
    .in(cond_wire29_in),
    .out(cond_wire29_out)
);
std_reg # (
    .WIDTH(1)
) cond30 (
    .clk(cond30_clk),
    .done(cond30_done),
    .in(cond30_in),
    .out(cond30_out),
    .reset(cond30_reset),
    .write_en(cond30_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire30 (
    .in(cond_wire30_in),
    .out(cond_wire30_out)
);
std_reg # (
    .WIDTH(1)
) cond31 (
    .clk(cond31_clk),
    .done(cond31_done),
    .in(cond31_in),
    .out(cond31_out),
    .reset(cond31_reset),
    .write_en(cond31_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire31 (
    .in(cond_wire31_in),
    .out(cond_wire31_out)
);
std_reg # (
    .WIDTH(1)
) cond32 (
    .clk(cond32_clk),
    .done(cond32_done),
    .in(cond32_in),
    .out(cond32_out),
    .reset(cond32_reset),
    .write_en(cond32_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire32 (
    .in(cond_wire32_in),
    .out(cond_wire32_out)
);
std_reg # (
    .WIDTH(1)
) cond33 (
    .clk(cond33_clk),
    .done(cond33_done),
    .in(cond33_in),
    .out(cond33_out),
    .reset(cond33_reset),
    .write_en(cond33_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire33 (
    .in(cond_wire33_in),
    .out(cond_wire33_out)
);
std_reg # (
    .WIDTH(1)
) cond34 (
    .clk(cond34_clk),
    .done(cond34_done),
    .in(cond34_in),
    .out(cond34_out),
    .reset(cond34_reset),
    .write_en(cond34_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire34 (
    .in(cond_wire34_in),
    .out(cond_wire34_out)
);
std_reg # (
    .WIDTH(1)
) cond35 (
    .clk(cond35_clk),
    .done(cond35_done),
    .in(cond35_in),
    .out(cond35_out),
    .reset(cond35_reset),
    .write_en(cond35_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire35 (
    .in(cond_wire35_in),
    .out(cond_wire35_out)
);
std_reg # (
    .WIDTH(1)
) cond36 (
    .clk(cond36_clk),
    .done(cond36_done),
    .in(cond36_in),
    .out(cond36_out),
    .reset(cond36_reset),
    .write_en(cond36_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire36 (
    .in(cond_wire36_in),
    .out(cond_wire36_out)
);
std_reg # (
    .WIDTH(1)
) cond37 (
    .clk(cond37_clk),
    .done(cond37_done),
    .in(cond37_in),
    .out(cond37_out),
    .reset(cond37_reset),
    .write_en(cond37_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire37 (
    .in(cond_wire37_in),
    .out(cond_wire37_out)
);
std_reg # (
    .WIDTH(1)
) cond38 (
    .clk(cond38_clk),
    .done(cond38_done),
    .in(cond38_in),
    .out(cond38_out),
    .reset(cond38_reset),
    .write_en(cond38_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire38 (
    .in(cond_wire38_in),
    .out(cond_wire38_out)
);
std_reg # (
    .WIDTH(1)
) cond39 (
    .clk(cond39_clk),
    .done(cond39_done),
    .in(cond39_in),
    .out(cond39_out),
    .reset(cond39_reset),
    .write_en(cond39_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire39 (
    .in(cond_wire39_in),
    .out(cond_wire39_out)
);
std_reg # (
    .WIDTH(1)
) cond40 (
    .clk(cond40_clk),
    .done(cond40_done),
    .in(cond40_in),
    .out(cond40_out),
    .reset(cond40_reset),
    .write_en(cond40_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire40 (
    .in(cond_wire40_in),
    .out(cond_wire40_out)
);
std_reg # (
    .WIDTH(1)
) cond41 (
    .clk(cond41_clk),
    .done(cond41_done),
    .in(cond41_in),
    .out(cond41_out),
    .reset(cond41_reset),
    .write_en(cond41_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire41 (
    .in(cond_wire41_in),
    .out(cond_wire41_out)
);
std_reg # (
    .WIDTH(1)
) cond42 (
    .clk(cond42_clk),
    .done(cond42_done),
    .in(cond42_in),
    .out(cond42_out),
    .reset(cond42_reset),
    .write_en(cond42_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire42 (
    .in(cond_wire42_in),
    .out(cond_wire42_out)
);
std_reg # (
    .WIDTH(1)
) cond43 (
    .clk(cond43_clk),
    .done(cond43_done),
    .in(cond43_in),
    .out(cond43_out),
    .reset(cond43_reset),
    .write_en(cond43_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire43 (
    .in(cond_wire43_in),
    .out(cond_wire43_out)
);
std_reg # (
    .WIDTH(1)
) cond44 (
    .clk(cond44_clk),
    .done(cond44_done),
    .in(cond44_in),
    .out(cond44_out),
    .reset(cond44_reset),
    .write_en(cond44_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire44 (
    .in(cond_wire44_in),
    .out(cond_wire44_out)
);
std_reg # (
    .WIDTH(1)
) cond45 (
    .clk(cond45_clk),
    .done(cond45_done),
    .in(cond45_in),
    .out(cond45_out),
    .reset(cond45_reset),
    .write_en(cond45_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire45 (
    .in(cond_wire45_in),
    .out(cond_wire45_out)
);
std_reg # (
    .WIDTH(1)
) cond46 (
    .clk(cond46_clk),
    .done(cond46_done),
    .in(cond46_in),
    .out(cond46_out),
    .reset(cond46_reset),
    .write_en(cond46_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire46 (
    .in(cond_wire46_in),
    .out(cond_wire46_out)
);
std_reg # (
    .WIDTH(1)
) cond47 (
    .clk(cond47_clk),
    .done(cond47_done),
    .in(cond47_in),
    .out(cond47_out),
    .reset(cond47_reset),
    .write_en(cond47_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire47 (
    .in(cond_wire47_in),
    .out(cond_wire47_out)
);
std_reg # (
    .WIDTH(1)
) cond48 (
    .clk(cond48_clk),
    .done(cond48_done),
    .in(cond48_in),
    .out(cond48_out),
    .reset(cond48_reset),
    .write_en(cond48_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire48 (
    .in(cond_wire48_in),
    .out(cond_wire48_out)
);
std_reg # (
    .WIDTH(1)
) cond49 (
    .clk(cond49_clk),
    .done(cond49_done),
    .in(cond49_in),
    .out(cond49_out),
    .reset(cond49_reset),
    .write_en(cond49_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire49 (
    .in(cond_wire49_in),
    .out(cond_wire49_out)
);
std_reg # (
    .WIDTH(1)
) cond50 (
    .clk(cond50_clk),
    .done(cond50_done),
    .in(cond50_in),
    .out(cond50_out),
    .reset(cond50_reset),
    .write_en(cond50_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire50 (
    .in(cond_wire50_in),
    .out(cond_wire50_out)
);
std_reg # (
    .WIDTH(1)
) cond51 (
    .clk(cond51_clk),
    .done(cond51_done),
    .in(cond51_in),
    .out(cond51_out),
    .reset(cond51_reset),
    .write_en(cond51_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire51 (
    .in(cond_wire51_in),
    .out(cond_wire51_out)
);
std_reg # (
    .WIDTH(1)
) cond52 (
    .clk(cond52_clk),
    .done(cond52_done),
    .in(cond52_in),
    .out(cond52_out),
    .reset(cond52_reset),
    .write_en(cond52_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire52 (
    .in(cond_wire52_in),
    .out(cond_wire52_out)
);
std_reg # (
    .WIDTH(1)
) cond53 (
    .clk(cond53_clk),
    .done(cond53_done),
    .in(cond53_in),
    .out(cond53_out),
    .reset(cond53_reset),
    .write_en(cond53_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire53 (
    .in(cond_wire53_in),
    .out(cond_wire53_out)
);
std_reg # (
    .WIDTH(1)
) cond54 (
    .clk(cond54_clk),
    .done(cond54_done),
    .in(cond54_in),
    .out(cond54_out),
    .reset(cond54_reset),
    .write_en(cond54_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire54 (
    .in(cond_wire54_in),
    .out(cond_wire54_out)
);
std_reg # (
    .WIDTH(1)
) cond55 (
    .clk(cond55_clk),
    .done(cond55_done),
    .in(cond55_in),
    .out(cond55_out),
    .reset(cond55_reset),
    .write_en(cond55_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire55 (
    .in(cond_wire55_in),
    .out(cond_wire55_out)
);
std_reg # (
    .WIDTH(1)
) cond56 (
    .clk(cond56_clk),
    .done(cond56_done),
    .in(cond56_in),
    .out(cond56_out),
    .reset(cond56_reset),
    .write_en(cond56_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire56 (
    .in(cond_wire56_in),
    .out(cond_wire56_out)
);
std_reg # (
    .WIDTH(1)
) cond57 (
    .clk(cond57_clk),
    .done(cond57_done),
    .in(cond57_in),
    .out(cond57_out),
    .reset(cond57_reset),
    .write_en(cond57_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire57 (
    .in(cond_wire57_in),
    .out(cond_wire57_out)
);
std_reg # (
    .WIDTH(1)
) cond58 (
    .clk(cond58_clk),
    .done(cond58_done),
    .in(cond58_in),
    .out(cond58_out),
    .reset(cond58_reset),
    .write_en(cond58_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire58 (
    .in(cond_wire58_in),
    .out(cond_wire58_out)
);
std_reg # (
    .WIDTH(1)
) cond59 (
    .clk(cond59_clk),
    .done(cond59_done),
    .in(cond59_in),
    .out(cond59_out),
    .reset(cond59_reset),
    .write_en(cond59_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire59 (
    .in(cond_wire59_in),
    .out(cond_wire59_out)
);
std_reg # (
    .WIDTH(1)
) cond60 (
    .clk(cond60_clk),
    .done(cond60_done),
    .in(cond60_in),
    .out(cond60_out),
    .reset(cond60_reset),
    .write_en(cond60_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire60 (
    .in(cond_wire60_in),
    .out(cond_wire60_out)
);
std_reg # (
    .WIDTH(1)
) cond61 (
    .clk(cond61_clk),
    .done(cond61_done),
    .in(cond61_in),
    .out(cond61_out),
    .reset(cond61_reset),
    .write_en(cond61_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire61 (
    .in(cond_wire61_in),
    .out(cond_wire61_out)
);
std_reg # (
    .WIDTH(1)
) cond62 (
    .clk(cond62_clk),
    .done(cond62_done),
    .in(cond62_in),
    .out(cond62_out),
    .reset(cond62_reset),
    .write_en(cond62_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire62 (
    .in(cond_wire62_in),
    .out(cond_wire62_out)
);
std_reg # (
    .WIDTH(1)
) cond63 (
    .clk(cond63_clk),
    .done(cond63_done),
    .in(cond63_in),
    .out(cond63_out),
    .reset(cond63_reset),
    .write_en(cond63_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire63 (
    .in(cond_wire63_in),
    .out(cond_wire63_out)
);
std_reg # (
    .WIDTH(1)
) cond64 (
    .clk(cond64_clk),
    .done(cond64_done),
    .in(cond64_in),
    .out(cond64_out),
    .reset(cond64_reset),
    .write_en(cond64_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire64 (
    .in(cond_wire64_in),
    .out(cond_wire64_out)
);
std_reg # (
    .WIDTH(1)
) cond65 (
    .clk(cond65_clk),
    .done(cond65_done),
    .in(cond65_in),
    .out(cond65_out),
    .reset(cond65_reset),
    .write_en(cond65_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire65 (
    .in(cond_wire65_in),
    .out(cond_wire65_out)
);
std_reg # (
    .WIDTH(1)
) cond66 (
    .clk(cond66_clk),
    .done(cond66_done),
    .in(cond66_in),
    .out(cond66_out),
    .reset(cond66_reset),
    .write_en(cond66_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire66 (
    .in(cond_wire66_in),
    .out(cond_wire66_out)
);
std_reg # (
    .WIDTH(1)
) cond67 (
    .clk(cond67_clk),
    .done(cond67_done),
    .in(cond67_in),
    .out(cond67_out),
    .reset(cond67_reset),
    .write_en(cond67_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire67 (
    .in(cond_wire67_in),
    .out(cond_wire67_out)
);
std_reg # (
    .WIDTH(1)
) cond68 (
    .clk(cond68_clk),
    .done(cond68_done),
    .in(cond68_in),
    .out(cond68_out),
    .reset(cond68_reset),
    .write_en(cond68_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire68 (
    .in(cond_wire68_in),
    .out(cond_wire68_out)
);
std_reg # (
    .WIDTH(1)
) fsm (
    .clk(fsm_clk),
    .done(fsm_done),
    .in(fsm_in),
    .out(fsm_out),
    .reset(fsm_reset),
    .write_en(fsm_write_en)
);
undef # (
    .WIDTH(1)
) ud (
    .out(ud_out)
);
std_add # (
    .WIDTH(1)
) adder (
    .left(adder_left),
    .out(adder_out),
    .right(adder_right)
);
undef # (
    .WIDTH(1)
) ud0 (
    .out(ud0_out)
);
std_add # (
    .WIDTH(1)
) adder0 (
    .left(adder0_left),
    .out(adder0_out),
    .right(adder0_right)
);
std_reg # (
    .WIDTH(1)
) signal_reg (
    .clk(signal_reg_clk),
    .done(signal_reg_done),
    .in(signal_reg_in),
    .out(signal_reg_out),
    .reset(signal_reg_reset),
    .write_en(signal_reg_write_en)
);
std_reg # (
    .WIDTH(2)
) fsm0 (
    .clk(fsm0_clk),
    .done(fsm0_done),
    .in(fsm0_in),
    .out(fsm0_out),
    .reset(fsm0_reset),
    .write_en(fsm0_write_en)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_go (
    .in(early_reset_static_par_go_in),
    .out(early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_done (
    .in(early_reset_static_par_done_in),
    .out(early_reset_static_par_done_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par0_go (
    .in(early_reset_static_par0_go_in),
    .out(early_reset_static_par0_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par0_done (
    .in(early_reset_static_par0_done_in),
    .out(early_reset_static_par0_done_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_go (
    .in(wrapper_early_reset_static_par_go_in),
    .out(wrapper_early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_done (
    .in(wrapper_early_reset_static_par_done_in),
    .out(wrapper_early_reset_static_par_done_out)
);
std_wire # (
    .WIDTH(1)
) while_wrapper_early_reset_static_par0_go (
    .in(while_wrapper_early_reset_static_par0_go_in),
    .out(while_wrapper_early_reset_static_par0_go_out)
);
std_wire # (
    .WIDTH(1)
) while_wrapper_early_reset_static_par0_done (
    .in(while_wrapper_early_reset_static_par0_done_in),
    .out(while_wrapper_early_reset_static_par0_done_out)
);
std_wire # (
    .WIDTH(1)
) tdcc_go (
    .in(tdcc_go_in),
    .out(tdcc_go_out)
);
std_wire # (
    .WIDTH(1)
) tdcc_done (
    .in(tdcc_done_in),
    .out(tdcc_done_out)
);
wire _guard0 = 1;
wire _guard1 = early_reset_static_par0_go_out;
wire _guard2 = early_reset_static_par0_go_out;
wire _guard3 = cond_wire14_out;
wire _guard4 = early_reset_static_par0_go_out;
wire _guard5 = _guard3 & _guard4;
wire _guard6 = cond_wire14_out;
wire _guard7 = early_reset_static_par0_go_out;
wire _guard8 = _guard6 & _guard7;
wire _guard9 = cond_wire19_out;
wire _guard10 = early_reset_static_par0_go_out;
wire _guard11 = _guard9 & _guard10;
wire _guard12 = cond_wire19_out;
wire _guard13 = early_reset_static_par0_go_out;
wire _guard14 = _guard12 & _guard13;
wire _guard15 = early_reset_static_par_go_out;
wire _guard16 = early_reset_static_par0_go_out;
wire _guard17 = _guard15 | _guard16;
wire _guard18 = early_reset_static_par0_go_out;
wire _guard19 = early_reset_static_par_go_out;
wire _guard20 = early_reset_static_par_go_out;
wire _guard21 = early_reset_static_par0_go_out;
wire _guard22 = _guard20 | _guard21;
wire _guard23 = early_reset_static_par0_go_out;
wire _guard24 = early_reset_static_par_go_out;
wire _guard25 = early_reset_static_par0_go_out;
wire _guard26 = ~_guard0;
wire _guard27 = early_reset_static_par0_go_out;
wire _guard28 = _guard26 & _guard27;
wire _guard29 = ~_guard0;
wire _guard30 = early_reset_static_par0_go_out;
wire _guard31 = _guard29 & _guard30;
wire _guard32 = early_reset_static_par0_go_out;
wire _guard33 = early_reset_static_par0_go_out;
wire _guard34 = ~_guard0;
wire _guard35 = early_reset_static_par0_go_out;
wire _guard36 = _guard34 & _guard35;
wire _guard37 = early_reset_static_par0_go_out;
wire _guard38 = ~_guard0;
wire _guard39 = early_reset_static_par0_go_out;
wire _guard40 = _guard38 & _guard39;
wire _guard41 = early_reset_static_par0_go_out;
wire _guard42 = ~_guard0;
wire _guard43 = early_reset_static_par0_go_out;
wire _guard44 = _guard42 & _guard43;
wire _guard45 = early_reset_static_par0_go_out;
wire _guard46 = early_reset_static_par0_go_out;
wire _guard47 = ~_guard0;
wire _guard48 = early_reset_static_par0_go_out;
wire _guard49 = _guard47 & _guard48;
wire _guard50 = early_reset_static_par0_go_out;
wire _guard51 = early_reset_static_par0_go_out;
wire _guard52 = early_reset_static_par0_go_out;
wire _guard53 = cond_wire11_out;
wire _guard54 = early_reset_static_par0_go_out;
wire _guard55 = _guard53 & _guard54;
wire _guard56 = cond_wire11_out;
wire _guard57 = early_reset_static_par0_go_out;
wire _guard58 = _guard56 & _guard57;
wire _guard59 = cond_wire1_out;
wire _guard60 = early_reset_static_par0_go_out;
wire _guard61 = _guard59 & _guard60;
wire _guard62 = cond_wire1_out;
wire _guard63 = early_reset_static_par0_go_out;
wire _guard64 = _guard62 & _guard63;
wire _guard65 = cond_wire30_out;
wire _guard66 = early_reset_static_par0_go_out;
wire _guard67 = _guard65 & _guard66;
wire _guard68 = cond_wire28_out;
wire _guard69 = early_reset_static_par0_go_out;
wire _guard70 = _guard68 & _guard69;
wire _guard71 = fsm_out == 1'd0;
wire _guard72 = cond_wire28_out;
wire _guard73 = _guard71 & _guard72;
wire _guard74 = fsm_out == 1'd0;
wire _guard75 = _guard73 & _guard74;
wire _guard76 = fsm_out == 1'd0;
wire _guard77 = cond_wire30_out;
wire _guard78 = _guard76 & _guard77;
wire _guard79 = fsm_out == 1'd0;
wire _guard80 = _guard78 & _guard79;
wire _guard81 = _guard75 | _guard80;
wire _guard82 = early_reset_static_par0_go_out;
wire _guard83 = _guard81 & _guard82;
wire _guard84 = fsm_out == 1'd0;
wire _guard85 = cond_wire28_out;
wire _guard86 = _guard84 & _guard85;
wire _guard87 = fsm_out == 1'd0;
wire _guard88 = _guard86 & _guard87;
wire _guard89 = fsm_out == 1'd0;
wire _guard90 = cond_wire30_out;
wire _guard91 = _guard89 & _guard90;
wire _guard92 = fsm_out == 1'd0;
wire _guard93 = _guard91 & _guard92;
wire _guard94 = _guard88 | _guard93;
wire _guard95 = early_reset_static_par0_go_out;
wire _guard96 = _guard94 & _guard95;
wire _guard97 = fsm_out == 1'd0;
wire _guard98 = cond_wire28_out;
wire _guard99 = _guard97 & _guard98;
wire _guard100 = fsm_out == 1'd0;
wire _guard101 = _guard99 & _guard100;
wire _guard102 = fsm_out == 1'd0;
wire _guard103 = cond_wire30_out;
wire _guard104 = _guard102 & _guard103;
wire _guard105 = fsm_out == 1'd0;
wire _guard106 = _guard104 & _guard105;
wire _guard107 = _guard101 | _guard106;
wire _guard108 = early_reset_static_par0_go_out;
wire _guard109 = _guard107 & _guard108;
wire _guard110 = cond_wire34_out;
wire _guard111 = early_reset_static_par0_go_out;
wire _guard112 = _guard110 & _guard111;
wire _guard113 = cond_wire32_out;
wire _guard114 = early_reset_static_par0_go_out;
wire _guard115 = _guard113 & _guard114;
wire _guard116 = fsm_out == 1'd0;
wire _guard117 = cond_wire32_out;
wire _guard118 = _guard116 & _guard117;
wire _guard119 = fsm_out == 1'd0;
wire _guard120 = _guard118 & _guard119;
wire _guard121 = fsm_out == 1'd0;
wire _guard122 = cond_wire34_out;
wire _guard123 = _guard121 & _guard122;
wire _guard124 = fsm_out == 1'd0;
wire _guard125 = _guard123 & _guard124;
wire _guard126 = _guard120 | _guard125;
wire _guard127 = early_reset_static_par0_go_out;
wire _guard128 = _guard126 & _guard127;
wire _guard129 = fsm_out == 1'd0;
wire _guard130 = cond_wire32_out;
wire _guard131 = _guard129 & _guard130;
wire _guard132 = fsm_out == 1'd0;
wire _guard133 = _guard131 & _guard132;
wire _guard134 = fsm_out == 1'd0;
wire _guard135 = cond_wire34_out;
wire _guard136 = _guard134 & _guard135;
wire _guard137 = fsm_out == 1'd0;
wire _guard138 = _guard136 & _guard137;
wire _guard139 = _guard133 | _guard138;
wire _guard140 = early_reset_static_par0_go_out;
wire _guard141 = _guard139 & _guard140;
wire _guard142 = fsm_out == 1'd0;
wire _guard143 = cond_wire32_out;
wire _guard144 = _guard142 & _guard143;
wire _guard145 = fsm_out == 1'd0;
wire _guard146 = _guard144 & _guard145;
wire _guard147 = fsm_out == 1'd0;
wire _guard148 = cond_wire34_out;
wire _guard149 = _guard147 & _guard148;
wire _guard150 = fsm_out == 1'd0;
wire _guard151 = _guard149 & _guard150;
wire _guard152 = _guard146 | _guard151;
wire _guard153 = early_reset_static_par0_go_out;
wire _guard154 = _guard152 & _guard153;
wire _guard155 = cond_wire29_out;
wire _guard156 = early_reset_static_par0_go_out;
wire _guard157 = _guard155 & _guard156;
wire _guard158 = cond_wire29_out;
wire _guard159 = early_reset_static_par0_go_out;
wire _guard160 = _guard158 & _guard159;
wire _guard161 = early_reset_static_par_go_out;
wire _guard162 = cond_wire53_out;
wire _guard163 = early_reset_static_par0_go_out;
wire _guard164 = _guard162 & _guard163;
wire _guard165 = _guard161 | _guard164;
wire _guard166 = cond_wire53_out;
wire _guard167 = early_reset_static_par0_go_out;
wire _guard168 = _guard166 & _guard167;
wire _guard169 = early_reset_static_par_go_out;
wire _guard170 = early_reset_static_par0_go_out;
wire _guard171 = early_reset_static_par0_go_out;
wire _guard172 = early_reset_static_par0_go_out;
wire _guard173 = early_reset_static_par0_go_out;
wire _guard174 = early_reset_static_par0_go_out;
wire _guard175 = early_reset_static_par0_go_out;
wire _guard176 = early_reset_static_par0_go_out;
wire _guard177 = early_reset_static_par0_go_out;
wire _guard178 = early_reset_static_par0_go_out;
wire _guard179 = early_reset_static_par0_go_out;
wire _guard180 = early_reset_static_par_go_out;
wire _guard181 = early_reset_static_par0_go_out;
wire _guard182 = _guard180 | _guard181;
wire _guard183 = early_reset_static_par0_go_out;
wire _guard184 = early_reset_static_par_go_out;
wire _guard185 = cond_wire9_out;
wire _guard186 = early_reset_static_par0_go_out;
wire _guard187 = _guard185 & _guard186;
wire _guard188 = tdcc_done_out;
wire _guard189 = cond_wire_out;
wire _guard190 = early_reset_static_par0_go_out;
wire _guard191 = _guard189 & _guard190;
wire _guard192 = cond_wire23_out;
wire _guard193 = early_reset_static_par0_go_out;
wire _guard194 = _guard192 & _guard193;
wire _guard195 = cond_wire31_out;
wire _guard196 = early_reset_static_par0_go_out;
wire _guard197 = _guard195 & _guard196;
wire _guard198 = cond_wire27_out;
wire _guard199 = early_reset_static_par0_go_out;
wire _guard200 = _guard198 & _guard199;
wire _guard201 = cond_wire35_out;
wire _guard202 = early_reset_static_par0_go_out;
wire _guard203 = _guard201 & _guard202;
wire _guard204 = cond_wire8_out;
wire _guard205 = early_reset_static_par0_go_out;
wire _guard206 = _guard204 & _guard205;
wire _guard207 = cond_wire18_out;
wire _guard208 = early_reset_static_par0_go_out;
wire _guard209 = _guard207 & _guard208;
wire _guard210 = cond_wire13_out;
wire _guard211 = early_reset_static_par0_go_out;
wire _guard212 = _guard210 & _guard211;
wire _guard213 = cond_wire3_out;
wire _guard214 = early_reset_static_par0_go_out;
wire _guard215 = _guard213 & _guard214;
wire _guard216 = cond_wire65_out;
wire _guard217 = early_reset_static_par0_go_out;
wire _guard218 = _guard216 & _guard217;
wire _guard219 = cond_wire57_out;
wire _guard220 = early_reset_static_par0_go_out;
wire _guard221 = _guard219 & _guard220;
wire _guard222 = cond_wire61_out;
wire _guard223 = early_reset_static_par0_go_out;
wire _guard224 = _guard222 & _guard223;
wire _guard225 = cond_wire68_out;
wire _guard226 = early_reset_static_par0_go_out;
wire _guard227 = _guard225 & _guard226;
wire _guard228 = cond_wire19_out;
wire _guard229 = early_reset_static_par0_go_out;
wire _guard230 = _guard228 & _guard229;
wire _guard231 = cond_wire53_out;
wire _guard232 = early_reset_static_par0_go_out;
wire _guard233 = _guard231 & _guard232;
wire _guard234 = cond_wire44_out;
wire _guard235 = early_reset_static_par0_go_out;
wire _guard236 = _guard234 & _guard235;
wire _guard237 = cond_wire52_out;
wire _guard238 = early_reset_static_par0_go_out;
wire _guard239 = _guard237 & _guard238;
wire _guard240 = cond_wire40_out;
wire _guard241 = early_reset_static_par0_go_out;
wire _guard242 = _guard240 & _guard241;
wire _guard243 = cond_wire48_out;
wire _guard244 = early_reset_static_par0_go_out;
wire _guard245 = _guard243 & _guard244;
wire _guard246 = cond_wire31_out;
wire _guard247 = early_reset_static_par0_go_out;
wire _guard248 = _guard246 & _guard247;
wire _guard249 = cond_wire35_out;
wire _guard250 = early_reset_static_par0_go_out;
wire _guard251 = _guard249 & _guard250;
wire _guard252 = cond_wire23_out;
wire _guard253 = early_reset_static_par0_go_out;
wire _guard254 = _guard252 & _guard253;
wire _guard255 = cond_wire27_out;
wire _guard256 = early_reset_static_par0_go_out;
wire _guard257 = _guard255 & _guard256;
wire _guard258 = fsm_out == 1'd0;
wire _guard259 = cond_wire23_out;
wire _guard260 = _guard258 & _guard259;
wire _guard261 = fsm_out == 1'd0;
wire _guard262 = _guard260 & _guard261;
wire _guard263 = fsm_out == 1'd0;
wire _guard264 = cond_wire27_out;
wire _guard265 = _guard263 & _guard264;
wire _guard266 = fsm_out == 1'd0;
wire _guard267 = _guard265 & _guard266;
wire _guard268 = _guard262 | _guard267;
wire _guard269 = fsm_out == 1'd0;
wire _guard270 = cond_wire31_out;
wire _guard271 = _guard269 & _guard270;
wire _guard272 = fsm_out == 1'd0;
wire _guard273 = _guard271 & _guard272;
wire _guard274 = _guard268 | _guard273;
wire _guard275 = fsm_out == 1'd0;
wire _guard276 = cond_wire35_out;
wire _guard277 = _guard275 & _guard276;
wire _guard278 = fsm_out == 1'd0;
wire _guard279 = _guard277 & _guard278;
wire _guard280 = _guard274 | _guard279;
wire _guard281 = early_reset_static_par0_go_out;
wire _guard282 = _guard280 & _guard281;
wire _guard283 = cond_wire_out;
wire _guard284 = early_reset_static_par0_go_out;
wire _guard285 = _guard283 & _guard284;
wire _guard286 = cond_wire4_out;
wire _guard287 = early_reset_static_par0_go_out;
wire _guard288 = _guard286 & _guard287;
wire _guard289 = fsm_out == 1'd0;
wire _guard290 = cond_wire3_out;
wire _guard291 = _guard289 & _guard290;
wire _guard292 = fsm_out == 1'd0;
wire _guard293 = _guard291 & _guard292;
wire _guard294 = fsm_out == 1'd0;
wire _guard295 = cond_wire8_out;
wire _guard296 = _guard294 & _guard295;
wire _guard297 = fsm_out == 1'd0;
wire _guard298 = _guard296 & _guard297;
wire _guard299 = _guard293 | _guard298;
wire _guard300 = fsm_out == 1'd0;
wire _guard301 = cond_wire13_out;
wire _guard302 = _guard300 & _guard301;
wire _guard303 = fsm_out == 1'd0;
wire _guard304 = _guard302 & _guard303;
wire _guard305 = _guard299 | _guard304;
wire _guard306 = fsm_out == 1'd0;
wire _guard307 = cond_wire18_out;
wire _guard308 = _guard306 & _guard307;
wire _guard309 = fsm_out == 1'd0;
wire _guard310 = _guard308 & _guard309;
wire _guard311 = _guard305 | _guard310;
wire _guard312 = early_reset_static_par0_go_out;
wire _guard313 = _guard311 & _guard312;
wire _guard314 = fsm_out == 1'd0;
wire _guard315 = cond_wire40_out;
wire _guard316 = _guard314 & _guard315;
wire _guard317 = fsm_out == 1'd0;
wire _guard318 = _guard316 & _guard317;
wire _guard319 = fsm_out == 1'd0;
wire _guard320 = cond_wire44_out;
wire _guard321 = _guard319 & _guard320;
wire _guard322 = fsm_out == 1'd0;
wire _guard323 = _guard321 & _guard322;
wire _guard324 = _guard318 | _guard323;
wire _guard325 = fsm_out == 1'd0;
wire _guard326 = cond_wire48_out;
wire _guard327 = _guard325 & _guard326;
wire _guard328 = fsm_out == 1'd0;
wire _guard329 = _guard327 & _guard328;
wire _guard330 = _guard324 | _guard329;
wire _guard331 = fsm_out == 1'd0;
wire _guard332 = cond_wire52_out;
wire _guard333 = _guard331 & _guard332;
wire _guard334 = fsm_out == 1'd0;
wire _guard335 = _guard333 & _guard334;
wire _guard336 = _guard330 | _guard335;
wire _guard337 = early_reset_static_par0_go_out;
wire _guard338 = _guard336 & _guard337;
wire _guard339 = fsm_out == 1'd0;
wire _guard340 = cond_wire57_out;
wire _guard341 = _guard339 & _guard340;
wire _guard342 = fsm_out == 1'd0;
wire _guard343 = _guard341 & _guard342;
wire _guard344 = fsm_out == 1'd0;
wire _guard345 = cond_wire61_out;
wire _guard346 = _guard344 & _guard345;
wire _guard347 = fsm_out == 1'd0;
wire _guard348 = _guard346 & _guard347;
wire _guard349 = _guard343 | _guard348;
wire _guard350 = fsm_out == 1'd0;
wire _guard351 = cond_wire65_out;
wire _guard352 = _guard350 & _guard351;
wire _guard353 = fsm_out == 1'd0;
wire _guard354 = _guard352 & _guard353;
wire _guard355 = _guard349 | _guard354;
wire _guard356 = fsm_out == 1'd0;
wire _guard357 = cond_wire68_out;
wire _guard358 = _guard356 & _guard357;
wire _guard359 = fsm_out == 1'd0;
wire _guard360 = _guard358 & _guard359;
wire _guard361 = _guard355 | _guard360;
wire _guard362 = early_reset_static_par0_go_out;
wire _guard363 = _guard361 & _guard362;
wire _guard364 = cond_wire36_out;
wire _guard365 = early_reset_static_par0_go_out;
wire _guard366 = _guard364 & _guard365;
wire _guard367 = cond_wire3_out;
wire _guard368 = early_reset_static_par0_go_out;
wire _guard369 = _guard367 & _guard368;
wire _guard370 = cond_wire13_out;
wire _guard371 = early_reset_static_par0_go_out;
wire _guard372 = _guard370 & _guard371;
wire _guard373 = cond_wire8_out;
wire _guard374 = early_reset_static_par0_go_out;
wire _guard375 = _guard373 & _guard374;
wire _guard376 = cond_wire18_out;
wire _guard377 = early_reset_static_par0_go_out;
wire _guard378 = _guard376 & _guard377;
wire _guard379 = cond_wire57_out;
wire _guard380 = early_reset_static_par0_go_out;
wire _guard381 = _guard379 & _guard380;
wire _guard382 = cond_wire65_out;
wire _guard383 = early_reset_static_par0_go_out;
wire _guard384 = _guard382 & _guard383;
wire _guard385 = cond_wire61_out;
wire _guard386 = early_reset_static_par0_go_out;
wire _guard387 = _guard385 & _guard386;
wire _guard388 = cond_wire68_out;
wire _guard389 = early_reset_static_par0_go_out;
wire _guard390 = _guard388 & _guard389;
wire _guard391 = cond_wire14_out;
wire _guard392 = early_reset_static_par0_go_out;
wire _guard393 = _guard391 & _guard392;
wire _guard394 = cond_wire40_out;
wire _guard395 = early_reset_static_par0_go_out;
wire _guard396 = _guard394 & _guard395;
wire _guard397 = cond_wire48_out;
wire _guard398 = early_reset_static_par0_go_out;
wire _guard399 = _guard397 & _guard398;
wire _guard400 = cond_wire44_out;
wire _guard401 = early_reset_static_par0_go_out;
wire _guard402 = _guard400 & _guard401;
wire _guard403 = cond_wire52_out;
wire _guard404 = early_reset_static_par0_go_out;
wire _guard405 = _guard403 & _guard404;
wire _guard406 = early_reset_static_par0_go_out;
wire _guard407 = ~_guard0;
wire _guard408 = early_reset_static_par0_go_out;
wire _guard409 = _guard407 & _guard408;
wire _guard410 = ~_guard0;
wire _guard411 = early_reset_static_par0_go_out;
wire _guard412 = _guard410 & _guard411;
wire _guard413 = early_reset_static_par0_go_out;
wire _guard414 = early_reset_static_par0_go_out;
wire _guard415 = early_reset_static_par0_go_out;
wire _guard416 = ~_guard0;
wire _guard417 = early_reset_static_par0_go_out;
wire _guard418 = _guard416 & _guard417;
wire _guard419 = early_reset_static_par0_go_out;
wire _guard420 = ~_guard0;
wire _guard421 = early_reset_static_par0_go_out;
wire _guard422 = _guard420 & _guard421;
wire _guard423 = early_reset_static_par0_go_out;
wire _guard424 = early_reset_static_par0_go_out;
wire _guard425 = early_reset_static_par0_go_out;
wire _guard426 = ~_guard0;
wire _guard427 = early_reset_static_par0_go_out;
wire _guard428 = _guard426 & _guard427;
wire _guard429 = early_reset_static_par0_go_out;
wire _guard430 = ~_guard0;
wire _guard431 = early_reset_static_par0_go_out;
wire _guard432 = _guard430 & _guard431;
wire _guard433 = early_reset_static_par0_go_out;
wire _guard434 = early_reset_static_par0_go_out;
wire _guard435 = early_reset_static_par0_go_out;
wire _guard436 = early_reset_static_par0_go_out;
wire _guard437 = early_reset_static_par0_go_out;
wire _guard438 = early_reset_static_par_go_out;
wire _guard439 = early_reset_static_par0_go_out;
wire _guard440 = _guard438 | _guard439;
wire _guard441 = fsm_out != 1'd0;
wire _guard442 = early_reset_static_par_go_out;
wire _guard443 = _guard441 & _guard442;
wire _guard444 = fsm_out == 1'd0;
wire _guard445 = early_reset_static_par_go_out;
wire _guard446 = _guard444 & _guard445;
wire _guard447 = fsm_out == 1'd0;
wire _guard448 = early_reset_static_par0_go_out;
wire _guard449 = _guard447 & _guard448;
wire _guard450 = _guard446 | _guard449;
wire _guard451 = fsm_out != 1'd0;
wire _guard452 = early_reset_static_par0_go_out;
wire _guard453 = _guard451 & _guard452;
wire _guard454 = early_reset_static_par_go_out;
wire _guard455 = early_reset_static_par_go_out;
wire _guard456 = while_wrapper_early_reset_static_par0_go_out;
wire _guard457 = early_reset_static_par0_go_out;
wire _guard458 = early_reset_static_par0_go_out;
wire _guard459 = early_reset_static_par0_go_out;
wire _guard460 = early_reset_static_par0_go_out;
wire _guard461 = early_reset_static_par_go_out;
wire _guard462 = cond_wire_out;
wire _guard463 = early_reset_static_par0_go_out;
wire _guard464 = _guard462 & _guard463;
wire _guard465 = _guard461 | _guard464;
wire _guard466 = cond_wire_out;
wire _guard467 = early_reset_static_par0_go_out;
wire _guard468 = _guard466 & _guard467;
wire _guard469 = early_reset_static_par_go_out;
wire _guard470 = early_reset_static_par0_go_out;
wire _guard471 = early_reset_static_par0_go_out;
wire _guard472 = early_reset_static_par0_go_out;
wire _guard473 = early_reset_static_par0_go_out;
wire _guard474 = early_reset_static_par_go_out;
wire _guard475 = early_reset_static_par0_go_out;
wire _guard476 = _guard474 | _guard475;
wire _guard477 = early_reset_static_par_go_out;
wire _guard478 = early_reset_static_par0_go_out;
wire _guard479 = early_reset_static_par0_go_out;
wire _guard480 = early_reset_static_par0_go_out;
wire _guard481 = early_reset_static_par0_go_out;
wire _guard482 = early_reset_static_par0_go_out;
wire _guard483 = ~_guard0;
wire _guard484 = early_reset_static_par0_go_out;
wire _guard485 = _guard483 & _guard484;
wire _guard486 = early_reset_static_par0_go_out;
wire _guard487 = early_reset_static_par0_go_out;
wire _guard488 = early_reset_static_par0_go_out;
wire _guard489 = ~_guard0;
wire _guard490 = early_reset_static_par0_go_out;
wire _guard491 = _guard489 & _guard490;
wire _guard492 = early_reset_static_par0_go_out;
wire _guard493 = early_reset_static_par0_go_out;
wire _guard494 = ~_guard0;
wire _guard495 = early_reset_static_par0_go_out;
wire _guard496 = _guard494 & _guard495;
wire _guard497 = early_reset_static_par0_go_out;
wire _guard498 = early_reset_static_par0_go_out;
wire _guard499 = ~_guard0;
wire _guard500 = early_reset_static_par0_go_out;
wire _guard501 = _guard499 & _guard500;
wire _guard502 = early_reset_static_par0_go_out;
wire _guard503 = early_reset_static_par0_go_out;
wire _guard504 = ~_guard0;
wire _guard505 = early_reset_static_par0_go_out;
wire _guard506 = _guard504 & _guard505;
wire _guard507 = cond_wire7_out;
wire _guard508 = early_reset_static_par0_go_out;
wire _guard509 = _guard507 & _guard508;
wire _guard510 = cond_wire5_out;
wire _guard511 = early_reset_static_par0_go_out;
wire _guard512 = _guard510 & _guard511;
wire _guard513 = fsm_out == 1'd0;
wire _guard514 = cond_wire5_out;
wire _guard515 = _guard513 & _guard514;
wire _guard516 = fsm_out == 1'd0;
wire _guard517 = _guard515 & _guard516;
wire _guard518 = fsm_out == 1'd0;
wire _guard519 = cond_wire7_out;
wire _guard520 = _guard518 & _guard519;
wire _guard521 = fsm_out == 1'd0;
wire _guard522 = _guard520 & _guard521;
wire _guard523 = _guard517 | _guard522;
wire _guard524 = early_reset_static_par0_go_out;
wire _guard525 = _guard523 & _guard524;
wire _guard526 = fsm_out == 1'd0;
wire _guard527 = cond_wire5_out;
wire _guard528 = _guard526 & _guard527;
wire _guard529 = fsm_out == 1'd0;
wire _guard530 = _guard528 & _guard529;
wire _guard531 = fsm_out == 1'd0;
wire _guard532 = cond_wire7_out;
wire _guard533 = _guard531 & _guard532;
wire _guard534 = fsm_out == 1'd0;
wire _guard535 = _guard533 & _guard534;
wire _guard536 = _guard530 | _guard535;
wire _guard537 = early_reset_static_par0_go_out;
wire _guard538 = _guard536 & _guard537;
wire _guard539 = fsm_out == 1'd0;
wire _guard540 = cond_wire5_out;
wire _guard541 = _guard539 & _guard540;
wire _guard542 = fsm_out == 1'd0;
wire _guard543 = _guard541 & _guard542;
wire _guard544 = fsm_out == 1'd0;
wire _guard545 = cond_wire7_out;
wire _guard546 = _guard544 & _guard545;
wire _guard547 = fsm_out == 1'd0;
wire _guard548 = _guard546 & _guard547;
wire _guard549 = _guard543 | _guard548;
wire _guard550 = early_reset_static_par0_go_out;
wire _guard551 = _guard549 & _guard550;
wire _guard552 = cond_wire25_out;
wire _guard553 = early_reset_static_par0_go_out;
wire _guard554 = _guard552 & _guard553;
wire _guard555 = cond_wire25_out;
wire _guard556 = early_reset_static_par0_go_out;
wire _guard557 = _guard555 & _guard556;
wire _guard558 = cond_wire42_out;
wire _guard559 = early_reset_static_par0_go_out;
wire _guard560 = _guard558 & _guard559;
wire _guard561 = cond_wire42_out;
wire _guard562 = early_reset_static_par0_go_out;
wire _guard563 = _guard561 & _guard562;
wire _guard564 = cond_wire53_out;
wire _guard565 = early_reset_static_par0_go_out;
wire _guard566 = _guard564 & _guard565;
wire _guard567 = cond_wire53_out;
wire _guard568 = early_reset_static_par0_go_out;
wire _guard569 = _guard567 & _guard568;
wire _guard570 = early_reset_static_par0_go_out;
wire _guard571 = early_reset_static_par0_go_out;
wire _guard572 = early_reset_static_par0_go_out;
wire _guard573 = early_reset_static_par0_go_out;
wire _guard574 = early_reset_static_par0_go_out;
wire _guard575 = early_reset_static_par0_go_out;
wire _guard576 = early_reset_static_par0_go_out;
wire _guard577 = early_reset_static_par0_go_out;
wire _guard578 = early_reset_static_par0_go_out;
wire _guard579 = early_reset_static_par0_go_out;
wire _guard580 = early_reset_static_par0_go_out;
wire _guard581 = early_reset_static_par0_go_out;
wire _guard582 = early_reset_static_par0_go_out;
wire _guard583 = ~_guard0;
wire _guard584 = early_reset_static_par0_go_out;
wire _guard585 = _guard583 & _guard584;
wire _guard586 = early_reset_static_par0_go_out;
wire _guard587 = early_reset_static_par0_go_out;
wire _guard588 = ~_guard0;
wire _guard589 = early_reset_static_par0_go_out;
wire _guard590 = _guard588 & _guard589;
wire _guard591 = early_reset_static_par0_go_out;
wire _guard592 = ~_guard0;
wire _guard593 = early_reset_static_par0_go_out;
wire _guard594 = _guard592 & _guard593;
wire _guard595 = early_reset_static_par0_go_out;
wire _guard596 = ~_guard0;
wire _guard597 = early_reset_static_par0_go_out;
wire _guard598 = _guard596 & _guard597;
wire _guard599 = early_reset_static_par0_go_out;
wire _guard600 = early_reset_static_par0_go_out;
wire _guard601 = early_reset_static_par0_go_out;
wire _guard602 = early_reset_static_par0_go_out;
wire _guard603 = early_reset_static_par0_go_out;
wire _guard604 = cond_wire22_out;
wire _guard605 = early_reset_static_par0_go_out;
wire _guard606 = _guard604 & _guard605;
wire _guard607 = cond_wire20_out;
wire _guard608 = early_reset_static_par0_go_out;
wire _guard609 = _guard607 & _guard608;
wire _guard610 = fsm_out == 1'd0;
wire _guard611 = cond_wire20_out;
wire _guard612 = _guard610 & _guard611;
wire _guard613 = fsm_out == 1'd0;
wire _guard614 = _guard612 & _guard613;
wire _guard615 = fsm_out == 1'd0;
wire _guard616 = cond_wire22_out;
wire _guard617 = _guard615 & _guard616;
wire _guard618 = fsm_out == 1'd0;
wire _guard619 = _guard617 & _guard618;
wire _guard620 = _guard614 | _guard619;
wire _guard621 = early_reset_static_par0_go_out;
wire _guard622 = _guard620 & _guard621;
wire _guard623 = fsm_out == 1'd0;
wire _guard624 = cond_wire20_out;
wire _guard625 = _guard623 & _guard624;
wire _guard626 = fsm_out == 1'd0;
wire _guard627 = _guard625 & _guard626;
wire _guard628 = fsm_out == 1'd0;
wire _guard629 = cond_wire22_out;
wire _guard630 = _guard628 & _guard629;
wire _guard631 = fsm_out == 1'd0;
wire _guard632 = _guard630 & _guard631;
wire _guard633 = _guard627 | _guard632;
wire _guard634 = early_reset_static_par0_go_out;
wire _guard635 = _guard633 & _guard634;
wire _guard636 = fsm_out == 1'd0;
wire _guard637 = cond_wire20_out;
wire _guard638 = _guard636 & _guard637;
wire _guard639 = fsm_out == 1'd0;
wire _guard640 = _guard638 & _guard639;
wire _guard641 = fsm_out == 1'd0;
wire _guard642 = cond_wire22_out;
wire _guard643 = _guard641 & _guard642;
wire _guard644 = fsm_out == 1'd0;
wire _guard645 = _guard643 & _guard644;
wire _guard646 = _guard640 | _guard645;
wire _guard647 = early_reset_static_par0_go_out;
wire _guard648 = _guard646 & _guard647;
wire _guard649 = cond_wire19_out;
wire _guard650 = early_reset_static_par0_go_out;
wire _guard651 = _guard649 & _guard650;
wire _guard652 = cond_wire19_out;
wire _guard653 = early_reset_static_par0_go_out;
wire _guard654 = _guard652 & _guard653;
wire _guard655 = cond_wire21_out;
wire _guard656 = early_reset_static_par0_go_out;
wire _guard657 = _guard655 & _guard656;
wire _guard658 = cond_wire21_out;
wire _guard659 = early_reset_static_par0_go_out;
wire _guard660 = _guard658 & _guard659;
wire _guard661 = cond_wire11_out;
wire _guard662 = early_reset_static_par0_go_out;
wire _guard663 = _guard661 & _guard662;
wire _guard664 = cond_wire11_out;
wire _guard665 = early_reset_static_par0_go_out;
wire _guard666 = _guard664 & _guard665;
wire _guard667 = cond_wire36_out;
wire _guard668 = early_reset_static_par0_go_out;
wire _guard669 = _guard667 & _guard668;
wire _guard670 = cond_wire36_out;
wire _guard671 = early_reset_static_par0_go_out;
wire _guard672 = _guard670 & _guard671;
wire _guard673 = cond_wire55_out;
wire _guard674 = early_reset_static_par0_go_out;
wire _guard675 = _guard673 & _guard674;
wire _guard676 = cond_wire55_out;
wire _guard677 = early_reset_static_par0_go_out;
wire _guard678 = _guard676 & _guard677;
wire _guard679 = cond_wire64_out;
wire _guard680 = early_reset_static_par0_go_out;
wire _guard681 = _guard679 & _guard680;
wire _guard682 = cond_wire62_out;
wire _guard683 = early_reset_static_par0_go_out;
wire _guard684 = _guard682 & _guard683;
wire _guard685 = fsm_out == 1'd0;
wire _guard686 = cond_wire62_out;
wire _guard687 = _guard685 & _guard686;
wire _guard688 = fsm_out == 1'd0;
wire _guard689 = _guard687 & _guard688;
wire _guard690 = fsm_out == 1'd0;
wire _guard691 = cond_wire64_out;
wire _guard692 = _guard690 & _guard691;
wire _guard693 = fsm_out == 1'd0;
wire _guard694 = _guard692 & _guard693;
wire _guard695 = _guard689 | _guard694;
wire _guard696 = early_reset_static_par0_go_out;
wire _guard697 = _guard695 & _guard696;
wire _guard698 = fsm_out == 1'd0;
wire _guard699 = cond_wire62_out;
wire _guard700 = _guard698 & _guard699;
wire _guard701 = fsm_out == 1'd0;
wire _guard702 = _guard700 & _guard701;
wire _guard703 = fsm_out == 1'd0;
wire _guard704 = cond_wire64_out;
wire _guard705 = _guard703 & _guard704;
wire _guard706 = fsm_out == 1'd0;
wire _guard707 = _guard705 & _guard706;
wire _guard708 = _guard702 | _guard707;
wire _guard709 = early_reset_static_par0_go_out;
wire _guard710 = _guard708 & _guard709;
wire _guard711 = fsm_out == 1'd0;
wire _guard712 = cond_wire62_out;
wire _guard713 = _guard711 & _guard712;
wire _guard714 = fsm_out == 1'd0;
wire _guard715 = _guard713 & _guard714;
wire _guard716 = fsm_out == 1'd0;
wire _guard717 = cond_wire64_out;
wire _guard718 = _guard716 & _guard717;
wire _guard719 = fsm_out == 1'd0;
wire _guard720 = _guard718 & _guard719;
wire _guard721 = _guard715 | _guard720;
wire _guard722 = early_reset_static_par0_go_out;
wire _guard723 = _guard721 & _guard722;
wire _guard724 = early_reset_static_par_go_out;
wire _guard725 = cond_wire4_out;
wire _guard726 = early_reset_static_par0_go_out;
wire _guard727 = _guard725 & _guard726;
wire _guard728 = _guard724 | _guard727;
wire _guard729 = cond_wire4_out;
wire _guard730 = early_reset_static_par0_go_out;
wire _guard731 = _guard729 & _guard730;
wire _guard732 = early_reset_static_par_go_out;
wire _guard733 = early_reset_static_par0_go_out;
wire _guard734 = early_reset_static_par0_go_out;
wire _guard735 = early_reset_static_par0_go_out;
wire _guard736 = early_reset_static_par0_go_out;
wire _guard737 = early_reset_static_par_go_out;
wire _guard738 = early_reset_static_par0_go_out;
wire _guard739 = _guard737 | _guard738;
wire _guard740 = early_reset_static_par_go_out;
wire _guard741 = early_reset_static_par0_go_out;
wire _guard742 = early_reset_static_par0_go_out;
wire _guard743 = early_reset_static_par0_go_out;
wire _guard744 = early_reset_static_par0_go_out;
wire _guard745 = early_reset_static_par0_go_out;
wire _guard746 = early_reset_static_par0_go_out;
wire _guard747 = early_reset_static_par0_go_out;
wire _guard748 = early_reset_static_par0_go_out;
wire _guard749 = ~_guard0;
wire _guard750 = early_reset_static_par0_go_out;
wire _guard751 = _guard749 & _guard750;
wire _guard752 = early_reset_static_par0_go_out;
wire _guard753 = ~_guard0;
wire _guard754 = early_reset_static_par0_go_out;
wire _guard755 = _guard753 & _guard754;
wire _guard756 = ~_guard0;
wire _guard757 = early_reset_static_par0_go_out;
wire _guard758 = _guard756 & _guard757;
wire _guard759 = early_reset_static_par0_go_out;
wire _guard760 = early_reset_static_par0_go_out;
wire _guard761 = ~_guard0;
wire _guard762 = early_reset_static_par0_go_out;
wire _guard763 = _guard761 & _guard762;
wire _guard764 = early_reset_static_par0_go_out;
wire _guard765 = early_reset_static_par0_go_out;
wire _guard766 = early_reset_static_par0_go_out;
wire _guard767 = early_reset_static_par0_go_out;
wire _guard768 = early_reset_static_par0_go_out;
wire _guard769 = early_reset_static_par0_go_out;
wire _guard770 = cond_wire_out;
wire _guard771 = early_reset_static_par0_go_out;
wire _guard772 = _guard770 & _guard771;
wire _guard773 = cond_wire_out;
wire _guard774 = early_reset_static_par0_go_out;
wire _guard775 = _guard773 & _guard774;
wire _guard776 = cond_wire17_out;
wire _guard777 = early_reset_static_par0_go_out;
wire _guard778 = _guard776 & _guard777;
wire _guard779 = cond_wire15_out;
wire _guard780 = early_reset_static_par0_go_out;
wire _guard781 = _guard779 & _guard780;
wire _guard782 = fsm_out == 1'd0;
wire _guard783 = cond_wire15_out;
wire _guard784 = _guard782 & _guard783;
wire _guard785 = fsm_out == 1'd0;
wire _guard786 = _guard784 & _guard785;
wire _guard787 = fsm_out == 1'd0;
wire _guard788 = cond_wire17_out;
wire _guard789 = _guard787 & _guard788;
wire _guard790 = fsm_out == 1'd0;
wire _guard791 = _guard789 & _guard790;
wire _guard792 = _guard786 | _guard791;
wire _guard793 = early_reset_static_par0_go_out;
wire _guard794 = _guard792 & _guard793;
wire _guard795 = fsm_out == 1'd0;
wire _guard796 = cond_wire15_out;
wire _guard797 = _guard795 & _guard796;
wire _guard798 = fsm_out == 1'd0;
wire _guard799 = _guard797 & _guard798;
wire _guard800 = fsm_out == 1'd0;
wire _guard801 = cond_wire17_out;
wire _guard802 = _guard800 & _guard801;
wire _guard803 = fsm_out == 1'd0;
wire _guard804 = _guard802 & _guard803;
wire _guard805 = _guard799 | _guard804;
wire _guard806 = early_reset_static_par0_go_out;
wire _guard807 = _guard805 & _guard806;
wire _guard808 = fsm_out == 1'd0;
wire _guard809 = cond_wire15_out;
wire _guard810 = _guard808 & _guard809;
wire _guard811 = fsm_out == 1'd0;
wire _guard812 = _guard810 & _guard811;
wire _guard813 = fsm_out == 1'd0;
wire _guard814 = cond_wire17_out;
wire _guard815 = _guard813 & _guard814;
wire _guard816 = fsm_out == 1'd0;
wire _guard817 = _guard815 & _guard816;
wire _guard818 = _guard812 | _guard817;
wire _guard819 = early_reset_static_par0_go_out;
wire _guard820 = _guard818 & _guard819;
wire _guard821 = cond_wire16_out;
wire _guard822 = early_reset_static_par0_go_out;
wire _guard823 = _guard821 & _guard822;
wire _guard824 = cond_wire16_out;
wire _guard825 = early_reset_static_par0_go_out;
wire _guard826 = _guard824 & _guard825;
wire _guard827 = cond_wire46_out;
wire _guard828 = early_reset_static_par0_go_out;
wire _guard829 = _guard827 & _guard828;
wire _guard830 = cond_wire46_out;
wire _guard831 = early_reset_static_par0_go_out;
wire _guard832 = _guard830 & _guard831;
wire _guard833 = cond_wire56_out;
wire _guard834 = early_reset_static_par0_go_out;
wire _guard835 = _guard833 & _guard834;
wire _guard836 = cond_wire54_out;
wire _guard837 = early_reset_static_par0_go_out;
wire _guard838 = _guard836 & _guard837;
wire _guard839 = fsm_out == 1'd0;
wire _guard840 = cond_wire54_out;
wire _guard841 = _guard839 & _guard840;
wire _guard842 = fsm_out == 1'd0;
wire _guard843 = _guard841 & _guard842;
wire _guard844 = fsm_out == 1'd0;
wire _guard845 = cond_wire56_out;
wire _guard846 = _guard844 & _guard845;
wire _guard847 = fsm_out == 1'd0;
wire _guard848 = _guard846 & _guard847;
wire _guard849 = _guard843 | _guard848;
wire _guard850 = early_reset_static_par0_go_out;
wire _guard851 = _guard849 & _guard850;
wire _guard852 = fsm_out == 1'd0;
wire _guard853 = cond_wire54_out;
wire _guard854 = _guard852 & _guard853;
wire _guard855 = fsm_out == 1'd0;
wire _guard856 = _guard854 & _guard855;
wire _guard857 = fsm_out == 1'd0;
wire _guard858 = cond_wire56_out;
wire _guard859 = _guard857 & _guard858;
wire _guard860 = fsm_out == 1'd0;
wire _guard861 = _guard859 & _guard860;
wire _guard862 = _guard856 | _guard861;
wire _guard863 = early_reset_static_par0_go_out;
wire _guard864 = _guard862 & _guard863;
wire _guard865 = fsm_out == 1'd0;
wire _guard866 = cond_wire54_out;
wire _guard867 = _guard865 & _guard866;
wire _guard868 = fsm_out == 1'd0;
wire _guard869 = _guard867 & _guard868;
wire _guard870 = fsm_out == 1'd0;
wire _guard871 = cond_wire56_out;
wire _guard872 = _guard870 & _guard871;
wire _guard873 = fsm_out == 1'd0;
wire _guard874 = _guard872 & _guard873;
wire _guard875 = _guard869 | _guard874;
wire _guard876 = early_reset_static_par0_go_out;
wire _guard877 = _guard875 & _guard876;
wire _guard878 = cond_wire46_out;
wire _guard879 = early_reset_static_par0_go_out;
wire _guard880 = _guard878 & _guard879;
wire _guard881 = cond_wire46_out;
wire _guard882 = early_reset_static_par0_go_out;
wire _guard883 = _guard881 & _guard882;
wire _guard884 = early_reset_static_par_go_out;
wire _guard885 = early_reset_static_par0_go_out;
wire _guard886 = _guard884 | _guard885;
wire _guard887 = early_reset_static_par0_go_out;
wire _guard888 = early_reset_static_par_go_out;
wire _guard889 = early_reset_static_par_go_out;
wire _guard890 = early_reset_static_par0_go_out;
wire _guard891 = _guard889 | _guard890;
wire _guard892 = early_reset_static_par_go_out;
wire _guard893 = early_reset_static_par0_go_out;
wire _guard894 = early_reset_static_par0_go_out;
wire _guard895 = early_reset_static_par0_go_out;
wire _guard896 = early_reset_static_par0_go_out;
wire _guard897 = early_reset_static_par0_go_out;
wire _guard898 = early_reset_static_par0_go_out;
wire _guard899 = ~_guard0;
wire _guard900 = early_reset_static_par0_go_out;
wire _guard901 = _guard899 & _guard900;
wire _guard902 = early_reset_static_par0_go_out;
wire _guard903 = early_reset_static_par0_go_out;
wire _guard904 = ~_guard0;
wire _guard905 = early_reset_static_par0_go_out;
wire _guard906 = _guard904 & _guard905;
wire _guard907 = early_reset_static_par0_go_out;
wire _guard908 = early_reset_static_par0_go_out;
wire _guard909 = early_reset_static_par0_go_out;
wire _guard910 = early_reset_static_par0_go_out;
wire _guard911 = early_reset_static_par0_go_out;
wire _guard912 = early_reset_static_par0_go_out;
wire _guard913 = early_reset_static_par0_go_out;
wire _guard914 = early_reset_static_par0_go_out;
wire _guard915 = ~_guard0;
wire _guard916 = early_reset_static_par0_go_out;
wire _guard917 = _guard915 & _guard916;
wire _guard918 = early_reset_static_par0_go_out;
wire _guard919 = ~_guard0;
wire _guard920 = early_reset_static_par0_go_out;
wire _guard921 = _guard919 & _guard920;
wire _guard922 = wrapper_early_reset_static_par_done_out;
wire _guard923 = ~_guard922;
wire _guard924 = fsm0_out == 2'd0;
wire _guard925 = _guard923 & _guard924;
wire _guard926 = tdcc_go_out;
wire _guard927 = _guard925 & _guard926;
wire _guard928 = early_reset_static_par0_go_out;
wire _guard929 = early_reset_static_par0_go_out;
wire _guard930 = cond_wire12_out;
wire _guard931 = early_reset_static_par0_go_out;
wire _guard932 = _guard930 & _guard931;
wire _guard933 = cond_wire10_out;
wire _guard934 = early_reset_static_par0_go_out;
wire _guard935 = _guard933 & _guard934;
wire _guard936 = fsm_out == 1'd0;
wire _guard937 = cond_wire10_out;
wire _guard938 = _guard936 & _guard937;
wire _guard939 = fsm_out == 1'd0;
wire _guard940 = _guard938 & _guard939;
wire _guard941 = fsm_out == 1'd0;
wire _guard942 = cond_wire12_out;
wire _guard943 = _guard941 & _guard942;
wire _guard944 = fsm_out == 1'd0;
wire _guard945 = _guard943 & _guard944;
wire _guard946 = _guard940 | _guard945;
wire _guard947 = early_reset_static_par0_go_out;
wire _guard948 = _guard946 & _guard947;
wire _guard949 = fsm_out == 1'd0;
wire _guard950 = cond_wire10_out;
wire _guard951 = _guard949 & _guard950;
wire _guard952 = fsm_out == 1'd0;
wire _guard953 = _guard951 & _guard952;
wire _guard954 = fsm_out == 1'd0;
wire _guard955 = cond_wire12_out;
wire _guard956 = _guard954 & _guard955;
wire _guard957 = fsm_out == 1'd0;
wire _guard958 = _guard956 & _guard957;
wire _guard959 = _guard953 | _guard958;
wire _guard960 = early_reset_static_par0_go_out;
wire _guard961 = _guard959 & _guard960;
wire _guard962 = fsm_out == 1'd0;
wire _guard963 = cond_wire10_out;
wire _guard964 = _guard962 & _guard963;
wire _guard965 = fsm_out == 1'd0;
wire _guard966 = _guard964 & _guard965;
wire _guard967 = fsm_out == 1'd0;
wire _guard968 = cond_wire12_out;
wire _guard969 = _guard967 & _guard968;
wire _guard970 = fsm_out == 1'd0;
wire _guard971 = _guard969 & _guard970;
wire _guard972 = _guard966 | _guard971;
wire _guard973 = early_reset_static_par0_go_out;
wire _guard974 = _guard972 & _guard973;
wire _guard975 = early_reset_static_par_go_out;
wire _guard976 = cond_wire_out;
wire _guard977 = early_reset_static_par0_go_out;
wire _guard978 = _guard976 & _guard977;
wire _guard979 = _guard975 | _guard978;
wire _guard980 = cond_wire_out;
wire _guard981 = early_reset_static_par0_go_out;
wire _guard982 = _guard980 & _guard981;
wire _guard983 = early_reset_static_par_go_out;
wire _guard984 = early_reset_static_par_go_out;
wire _guard985 = cond_wire19_out;
wire _guard986 = early_reset_static_par0_go_out;
wire _guard987 = _guard985 & _guard986;
wire _guard988 = _guard984 | _guard987;
wire _guard989 = cond_wire19_out;
wire _guard990 = early_reset_static_par0_go_out;
wire _guard991 = _guard989 & _guard990;
wire _guard992 = early_reset_static_par_go_out;
wire _guard993 = early_reset_static_par0_go_out;
wire _guard994 = early_reset_static_par0_go_out;
wire _guard995 = early_reset_static_par0_go_out;
wire _guard996 = early_reset_static_par0_go_out;
wire _guard997 = early_reset_static_par0_go_out;
wire _guard998 = early_reset_static_par0_go_out;
wire _guard999 = early_reset_static_par_go_out;
wire _guard1000 = early_reset_static_par0_go_out;
wire _guard1001 = _guard999 | _guard1000;
wire _guard1002 = early_reset_static_par0_go_out;
wire _guard1003 = early_reset_static_par_go_out;
wire _guard1004 = early_reset_static_par0_go_out;
wire _guard1005 = early_reset_static_par0_go_out;
wire _guard1006 = early_reset_static_par0_go_out;
wire _guard1007 = early_reset_static_par0_go_out;
wire _guard1008 = early_reset_static_par0_go_out;
wire _guard1009 = early_reset_static_par0_go_out;
wire _guard1010 = early_reset_static_par0_go_out;
wire _guard1011 = early_reset_static_par0_go_out;
wire _guard1012 = early_reset_static_par0_go_out;
wire _guard1013 = early_reset_static_par0_go_out;
wire _guard1014 = early_reset_static_par0_go_out;
wire _guard1015 = early_reset_static_par0_go_out;
wire _guard1016 = early_reset_static_par0_go_out;
wire _guard1017 = early_reset_static_par0_go_out;
wire _guard1018 = early_reset_static_par0_go_out;
wire _guard1019 = early_reset_static_par0_go_out;
wire _guard1020 = fsm_out == 1'd0;
wire _guard1021 = signal_reg_out;
wire _guard1022 = _guard1020 & _guard1021;
wire _guard1023 = cond_wire43_out;
wire _guard1024 = early_reset_static_par0_go_out;
wire _guard1025 = _guard1023 & _guard1024;
wire _guard1026 = cond_wire41_out;
wire _guard1027 = early_reset_static_par0_go_out;
wire _guard1028 = _guard1026 & _guard1027;
wire _guard1029 = fsm_out == 1'd0;
wire _guard1030 = cond_wire41_out;
wire _guard1031 = _guard1029 & _guard1030;
wire _guard1032 = fsm_out == 1'd0;
wire _guard1033 = _guard1031 & _guard1032;
wire _guard1034 = fsm_out == 1'd0;
wire _guard1035 = cond_wire43_out;
wire _guard1036 = _guard1034 & _guard1035;
wire _guard1037 = fsm_out == 1'd0;
wire _guard1038 = _guard1036 & _guard1037;
wire _guard1039 = _guard1033 | _guard1038;
wire _guard1040 = early_reset_static_par0_go_out;
wire _guard1041 = _guard1039 & _guard1040;
wire _guard1042 = fsm_out == 1'd0;
wire _guard1043 = cond_wire41_out;
wire _guard1044 = _guard1042 & _guard1043;
wire _guard1045 = fsm_out == 1'd0;
wire _guard1046 = _guard1044 & _guard1045;
wire _guard1047 = fsm_out == 1'd0;
wire _guard1048 = cond_wire43_out;
wire _guard1049 = _guard1047 & _guard1048;
wire _guard1050 = fsm_out == 1'd0;
wire _guard1051 = _guard1049 & _guard1050;
wire _guard1052 = _guard1046 | _guard1051;
wire _guard1053 = early_reset_static_par0_go_out;
wire _guard1054 = _guard1052 & _guard1053;
wire _guard1055 = fsm_out == 1'd0;
wire _guard1056 = cond_wire41_out;
wire _guard1057 = _guard1055 & _guard1056;
wire _guard1058 = fsm_out == 1'd0;
wire _guard1059 = _guard1057 & _guard1058;
wire _guard1060 = fsm_out == 1'd0;
wire _guard1061 = cond_wire43_out;
wire _guard1062 = _guard1060 & _guard1061;
wire _guard1063 = fsm_out == 1'd0;
wire _guard1064 = _guard1062 & _guard1063;
wire _guard1065 = _guard1059 | _guard1064;
wire _guard1066 = early_reset_static_par0_go_out;
wire _guard1067 = _guard1065 & _guard1066;
wire _guard1068 = cond_wire51_out;
wire _guard1069 = early_reset_static_par0_go_out;
wire _guard1070 = _guard1068 & _guard1069;
wire _guard1071 = cond_wire49_out;
wire _guard1072 = early_reset_static_par0_go_out;
wire _guard1073 = _guard1071 & _guard1072;
wire _guard1074 = fsm_out == 1'd0;
wire _guard1075 = cond_wire49_out;
wire _guard1076 = _guard1074 & _guard1075;
wire _guard1077 = fsm_out == 1'd0;
wire _guard1078 = _guard1076 & _guard1077;
wire _guard1079 = fsm_out == 1'd0;
wire _guard1080 = cond_wire51_out;
wire _guard1081 = _guard1079 & _guard1080;
wire _guard1082 = fsm_out == 1'd0;
wire _guard1083 = _guard1081 & _guard1082;
wire _guard1084 = _guard1078 | _guard1083;
wire _guard1085 = early_reset_static_par0_go_out;
wire _guard1086 = _guard1084 & _guard1085;
wire _guard1087 = fsm_out == 1'd0;
wire _guard1088 = cond_wire49_out;
wire _guard1089 = _guard1087 & _guard1088;
wire _guard1090 = fsm_out == 1'd0;
wire _guard1091 = _guard1089 & _guard1090;
wire _guard1092 = fsm_out == 1'd0;
wire _guard1093 = cond_wire51_out;
wire _guard1094 = _guard1092 & _guard1093;
wire _guard1095 = fsm_out == 1'd0;
wire _guard1096 = _guard1094 & _guard1095;
wire _guard1097 = _guard1091 | _guard1096;
wire _guard1098 = early_reset_static_par0_go_out;
wire _guard1099 = _guard1097 & _guard1098;
wire _guard1100 = fsm_out == 1'd0;
wire _guard1101 = cond_wire49_out;
wire _guard1102 = _guard1100 & _guard1101;
wire _guard1103 = fsm_out == 1'd0;
wire _guard1104 = _guard1102 & _guard1103;
wire _guard1105 = fsm_out == 1'd0;
wire _guard1106 = cond_wire51_out;
wire _guard1107 = _guard1105 & _guard1106;
wire _guard1108 = fsm_out == 1'd0;
wire _guard1109 = _guard1107 & _guard1108;
wire _guard1110 = _guard1104 | _guard1109;
wire _guard1111 = early_reset_static_par0_go_out;
wire _guard1112 = _guard1110 & _guard1111;
wire _guard1113 = cond_wire60_out;
wire _guard1114 = early_reset_static_par0_go_out;
wire _guard1115 = _guard1113 & _guard1114;
wire _guard1116 = cond_wire58_out;
wire _guard1117 = early_reset_static_par0_go_out;
wire _guard1118 = _guard1116 & _guard1117;
wire _guard1119 = fsm_out == 1'd0;
wire _guard1120 = cond_wire58_out;
wire _guard1121 = _guard1119 & _guard1120;
wire _guard1122 = fsm_out == 1'd0;
wire _guard1123 = _guard1121 & _guard1122;
wire _guard1124 = fsm_out == 1'd0;
wire _guard1125 = cond_wire60_out;
wire _guard1126 = _guard1124 & _guard1125;
wire _guard1127 = fsm_out == 1'd0;
wire _guard1128 = _guard1126 & _guard1127;
wire _guard1129 = _guard1123 | _guard1128;
wire _guard1130 = early_reset_static_par0_go_out;
wire _guard1131 = _guard1129 & _guard1130;
wire _guard1132 = fsm_out == 1'd0;
wire _guard1133 = cond_wire58_out;
wire _guard1134 = _guard1132 & _guard1133;
wire _guard1135 = fsm_out == 1'd0;
wire _guard1136 = _guard1134 & _guard1135;
wire _guard1137 = fsm_out == 1'd0;
wire _guard1138 = cond_wire60_out;
wire _guard1139 = _guard1137 & _guard1138;
wire _guard1140 = fsm_out == 1'd0;
wire _guard1141 = _guard1139 & _guard1140;
wire _guard1142 = _guard1136 | _guard1141;
wire _guard1143 = early_reset_static_par0_go_out;
wire _guard1144 = _guard1142 & _guard1143;
wire _guard1145 = fsm_out == 1'd0;
wire _guard1146 = cond_wire58_out;
wire _guard1147 = _guard1145 & _guard1146;
wire _guard1148 = fsm_out == 1'd0;
wire _guard1149 = _guard1147 & _guard1148;
wire _guard1150 = fsm_out == 1'd0;
wire _guard1151 = cond_wire60_out;
wire _guard1152 = _guard1150 & _guard1151;
wire _guard1153 = fsm_out == 1'd0;
wire _guard1154 = _guard1152 & _guard1153;
wire _guard1155 = _guard1149 | _guard1154;
wire _guard1156 = early_reset_static_par0_go_out;
wire _guard1157 = _guard1155 & _guard1156;
wire _guard1158 = early_reset_static_par_go_out;
wire _guard1159 = early_reset_static_par0_go_out;
wire _guard1160 = early_reset_static_par_go_out;
wire _guard1161 = early_reset_static_par0_go_out;
wire _guard1162 = early_reset_static_par0_go_out;
wire _guard1163 = early_reset_static_par0_go_out;
wire _guard1164 = early_reset_static_par0_go_out;
wire _guard1165 = early_reset_static_par0_go_out;
wire _guard1166 = early_reset_static_par0_go_out;
wire _guard1167 = early_reset_static_par0_go_out;
wire _guard1168 = early_reset_static_par0_go_out;
wire _guard1169 = early_reset_static_par0_go_out;
wire _guard1170 = early_reset_static_par0_go_out;
wire _guard1171 = ~_guard0;
wire _guard1172 = early_reset_static_par0_go_out;
wire _guard1173 = _guard1171 & _guard1172;
wire _guard1174 = early_reset_static_par0_go_out;
wire _guard1175 = early_reset_static_par0_go_out;
wire _guard1176 = early_reset_static_par0_go_out;
wire _guard1177 = early_reset_static_par0_go_out;
wire _guard1178 = ~_guard0;
wire _guard1179 = early_reset_static_par0_go_out;
wire _guard1180 = _guard1178 & _guard1179;
wire _guard1181 = early_reset_static_par0_go_out;
wire _guard1182 = early_reset_static_par0_go_out;
wire _guard1183 = early_reset_static_par0_go_out;
wire _guard1184 = early_reset_static_par0_go_out;
wire _guard1185 = early_reset_static_par0_go_out;
wire _guard1186 = early_reset_static_par0_go_out;
wire _guard1187 = early_reset_static_par0_go_out;
wire _guard1188 = fsm0_out == 2'd2;
wire _guard1189 = fsm0_out == 2'd0;
wire _guard1190 = wrapper_early_reset_static_par_done_out;
wire _guard1191 = _guard1189 & _guard1190;
wire _guard1192 = tdcc_go_out;
wire _guard1193 = _guard1191 & _guard1192;
wire _guard1194 = _guard1188 | _guard1193;
wire _guard1195 = fsm0_out == 2'd1;
wire _guard1196 = while_wrapper_early_reset_static_par0_done_out;
wire _guard1197 = _guard1195 & _guard1196;
wire _guard1198 = tdcc_go_out;
wire _guard1199 = _guard1197 & _guard1198;
wire _guard1200 = _guard1194 | _guard1199;
wire _guard1201 = fsm0_out == 2'd0;
wire _guard1202 = wrapper_early_reset_static_par_done_out;
wire _guard1203 = _guard1201 & _guard1202;
wire _guard1204 = tdcc_go_out;
wire _guard1205 = _guard1203 & _guard1204;
wire _guard1206 = fsm0_out == 2'd2;
wire _guard1207 = fsm0_out == 2'd1;
wire _guard1208 = while_wrapper_early_reset_static_par0_done_out;
wire _guard1209 = _guard1207 & _guard1208;
wire _guard1210 = tdcc_go_out;
wire _guard1211 = _guard1209 & _guard1210;
wire _guard1212 = early_reset_static_par0_go_out;
wire _guard1213 = early_reset_static_par_go_out;
wire _guard1214 = early_reset_static_par_go_out;
wire _guard1215 = early_reset_static_par0_go_out;
wire _guard1216 = early_reset_static_par0_go_out;
wire _guard1217 = early_reset_static_par0_go_out;
wire _guard1218 = early_reset_static_par0_go_out;
wire _guard1219 = early_reset_static_par0_go_out;
wire _guard1220 = cond_wire21_out;
wire _guard1221 = early_reset_static_par0_go_out;
wire _guard1222 = _guard1220 & _guard1221;
wire _guard1223 = cond_wire21_out;
wire _guard1224 = early_reset_static_par0_go_out;
wire _guard1225 = _guard1223 & _guard1224;
wire _guard1226 = cond_wire38_out;
wire _guard1227 = early_reset_static_par0_go_out;
wire _guard1228 = _guard1226 & _guard1227;
wire _guard1229 = cond_wire38_out;
wire _guard1230 = early_reset_static_par0_go_out;
wire _guard1231 = _guard1229 & _guard1230;
wire _guard1232 = cond_wire42_out;
wire _guard1233 = early_reset_static_par0_go_out;
wire _guard1234 = _guard1232 & _guard1233;
wire _guard1235 = cond_wire42_out;
wire _guard1236 = early_reset_static_par0_go_out;
wire _guard1237 = _guard1235 & _guard1236;
wire _guard1238 = early_reset_static_par_go_out;
wire _guard1239 = early_reset_static_par0_go_out;
wire _guard1240 = _guard1238 | _guard1239;
wire _guard1241 = early_reset_static_par_go_out;
wire _guard1242 = early_reset_static_par0_go_out;
wire _guard1243 = early_reset_static_par_go_out;
wire _guard1244 = early_reset_static_par0_go_out;
wire _guard1245 = _guard1243 | _guard1244;
wire _guard1246 = early_reset_static_par0_go_out;
wire _guard1247 = early_reset_static_par_go_out;
wire _guard1248 = early_reset_static_par0_go_out;
wire _guard1249 = early_reset_static_par0_go_out;
wire _guard1250 = early_reset_static_par_go_out;
wire _guard1251 = early_reset_static_par0_go_out;
wire _guard1252 = _guard1250 | _guard1251;
wire _guard1253 = early_reset_static_par_go_out;
wire _guard1254 = early_reset_static_par0_go_out;
wire _guard1255 = early_reset_static_par0_go_out;
wire _guard1256 = early_reset_static_par0_go_out;
wire _guard1257 = early_reset_static_par0_go_out;
wire _guard1258 = early_reset_static_par0_go_out;
wire _guard1259 = early_reset_static_par0_go_out;
wire _guard1260 = early_reset_static_par0_go_out;
wire _guard1261 = early_reset_static_par_go_out;
wire _guard1262 = early_reset_static_par0_go_out;
wire _guard1263 = _guard1261 | _guard1262;
wire _guard1264 = early_reset_static_par_go_out;
wire _guard1265 = early_reset_static_par0_go_out;
wire _guard1266 = early_reset_static_par0_go_out;
wire _guard1267 = early_reset_static_par0_go_out;
wire _guard1268 = early_reset_static_par0_go_out;
wire _guard1269 = early_reset_static_par0_go_out;
wire _guard1270 = early_reset_static_par0_go_out;
wire _guard1271 = early_reset_static_par0_go_out;
wire _guard1272 = early_reset_static_par0_go_out;
wire _guard1273 = early_reset_static_par0_go_out;
wire _guard1274 = early_reset_static_par0_go_out;
wire _guard1275 = ~_guard0;
wire _guard1276 = early_reset_static_par0_go_out;
wire _guard1277 = _guard1275 & _guard1276;
wire _guard1278 = early_reset_static_par0_go_out;
wire _guard1279 = early_reset_static_par0_go_out;
wire _guard1280 = early_reset_static_par0_go_out;
wire _guard1281 = early_reset_static_par0_go_out;
wire _guard1282 = ~_guard0;
wire _guard1283 = early_reset_static_par0_go_out;
wire _guard1284 = _guard1282 & _guard1283;
wire _guard1285 = early_reset_static_par0_go_out;
wire _guard1286 = early_reset_static_par0_go_out;
wire _guard1287 = early_reset_static_par0_go_out;
wire _guard1288 = early_reset_static_par0_go_out;
wire _guard1289 = early_reset_static_par0_go_out;
wire _guard1290 = early_reset_static_par0_go_out;
wire _guard1291 = ~_guard0;
wire _guard1292 = early_reset_static_par0_go_out;
wire _guard1293 = _guard1291 & _guard1292;
wire _guard1294 = early_reset_static_par0_go_out;
wire _guard1295 = early_reset_static_par0_go_out;
wire _guard1296 = ~_guard0;
wire _guard1297 = early_reset_static_par0_go_out;
wire _guard1298 = _guard1296 & _guard1297;
wire _guard1299 = early_reset_static_par0_go_out;
wire _guard1300 = ~_guard0;
wire _guard1301 = early_reset_static_par0_go_out;
wire _guard1302 = _guard1300 & _guard1301;
wire _guard1303 = early_reset_static_par0_go_out;
wire _guard1304 = early_reset_static_par_go_out;
wire _guard1305 = lt_iter_limit_out;
wire _guard1306 = early_reset_static_par_go_out;
wire _guard1307 = _guard1305 & _guard1306;
wire _guard1308 = lt_iter_limit_out;
wire _guard1309 = ~_guard1308;
wire _guard1310 = early_reset_static_par_go_out;
wire _guard1311 = _guard1309 & _guard1310;
wire _guard1312 = early_reset_static_par0_go_out;
wire _guard1313 = early_reset_static_par0_go_out;
wire _guard1314 = cond_wire4_out;
wire _guard1315 = early_reset_static_par0_go_out;
wire _guard1316 = _guard1314 & _guard1315;
wire _guard1317 = cond_wire4_out;
wire _guard1318 = early_reset_static_par0_go_out;
wire _guard1319 = _guard1317 & _guard1318;
wire _guard1320 = cond_wire6_out;
wire _guard1321 = early_reset_static_par0_go_out;
wire _guard1322 = _guard1320 & _guard1321;
wire _guard1323 = cond_wire6_out;
wire _guard1324 = early_reset_static_par0_go_out;
wire _guard1325 = _guard1323 & _guard1324;
wire _guard1326 = cond_wire33_out;
wire _guard1327 = early_reset_static_par0_go_out;
wire _guard1328 = _guard1326 & _guard1327;
wire _guard1329 = cond_wire33_out;
wire _guard1330 = early_reset_static_par0_go_out;
wire _guard1331 = _guard1329 & _guard1330;
wire _guard1332 = cond_wire53_out;
wire _guard1333 = early_reset_static_par0_go_out;
wire _guard1334 = _guard1332 & _guard1333;
wire _guard1335 = cond_wire53_out;
wire _guard1336 = early_reset_static_par0_go_out;
wire _guard1337 = _guard1335 & _guard1336;
wire _guard1338 = early_reset_static_par_go_out;
wire _guard1339 = early_reset_static_par0_go_out;
wire _guard1340 = _guard1338 | _guard1339;
wire _guard1341 = early_reset_static_par0_go_out;
wire _guard1342 = early_reset_static_par_go_out;
wire _guard1343 = early_reset_static_par0_go_out;
wire _guard1344 = early_reset_static_par0_go_out;
wire _guard1345 = early_reset_static_par_go_out;
wire _guard1346 = early_reset_static_par0_go_out;
wire _guard1347 = _guard1345 | _guard1346;
wire _guard1348 = early_reset_static_par_go_out;
wire _guard1349 = early_reset_static_par0_go_out;
wire _guard1350 = early_reset_static_par0_go_out;
wire _guard1351 = early_reset_static_par0_go_out;
wire _guard1352 = early_reset_static_par0_go_out;
wire _guard1353 = early_reset_static_par0_go_out;
wire _guard1354 = early_reset_static_par0_go_out;
wire _guard1355 = early_reset_static_par0_go_out;
wire _guard1356 = ~_guard0;
wire _guard1357 = early_reset_static_par0_go_out;
wire _guard1358 = _guard1356 & _guard1357;
wire _guard1359 = early_reset_static_par0_go_out;
wire _guard1360 = early_reset_static_par0_go_out;
wire _guard1361 = early_reset_static_par0_go_out;
wire _guard1362 = ~_guard0;
wire _guard1363 = early_reset_static_par0_go_out;
wire _guard1364 = _guard1362 & _guard1363;
wire _guard1365 = early_reset_static_par0_go_out;
wire _guard1366 = early_reset_static_par0_go_out;
wire _guard1367 = early_reset_static_par0_go_out;
wire _guard1368 = ~_guard0;
wire _guard1369 = early_reset_static_par0_go_out;
wire _guard1370 = _guard1368 & _guard1369;
wire _guard1371 = early_reset_static_par0_go_out;
wire _guard1372 = early_reset_static_par0_go_out;
wire _guard1373 = early_reset_static_par0_go_out;
wire _guard1374 = early_reset_static_par0_go_out;
wire _guard1375 = ~_guard0;
wire _guard1376 = early_reset_static_par0_go_out;
wire _guard1377 = _guard1375 & _guard1376;
wire _guard1378 = early_reset_static_par0_go_out;
wire _guard1379 = early_reset_static_par0_go_out;
wire _guard1380 = early_reset_static_par0_go_out;
wire _guard1381 = early_reset_static_par0_go_out;
wire _guard1382 = cond_wire9_out;
wire _guard1383 = early_reset_static_par0_go_out;
wire _guard1384 = _guard1382 & _guard1383;
wire _guard1385 = cond_wire9_out;
wire _guard1386 = early_reset_static_par0_go_out;
wire _guard1387 = _guard1385 & _guard1386;
wire _guard1388 = cond_wire6_out;
wire _guard1389 = early_reset_static_par0_go_out;
wire _guard1390 = _guard1388 & _guard1389;
wire _guard1391 = cond_wire6_out;
wire _guard1392 = early_reset_static_par0_go_out;
wire _guard1393 = _guard1391 & _guard1392;
wire _guard1394 = cond_wire59_out;
wire _guard1395 = early_reset_static_par0_go_out;
wire _guard1396 = _guard1394 & _guard1395;
wire _guard1397 = cond_wire59_out;
wire _guard1398 = early_reset_static_par0_go_out;
wire _guard1399 = _guard1397 & _guard1398;
wire _guard1400 = cond_wire_out;
wire _guard1401 = early_reset_static_par0_go_out;
wire _guard1402 = _guard1400 & _guard1401;
wire _guard1403 = cond_wire_out;
wire _guard1404 = early_reset_static_par0_go_out;
wire _guard1405 = _guard1403 & _guard1404;
wire _guard1406 = cond_wire_out;
wire _guard1407 = early_reset_static_par0_go_out;
wire _guard1408 = _guard1406 & _guard1407;
wire _guard1409 = cond_wire_out;
wire _guard1410 = early_reset_static_par0_go_out;
wire _guard1411 = _guard1409 & _guard1410;
wire _guard1412 = early_reset_static_par0_go_out;
wire _guard1413 = early_reset_static_par0_go_out;
wire _guard1414 = early_reset_static_par0_go_out;
wire _guard1415 = early_reset_static_par0_go_out;
wire _guard1416 = early_reset_static_par0_go_out;
wire _guard1417 = early_reset_static_par0_go_out;
wire _guard1418 = early_reset_static_par0_go_out;
wire _guard1419 = early_reset_static_par0_go_out;
wire _guard1420 = ~_guard0;
wire _guard1421 = early_reset_static_par0_go_out;
wire _guard1422 = _guard1420 & _guard1421;
wire _guard1423 = early_reset_static_par0_go_out;
wire _guard1424 = ~_guard0;
wire _guard1425 = early_reset_static_par0_go_out;
wire _guard1426 = _guard1424 & _guard1425;
wire _guard1427 = early_reset_static_par0_go_out;
wire _guard1428 = early_reset_static_par0_go_out;
wire _guard1429 = early_reset_static_par0_go_out;
wire _guard1430 = ~_guard0;
wire _guard1431 = early_reset_static_par0_go_out;
wire _guard1432 = _guard1430 & _guard1431;
wire _guard1433 = early_reset_static_par0_go_out;
wire _guard1434 = early_reset_static_par0_go_out;
wire _guard1435 = early_reset_static_par0_go_out;
wire _guard1436 = early_reset_static_par0_go_out;
wire _guard1437 = early_reset_static_par0_go_out;
wire _guard1438 = early_reset_static_par0_go_out;
wire _guard1439 = early_reset_static_par0_go_out;
wire _guard1440 = early_reset_static_par0_go_out;
wire _guard1441 = early_reset_static_par0_go_out;
wire _guard1442 = ~_guard0;
wire _guard1443 = early_reset_static_par0_go_out;
wire _guard1444 = _guard1442 & _guard1443;
wire _guard1445 = early_reset_static_par0_go_out;
wire _guard1446 = ~_guard0;
wire _guard1447 = early_reset_static_par0_go_out;
wire _guard1448 = _guard1446 & _guard1447;
wire _guard1449 = early_reset_static_par0_go_out;
wire _guard1450 = early_reset_static_par0_go_out;
wire _guard1451 = early_reset_static_par0_go_out;
wire _guard1452 = early_reset_static_par0_go_out;
wire _guard1453 = ~_guard0;
wire _guard1454 = early_reset_static_par0_go_out;
wire _guard1455 = _guard1453 & _guard1454;
wire _guard1456 = ~_guard0;
wire _guard1457 = early_reset_static_par0_go_out;
wire _guard1458 = _guard1456 & _guard1457;
wire _guard1459 = early_reset_static_par0_go_out;
wire _guard1460 = early_reset_static_par0_go_out;
wire _guard1461 = early_reset_static_par0_go_out;
wire _guard1462 = fsm_out == 1'd0;
wire _guard1463 = signal_reg_out;
wire _guard1464 = _guard1462 & _guard1463;
wire _guard1465 = fsm_out == 1'd0;
wire _guard1466 = signal_reg_out;
wire _guard1467 = ~_guard1466;
wire _guard1468 = _guard1465 & _guard1467;
wire _guard1469 = wrapper_early_reset_static_par_go_out;
wire _guard1470 = _guard1468 & _guard1469;
wire _guard1471 = _guard1464 | _guard1470;
wire _guard1472 = fsm_out == 1'd0;
wire _guard1473 = signal_reg_out;
wire _guard1474 = ~_guard1473;
wire _guard1475 = _guard1472 & _guard1474;
wire _guard1476 = wrapper_early_reset_static_par_go_out;
wire _guard1477 = _guard1475 & _guard1476;
wire _guard1478 = fsm_out == 1'd0;
wire _guard1479 = signal_reg_out;
wire _guard1480 = _guard1478 & _guard1479;
wire _guard1481 = early_reset_static_par0_go_out;
wire _guard1482 = early_reset_static_par0_go_out;
wire _guard1483 = early_reset_static_par0_go_out;
wire _guard1484 = early_reset_static_par0_go_out;
wire _guard1485 = cond_wire39_out;
wire _guard1486 = early_reset_static_par0_go_out;
wire _guard1487 = _guard1485 & _guard1486;
wire _guard1488 = cond_wire37_out;
wire _guard1489 = early_reset_static_par0_go_out;
wire _guard1490 = _guard1488 & _guard1489;
wire _guard1491 = fsm_out == 1'd0;
wire _guard1492 = cond_wire37_out;
wire _guard1493 = _guard1491 & _guard1492;
wire _guard1494 = fsm_out == 1'd0;
wire _guard1495 = _guard1493 & _guard1494;
wire _guard1496 = fsm_out == 1'd0;
wire _guard1497 = cond_wire39_out;
wire _guard1498 = _guard1496 & _guard1497;
wire _guard1499 = fsm_out == 1'd0;
wire _guard1500 = _guard1498 & _guard1499;
wire _guard1501 = _guard1495 | _guard1500;
wire _guard1502 = early_reset_static_par0_go_out;
wire _guard1503 = _guard1501 & _guard1502;
wire _guard1504 = fsm_out == 1'd0;
wire _guard1505 = cond_wire37_out;
wire _guard1506 = _guard1504 & _guard1505;
wire _guard1507 = fsm_out == 1'd0;
wire _guard1508 = _guard1506 & _guard1507;
wire _guard1509 = fsm_out == 1'd0;
wire _guard1510 = cond_wire39_out;
wire _guard1511 = _guard1509 & _guard1510;
wire _guard1512 = fsm_out == 1'd0;
wire _guard1513 = _guard1511 & _guard1512;
wire _guard1514 = _guard1508 | _guard1513;
wire _guard1515 = early_reset_static_par0_go_out;
wire _guard1516 = _guard1514 & _guard1515;
wire _guard1517 = fsm_out == 1'd0;
wire _guard1518 = cond_wire37_out;
wire _guard1519 = _guard1517 & _guard1518;
wire _guard1520 = fsm_out == 1'd0;
wire _guard1521 = _guard1519 & _guard1520;
wire _guard1522 = fsm_out == 1'd0;
wire _guard1523 = cond_wire39_out;
wire _guard1524 = _guard1522 & _guard1523;
wire _guard1525 = fsm_out == 1'd0;
wire _guard1526 = _guard1524 & _guard1525;
wire _guard1527 = _guard1521 | _guard1526;
wire _guard1528 = early_reset_static_par0_go_out;
wire _guard1529 = _guard1527 & _guard1528;
wire _guard1530 = cond_wire38_out;
wire _guard1531 = early_reset_static_par0_go_out;
wire _guard1532 = _guard1530 & _guard1531;
wire _guard1533 = cond_wire38_out;
wire _guard1534 = early_reset_static_par0_go_out;
wire _guard1535 = _guard1533 & _guard1534;
wire _guard1536 = cond_wire29_out;
wire _guard1537 = early_reset_static_par0_go_out;
wire _guard1538 = _guard1536 & _guard1537;
wire _guard1539 = cond_wire29_out;
wire _guard1540 = early_reset_static_par0_go_out;
wire _guard1541 = _guard1539 & _guard1540;
wire _guard1542 = cond_wire4_out;
wire _guard1543 = early_reset_static_par0_go_out;
wire _guard1544 = _guard1542 & _guard1543;
wire _guard1545 = cond_wire4_out;
wire _guard1546 = early_reset_static_par0_go_out;
wire _guard1547 = _guard1545 & _guard1546;
wire _guard1548 = early_reset_static_par_go_out;
wire _guard1549 = cond_wire14_out;
wire _guard1550 = early_reset_static_par0_go_out;
wire _guard1551 = _guard1549 & _guard1550;
wire _guard1552 = _guard1548 | _guard1551;
wire _guard1553 = cond_wire14_out;
wire _guard1554 = early_reset_static_par0_go_out;
wire _guard1555 = _guard1553 & _guard1554;
wire _guard1556 = early_reset_static_par_go_out;
wire _guard1557 = early_reset_static_par0_go_out;
wire _guard1558 = early_reset_static_par0_go_out;
wire _guard1559 = early_reset_static_par0_go_out;
wire _guard1560 = early_reset_static_par0_go_out;
wire _guard1561 = early_reset_static_par0_go_out;
wire _guard1562 = early_reset_static_par0_go_out;
wire _guard1563 = early_reset_static_par_go_out;
wire _guard1564 = early_reset_static_par0_go_out;
wire _guard1565 = _guard1563 | _guard1564;
wire _guard1566 = early_reset_static_par0_go_out;
wire _guard1567 = early_reset_static_par_go_out;
wire _guard1568 = early_reset_static_par0_go_out;
wire _guard1569 = early_reset_static_par0_go_out;
wire _guard1570 = early_reset_static_par0_go_out;
wire _guard1571 = early_reset_static_par0_go_out;
wire _guard1572 = early_reset_static_par_go_out;
wire _guard1573 = early_reset_static_par0_go_out;
wire _guard1574 = _guard1572 | _guard1573;
wire _guard1575 = early_reset_static_par_go_out;
wire _guard1576 = early_reset_static_par0_go_out;
wire _guard1577 = early_reset_static_par0_go_out;
wire _guard1578 = early_reset_static_par0_go_out;
wire _guard1579 = early_reset_static_par_go_out;
wire _guard1580 = early_reset_static_par0_go_out;
wire _guard1581 = _guard1579 | _guard1580;
wire _guard1582 = early_reset_static_par_go_out;
wire _guard1583 = early_reset_static_par0_go_out;
wire _guard1584 = ~_guard0;
wire _guard1585 = early_reset_static_par0_go_out;
wire _guard1586 = _guard1584 & _guard1585;
wire _guard1587 = early_reset_static_par0_go_out;
wire _guard1588 = ~_guard0;
wire _guard1589 = early_reset_static_par0_go_out;
wire _guard1590 = _guard1588 & _guard1589;
wire _guard1591 = early_reset_static_par0_go_out;
wire _guard1592 = early_reset_static_par0_go_out;
wire _guard1593 = early_reset_static_par0_go_out;
wire _guard1594 = early_reset_static_par0_go_out;
wire _guard1595 = early_reset_static_par0_go_out;
wire _guard1596 = early_reset_static_par0_go_out;
wire _guard1597 = ~_guard0;
wire _guard1598 = early_reset_static_par0_go_out;
wire _guard1599 = _guard1597 & _guard1598;
wire _guard1600 = early_reset_static_par0_go_out;
wire _guard1601 = ~_guard0;
wire _guard1602 = early_reset_static_par0_go_out;
wire _guard1603 = _guard1601 & _guard1602;
wire _guard1604 = early_reset_static_par0_go_out;
wire _guard1605 = early_reset_static_par0_go_out;
wire _guard1606 = cond_wire2_out;
wire _guard1607 = early_reset_static_par0_go_out;
wire _guard1608 = _guard1606 & _guard1607;
wire _guard1609 = cond_wire0_out;
wire _guard1610 = early_reset_static_par0_go_out;
wire _guard1611 = _guard1609 & _guard1610;
wire _guard1612 = fsm_out == 1'd0;
wire _guard1613 = cond_wire0_out;
wire _guard1614 = _guard1612 & _guard1613;
wire _guard1615 = fsm_out == 1'd0;
wire _guard1616 = _guard1614 & _guard1615;
wire _guard1617 = fsm_out == 1'd0;
wire _guard1618 = cond_wire2_out;
wire _guard1619 = _guard1617 & _guard1618;
wire _guard1620 = fsm_out == 1'd0;
wire _guard1621 = _guard1619 & _guard1620;
wire _guard1622 = _guard1616 | _guard1621;
wire _guard1623 = early_reset_static_par0_go_out;
wire _guard1624 = _guard1622 & _guard1623;
wire _guard1625 = fsm_out == 1'd0;
wire _guard1626 = cond_wire0_out;
wire _guard1627 = _guard1625 & _guard1626;
wire _guard1628 = fsm_out == 1'd0;
wire _guard1629 = _guard1627 & _guard1628;
wire _guard1630 = fsm_out == 1'd0;
wire _guard1631 = cond_wire2_out;
wire _guard1632 = _guard1630 & _guard1631;
wire _guard1633 = fsm_out == 1'd0;
wire _guard1634 = _guard1632 & _guard1633;
wire _guard1635 = _guard1629 | _guard1634;
wire _guard1636 = early_reset_static_par0_go_out;
wire _guard1637 = _guard1635 & _guard1636;
wire _guard1638 = fsm_out == 1'd0;
wire _guard1639 = cond_wire0_out;
wire _guard1640 = _guard1638 & _guard1639;
wire _guard1641 = fsm_out == 1'd0;
wire _guard1642 = _guard1640 & _guard1641;
wire _guard1643 = fsm_out == 1'd0;
wire _guard1644 = cond_wire2_out;
wire _guard1645 = _guard1643 & _guard1644;
wire _guard1646 = fsm_out == 1'd0;
wire _guard1647 = _guard1645 & _guard1646;
wire _guard1648 = _guard1642 | _guard1647;
wire _guard1649 = early_reset_static_par0_go_out;
wire _guard1650 = _guard1648 & _guard1649;
wire _guard1651 = cond_wire67_out;
wire _guard1652 = early_reset_static_par0_go_out;
wire _guard1653 = _guard1651 & _guard1652;
wire _guard1654 = cond_wire66_out;
wire _guard1655 = early_reset_static_par0_go_out;
wire _guard1656 = _guard1654 & _guard1655;
wire _guard1657 = fsm_out == 1'd0;
wire _guard1658 = cond_wire66_out;
wire _guard1659 = _guard1657 & _guard1658;
wire _guard1660 = fsm_out == 1'd0;
wire _guard1661 = _guard1659 & _guard1660;
wire _guard1662 = fsm_out == 1'd0;
wire _guard1663 = cond_wire67_out;
wire _guard1664 = _guard1662 & _guard1663;
wire _guard1665 = fsm_out == 1'd0;
wire _guard1666 = _guard1664 & _guard1665;
wire _guard1667 = _guard1661 | _guard1666;
wire _guard1668 = early_reset_static_par0_go_out;
wire _guard1669 = _guard1667 & _guard1668;
wire _guard1670 = fsm_out == 1'd0;
wire _guard1671 = cond_wire66_out;
wire _guard1672 = _guard1670 & _guard1671;
wire _guard1673 = fsm_out == 1'd0;
wire _guard1674 = _guard1672 & _guard1673;
wire _guard1675 = fsm_out == 1'd0;
wire _guard1676 = cond_wire67_out;
wire _guard1677 = _guard1675 & _guard1676;
wire _guard1678 = fsm_out == 1'd0;
wire _guard1679 = _guard1677 & _guard1678;
wire _guard1680 = _guard1674 | _guard1679;
wire _guard1681 = early_reset_static_par0_go_out;
wire _guard1682 = _guard1680 & _guard1681;
wire _guard1683 = fsm_out == 1'd0;
wire _guard1684 = cond_wire66_out;
wire _guard1685 = _guard1683 & _guard1684;
wire _guard1686 = fsm_out == 1'd0;
wire _guard1687 = _guard1685 & _guard1686;
wire _guard1688 = fsm_out == 1'd0;
wire _guard1689 = cond_wire67_out;
wire _guard1690 = _guard1688 & _guard1689;
wire _guard1691 = fsm_out == 1'd0;
wire _guard1692 = _guard1690 & _guard1691;
wire _guard1693 = _guard1687 | _guard1692;
wire _guard1694 = early_reset_static_par0_go_out;
wire _guard1695 = _guard1693 & _guard1694;
wire _guard1696 = cond_wire50_out;
wire _guard1697 = early_reset_static_par0_go_out;
wire _guard1698 = _guard1696 & _guard1697;
wire _guard1699 = cond_wire50_out;
wire _guard1700 = early_reset_static_par0_go_out;
wire _guard1701 = _guard1699 & _guard1700;
wire _guard1702 = cond_wire9_out;
wire _guard1703 = early_reset_static_par0_go_out;
wire _guard1704 = _guard1702 & _guard1703;
wire _guard1705 = cond_wire9_out;
wire _guard1706 = early_reset_static_par0_go_out;
wire _guard1707 = _guard1705 & _guard1706;
wire _guard1708 = early_reset_static_par_go_out;
wire _guard1709 = early_reset_static_par0_go_out;
wire _guard1710 = _guard1708 | _guard1709;
wire _guard1711 = early_reset_static_par0_go_out;
wire _guard1712 = early_reset_static_par_go_out;
wire _guard1713 = early_reset_static_par_go_out;
wire _guard1714 = early_reset_static_par0_go_out;
wire _guard1715 = _guard1713 | _guard1714;
wire _guard1716 = early_reset_static_par_go_out;
wire _guard1717 = early_reset_static_par0_go_out;
wire _guard1718 = early_reset_static_par0_go_out;
wire _guard1719 = early_reset_static_par0_go_out;
wire _guard1720 = early_reset_static_par_go_out;
wire _guard1721 = early_reset_static_par0_go_out;
wire _guard1722 = _guard1720 | _guard1721;
wire _guard1723 = early_reset_static_par_go_out;
wire _guard1724 = early_reset_static_par0_go_out;
wire _guard1725 = early_reset_static_par0_go_out;
wire _guard1726 = early_reset_static_par0_go_out;
wire _guard1727 = early_reset_static_par_go_out;
wire _guard1728 = early_reset_static_par0_go_out;
wire _guard1729 = _guard1727 | _guard1728;
wire _guard1730 = early_reset_static_par_go_out;
wire _guard1731 = early_reset_static_par0_go_out;
wire _guard1732 = early_reset_static_par0_go_out;
wire _guard1733 = early_reset_static_par0_go_out;
wire _guard1734 = early_reset_static_par0_go_out;
wire _guard1735 = early_reset_static_par0_go_out;
wire _guard1736 = early_reset_static_par_go_out;
wire _guard1737 = early_reset_static_par0_go_out;
wire _guard1738 = _guard1736 | _guard1737;
wire _guard1739 = early_reset_static_par0_go_out;
wire _guard1740 = early_reset_static_par_go_out;
wire _guard1741 = early_reset_static_par0_go_out;
wire _guard1742 = early_reset_static_par0_go_out;
wire _guard1743 = early_reset_static_par0_go_out;
wire _guard1744 = early_reset_static_par0_go_out;
wire _guard1745 = early_reset_static_par0_go_out;
wire _guard1746 = early_reset_static_par0_go_out;
wire _guard1747 = early_reset_static_par_go_out;
wire _guard1748 = early_reset_static_par0_go_out;
wire _guard1749 = _guard1747 | _guard1748;
wire _guard1750 = early_reset_static_par_go_out;
wire _guard1751 = early_reset_static_par0_go_out;
wire _guard1752 = early_reset_static_par0_go_out;
wire _guard1753 = early_reset_static_par0_go_out;
wire _guard1754 = early_reset_static_par0_go_out;
wire _guard1755 = early_reset_static_par0_go_out;
wire _guard1756 = early_reset_static_par0_go_out;
wire _guard1757 = early_reset_static_par0_go_out;
wire _guard1758 = ~_guard0;
wire _guard1759 = early_reset_static_par0_go_out;
wire _guard1760 = _guard1758 & _guard1759;
wire _guard1761 = early_reset_static_par0_go_out;
wire _guard1762 = early_reset_static_par0_go_out;
wire _guard1763 = ~_guard0;
wire _guard1764 = early_reset_static_par0_go_out;
wire _guard1765 = _guard1763 & _guard1764;
wire _guard1766 = early_reset_static_par0_go_out;
wire _guard1767 = ~_guard0;
wire _guard1768 = early_reset_static_par0_go_out;
wire _guard1769 = _guard1767 & _guard1768;
wire _guard1770 = ~_guard0;
wire _guard1771 = early_reset_static_par0_go_out;
wire _guard1772 = _guard1770 & _guard1771;
wire _guard1773 = early_reset_static_par0_go_out;
wire _guard1774 = ~_guard0;
wire _guard1775 = early_reset_static_par0_go_out;
wire _guard1776 = _guard1774 & _guard1775;
wire _guard1777 = early_reset_static_par0_go_out;
wire _guard1778 = early_reset_static_par0_go_out;
wire _guard1779 = ~_guard0;
wire _guard1780 = early_reset_static_par0_go_out;
wire _guard1781 = _guard1779 & _guard1780;
wire _guard1782 = ~_guard0;
wire _guard1783 = early_reset_static_par0_go_out;
wire _guard1784 = _guard1782 & _guard1783;
wire _guard1785 = early_reset_static_par0_go_out;
wire _guard1786 = early_reset_static_par0_go_out;
wire _guard1787 = early_reset_static_par0_go_out;
wire _guard1788 = early_reset_static_par0_go_out;
wire _guard1789 = ~_guard0;
wire _guard1790 = early_reset_static_par0_go_out;
wire _guard1791 = _guard1789 & _guard1790;
wire _guard1792 = early_reset_static_par0_go_out;
wire _guard1793 = early_reset_static_par0_go_out;
wire _guard1794 = early_reset_static_par0_go_out;
wire _guard1795 = early_reset_static_par0_go_out;
wire _guard1796 = early_reset_static_par0_go_out;
wire _guard1797 = early_reset_static_par0_go_out;
wire _guard1798 = fsm0_out == 2'd2;
wire _guard1799 = cond_wire14_out;
wire _guard1800 = early_reset_static_par0_go_out;
wire _guard1801 = _guard1799 & _guard1800;
wire _guard1802 = cond_wire14_out;
wire _guard1803 = early_reset_static_par0_go_out;
wire _guard1804 = _guard1802 & _guard1803;
wire _guard1805 = cond_wire25_out;
wire _guard1806 = early_reset_static_par0_go_out;
wire _guard1807 = _guard1805 & _guard1806;
wire _guard1808 = cond_wire25_out;
wire _guard1809 = early_reset_static_par0_go_out;
wire _guard1810 = _guard1808 & _guard1809;
wire _guard1811 = cond_wire63_out;
wire _guard1812 = early_reset_static_par0_go_out;
wire _guard1813 = _guard1811 & _guard1812;
wire _guard1814 = cond_wire63_out;
wire _guard1815 = early_reset_static_par0_go_out;
wire _guard1816 = _guard1814 & _guard1815;
wire _guard1817 = early_reset_static_par_go_out;
wire _guard1818 = cond_wire9_out;
wire _guard1819 = early_reset_static_par0_go_out;
wire _guard1820 = _guard1818 & _guard1819;
wire _guard1821 = _guard1817 | _guard1820;
wire _guard1822 = cond_wire9_out;
wire _guard1823 = early_reset_static_par0_go_out;
wire _guard1824 = _guard1822 & _guard1823;
wire _guard1825 = early_reset_static_par_go_out;
wire _guard1826 = early_reset_static_par_go_out;
wire _guard1827 = cond_wire36_out;
wire _guard1828 = early_reset_static_par0_go_out;
wire _guard1829 = _guard1827 & _guard1828;
wire _guard1830 = _guard1826 | _guard1829;
wire _guard1831 = early_reset_static_par_go_out;
wire _guard1832 = cond_wire36_out;
wire _guard1833 = early_reset_static_par0_go_out;
wire _guard1834 = _guard1832 & _guard1833;
wire _guard1835 = early_reset_static_par0_go_out;
wire _guard1836 = early_reset_static_par0_go_out;
wire _guard1837 = early_reset_static_par0_go_out;
wire _guard1838 = early_reset_static_par0_go_out;
wire _guard1839 = early_reset_static_par0_go_out;
wire _guard1840 = early_reset_static_par0_go_out;
wire _guard1841 = early_reset_static_par_go_out;
wire _guard1842 = early_reset_static_par0_go_out;
wire _guard1843 = _guard1841 | _guard1842;
wire _guard1844 = early_reset_static_par0_go_out;
wire _guard1845 = early_reset_static_par_go_out;
wire _guard1846 = early_reset_static_par0_go_out;
wire _guard1847 = early_reset_static_par0_go_out;
wire _guard1848 = early_reset_static_par0_go_out;
wire _guard1849 = early_reset_static_par0_go_out;
wire _guard1850 = ~_guard0;
wire _guard1851 = early_reset_static_par0_go_out;
wire _guard1852 = _guard1850 & _guard1851;
wire _guard1853 = early_reset_static_par0_go_out;
wire _guard1854 = early_reset_static_par0_go_out;
wire _guard1855 = early_reset_static_par0_go_out;
wire _guard1856 = early_reset_static_par0_go_out;
wire _guard1857 = early_reset_static_par0_go_out;
wire _guard1858 = ~_guard0;
wire _guard1859 = early_reset_static_par0_go_out;
wire _guard1860 = _guard1858 & _guard1859;
wire _guard1861 = early_reset_static_par0_go_out;
wire _guard1862 = early_reset_static_par0_go_out;
wire _guard1863 = early_reset_static_par0_go_out;
wire _guard1864 = early_reset_static_par0_go_out;
wire _guard1865 = early_reset_static_par0_go_out;
wire _guard1866 = ~_guard0;
wire _guard1867 = early_reset_static_par0_go_out;
wire _guard1868 = _guard1866 & _guard1867;
wire _guard1869 = early_reset_static_par0_go_out;
wire _guard1870 = ~_guard0;
wire _guard1871 = early_reset_static_par0_go_out;
wire _guard1872 = _guard1870 & _guard1871;
wire _guard1873 = early_reset_static_par0_go_out;
wire _guard1874 = wrapper_early_reset_static_par_go_out;
wire _guard1875 = early_reset_static_par_go_out;
wire _guard1876 = early_reset_static_par_go_out;
wire _guard1877 = early_reset_static_par0_go_out;
wire _guard1878 = early_reset_static_par0_go_out;
wire _guard1879 = early_reset_static_par0_go_out;
wire _guard1880 = early_reset_static_par0_go_out;
wire _guard1881 = early_reset_static_par0_go_out;
wire _guard1882 = early_reset_static_par0_go_out;
wire _guard1883 = early_reset_static_par0_go_out;
wire _guard1884 = early_reset_static_par0_go_out;
wire _guard1885 = cond_wire_out;
wire _guard1886 = early_reset_static_par0_go_out;
wire _guard1887 = _guard1885 & _guard1886;
wire _guard1888 = cond_wire_out;
wire _guard1889 = early_reset_static_par0_go_out;
wire _guard1890 = _guard1888 & _guard1889;
wire _guard1891 = cond_wire26_out;
wire _guard1892 = early_reset_static_par0_go_out;
wire _guard1893 = _guard1891 & _guard1892;
wire _guard1894 = cond_wire24_out;
wire _guard1895 = early_reset_static_par0_go_out;
wire _guard1896 = _guard1894 & _guard1895;
wire _guard1897 = fsm_out == 1'd0;
wire _guard1898 = cond_wire24_out;
wire _guard1899 = _guard1897 & _guard1898;
wire _guard1900 = fsm_out == 1'd0;
wire _guard1901 = _guard1899 & _guard1900;
wire _guard1902 = fsm_out == 1'd0;
wire _guard1903 = cond_wire26_out;
wire _guard1904 = _guard1902 & _guard1903;
wire _guard1905 = fsm_out == 1'd0;
wire _guard1906 = _guard1904 & _guard1905;
wire _guard1907 = _guard1901 | _guard1906;
wire _guard1908 = early_reset_static_par0_go_out;
wire _guard1909 = _guard1907 & _guard1908;
wire _guard1910 = fsm_out == 1'd0;
wire _guard1911 = cond_wire24_out;
wire _guard1912 = _guard1910 & _guard1911;
wire _guard1913 = fsm_out == 1'd0;
wire _guard1914 = _guard1912 & _guard1913;
wire _guard1915 = fsm_out == 1'd0;
wire _guard1916 = cond_wire26_out;
wire _guard1917 = _guard1915 & _guard1916;
wire _guard1918 = fsm_out == 1'd0;
wire _guard1919 = _guard1917 & _guard1918;
wire _guard1920 = _guard1914 | _guard1919;
wire _guard1921 = early_reset_static_par0_go_out;
wire _guard1922 = _guard1920 & _guard1921;
wire _guard1923 = fsm_out == 1'd0;
wire _guard1924 = cond_wire24_out;
wire _guard1925 = _guard1923 & _guard1924;
wire _guard1926 = fsm_out == 1'd0;
wire _guard1927 = _guard1925 & _guard1926;
wire _guard1928 = fsm_out == 1'd0;
wire _guard1929 = cond_wire26_out;
wire _guard1930 = _guard1928 & _guard1929;
wire _guard1931 = fsm_out == 1'd0;
wire _guard1932 = _guard1930 & _guard1931;
wire _guard1933 = _guard1927 | _guard1932;
wire _guard1934 = early_reset_static_par0_go_out;
wire _guard1935 = _guard1933 & _guard1934;
wire _guard1936 = early_reset_static_par0_go_out;
wire _guard1937 = early_reset_static_par0_go_out;
wire _guard1938 = early_reset_static_par0_go_out;
wire _guard1939 = early_reset_static_par0_go_out;
wire _guard1940 = early_reset_static_par0_go_out;
wire _guard1941 = early_reset_static_par0_go_out;
wire _guard1942 = early_reset_static_par0_go_out;
wire _guard1943 = early_reset_static_par0_go_out;
wire _guard1944 = early_reset_static_par_go_out;
wire _guard1945 = early_reset_static_par0_go_out;
wire _guard1946 = _guard1944 | _guard1945;
wire _guard1947 = early_reset_static_par_go_out;
wire _guard1948 = early_reset_static_par0_go_out;
wire _guard1949 = early_reset_static_par0_go_out;
wire _guard1950 = early_reset_static_par0_go_out;
wire _guard1951 = early_reset_static_par0_go_out;
wire _guard1952 = ~_guard0;
wire _guard1953 = early_reset_static_par0_go_out;
wire _guard1954 = _guard1952 & _guard1953;
wire _guard1955 = early_reset_static_par0_go_out;
wire _guard1956 = early_reset_static_par0_go_out;
wire _guard1957 = early_reset_static_par0_go_out;
wire _guard1958 = early_reset_static_par0_go_out;
wire _guard1959 = early_reset_static_par0_go_out;
wire _guard1960 = early_reset_static_par0_go_out;
wire _guard1961 = early_reset_static_par0_go_out;
wire _guard1962 = ~_guard0;
wire _guard1963 = early_reset_static_par0_go_out;
wire _guard1964 = _guard1962 & _guard1963;
wire _guard1965 = ~_guard0;
wire _guard1966 = early_reset_static_par0_go_out;
wire _guard1967 = _guard1965 & _guard1966;
wire _guard1968 = early_reset_static_par0_go_out;
wire _guard1969 = early_reset_static_par0_go_out;
wire _guard1970 = early_reset_static_par0_go_out;
wire _guard1971 = ~_guard0;
wire _guard1972 = early_reset_static_par0_go_out;
wire _guard1973 = _guard1971 & _guard1972;
wire _guard1974 = early_reset_static_par0_go_out;
wire _guard1975 = cond_wire1_out;
wire _guard1976 = early_reset_static_par0_go_out;
wire _guard1977 = _guard1975 & _guard1976;
wire _guard1978 = cond_wire1_out;
wire _guard1979 = early_reset_static_par0_go_out;
wire _guard1980 = _guard1978 & _guard1979;
wire _guard1981 = cond_wire47_out;
wire _guard1982 = early_reset_static_par0_go_out;
wire _guard1983 = _guard1981 & _guard1982;
wire _guard1984 = cond_wire45_out;
wire _guard1985 = early_reset_static_par0_go_out;
wire _guard1986 = _guard1984 & _guard1985;
wire _guard1987 = fsm_out == 1'd0;
wire _guard1988 = cond_wire45_out;
wire _guard1989 = _guard1987 & _guard1988;
wire _guard1990 = fsm_out == 1'd0;
wire _guard1991 = _guard1989 & _guard1990;
wire _guard1992 = fsm_out == 1'd0;
wire _guard1993 = cond_wire47_out;
wire _guard1994 = _guard1992 & _guard1993;
wire _guard1995 = fsm_out == 1'd0;
wire _guard1996 = _guard1994 & _guard1995;
wire _guard1997 = _guard1991 | _guard1996;
wire _guard1998 = early_reset_static_par0_go_out;
wire _guard1999 = _guard1997 & _guard1998;
wire _guard2000 = fsm_out == 1'd0;
wire _guard2001 = cond_wire45_out;
wire _guard2002 = _guard2000 & _guard2001;
wire _guard2003 = fsm_out == 1'd0;
wire _guard2004 = _guard2002 & _guard2003;
wire _guard2005 = fsm_out == 1'd0;
wire _guard2006 = cond_wire47_out;
wire _guard2007 = _guard2005 & _guard2006;
wire _guard2008 = fsm_out == 1'd0;
wire _guard2009 = _guard2007 & _guard2008;
wire _guard2010 = _guard2004 | _guard2009;
wire _guard2011 = early_reset_static_par0_go_out;
wire _guard2012 = _guard2010 & _guard2011;
wire _guard2013 = fsm_out == 1'd0;
wire _guard2014 = cond_wire45_out;
wire _guard2015 = _guard2013 & _guard2014;
wire _guard2016 = fsm_out == 1'd0;
wire _guard2017 = _guard2015 & _guard2016;
wire _guard2018 = fsm_out == 1'd0;
wire _guard2019 = cond_wire47_out;
wire _guard2020 = _guard2018 & _guard2019;
wire _guard2021 = fsm_out == 1'd0;
wire _guard2022 = _guard2020 & _guard2021;
wire _guard2023 = _guard2017 | _guard2022;
wire _guard2024 = early_reset_static_par0_go_out;
wire _guard2025 = _guard2023 & _guard2024;
wire _guard2026 = cond_wire36_out;
wire _guard2027 = early_reset_static_par0_go_out;
wire _guard2028 = _guard2026 & _guard2027;
wire _guard2029 = cond_wire36_out;
wire _guard2030 = early_reset_static_par0_go_out;
wire _guard2031 = _guard2029 & _guard2030;
wire _guard2032 = early_reset_static_par_go_out;
wire _guard2033 = early_reset_static_par0_go_out;
wire _guard2034 = _guard2032 | _guard2033;
wire _guard2035 = early_reset_static_par_go_out;
wire _guard2036 = early_reset_static_par0_go_out;
wire _guard2037 = early_reset_static_par0_go_out;
wire _guard2038 = early_reset_static_par0_go_out;
wire _guard2039 = early_reset_static_par0_go_out;
wire _guard2040 = early_reset_static_par0_go_out;
wire _guard2041 = early_reset_static_par_go_out;
wire _guard2042 = early_reset_static_par0_go_out;
wire _guard2043 = _guard2041 | _guard2042;
wire _guard2044 = early_reset_static_par0_go_out;
wire _guard2045 = early_reset_static_par_go_out;
wire _guard2046 = early_reset_static_par0_go_out;
wire _guard2047 = early_reset_static_par0_go_out;
wire _guard2048 = early_reset_static_par0_go_out;
wire _guard2049 = early_reset_static_par0_go_out;
wire _guard2050 = early_reset_static_par_go_out;
wire _guard2051 = early_reset_static_par0_go_out;
wire _guard2052 = _guard2050 | _guard2051;
wire _guard2053 = early_reset_static_par0_go_out;
wire _guard2054 = early_reset_static_par_go_out;
wire _guard2055 = ~_guard0;
wire _guard2056 = early_reset_static_par0_go_out;
wire _guard2057 = _guard2055 & _guard2056;
wire _guard2058 = early_reset_static_par0_go_out;
wire _guard2059 = ~_guard0;
wire _guard2060 = early_reset_static_par0_go_out;
wire _guard2061 = _guard2059 & _guard2060;
wire _guard2062 = early_reset_static_par0_go_out;
wire _guard2063 = early_reset_static_par0_go_out;
wire _guard2064 = early_reset_static_par0_go_out;
wire _guard2065 = early_reset_static_par0_go_out;
wire _guard2066 = early_reset_static_par0_go_out;
wire _guard2067 = ~_guard0;
wire _guard2068 = early_reset_static_par0_go_out;
wire _guard2069 = _guard2067 & _guard2068;
wire _guard2070 = early_reset_static_par0_go_out;
wire _guard2071 = early_reset_static_par0_go_out;
wire _guard2072 = early_reset_static_par0_go_out;
wire _guard2073 = while_wrapper_early_reset_static_par0_done_out;
wire _guard2074 = ~_guard2073;
wire _guard2075 = fsm0_out == 2'd1;
wire _guard2076 = _guard2074 & _guard2075;
wire _guard2077 = tdcc_go_out;
wire _guard2078 = _guard2076 & _guard2077;
wire _guard2079 = cond_reg_out;
wire _guard2080 = ~_guard2079;
wire _guard2081 = fsm_out == 1'd0;
wire _guard2082 = _guard2080 & _guard2081;
assign min_depth_4_plus_5_left = min_depth_4_out;
assign min_depth_4_plus_5_right = 32'd5;
assign t3_add_left = 3'd1;
assign t3_add_right = t3_idx_out;
assign l1_add_left = 3'd1;
assign l1_add_right = l1_idx_out;
assign idx_between_depth_plus_8_depth_plus_9_reg_write_en = _guard17;
assign idx_between_depth_plus_8_depth_plus_9_reg_clk = clk;
assign idx_between_depth_plus_8_depth_plus_9_reg_reset = reset;
assign idx_between_depth_plus_8_depth_plus_9_reg_in =
  _guard18 ? idx_between_depth_plus_8_depth_plus_9_comb_out :
  _guard19 ? 1'd0 :
  'x;
assign idx_between_11_depth_plus_11_reg_write_en = _guard22;
assign idx_between_11_depth_plus_11_reg_clk = clk;
assign idx_between_11_depth_plus_11_reg_reset = reset;
assign idx_between_11_depth_plus_11_reg_in =
  _guard23 ? idx_between_11_depth_plus_11_comb_out :
  _guard24 ? 1'd0 :
  'x;
assign cond_wire3_in =
  _guard25 ? idx_between_depth_plus_5_depth_plus_6_reg_out :
  _guard28 ? cond3_out :
  1'd0;
assign cond_wire30_in =
  _guard31 ? cond30_out :
  _guard32 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire38_in =
  _guard33 ? idx_between_3_depth_plus_3_reg_out :
  _guard36 ? cond38_out :
  1'd0;
assign cond_wire39_in =
  _guard37 ? idx_between_7_depth_plus_7_reg_out :
  _guard40 ? cond39_out :
  1'd0;
assign cond_wire47_in =
  _guard41 ? idx_between_9_depth_plus_9_reg_out :
  _guard44 ? cond47_out :
  1'd0;
assign cond53_write_en = _guard45;
assign cond53_clk = clk;
assign cond53_reset = reset;
assign cond53_in =
  _guard46 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond_wire54_in =
  _guard49 ? cond54_out :
  _guard50 ? idx_between_4_min_depth_4_plus_4_reg_out :
  1'd0;
assign cond65_write_en = _guard51;
assign cond65_clk = clk;
assign cond65_reset = reset;
assign cond65_in =
  _guard52 ? idx_between_depth_plus_10_depth_plus_11_reg_out :
  1'd0;
assign left_0_3_write_en = _guard55;
assign left_0_3_clk = clk;
assign left_0_3_reset = reset;
assign left_0_3_in = left_0_2_out;
assign top_1_0_write_en = _guard61;
assign top_1_0_clk = clk;
assign top_1_0_reset = reset;
assign top_1_0_in = top_0_0_out;
assign pe_1_2_mul_ready =
  _guard67 ? 1'd1 :
  _guard70 ? 1'd0 :
  1'd0;
assign pe_1_2_clk = clk;
assign pe_1_2_top =
  _guard83 ? top_1_2_out :
  32'd0;
assign pe_1_2_left =
  _guard96 ? left_1_2_out :
  32'd0;
assign pe_1_2_reset = reset;
assign pe_1_2_go = _guard109;
assign pe_1_3_mul_ready =
  _guard112 ? 1'd1 :
  _guard115 ? 1'd0 :
  1'd0;
assign pe_1_3_clk = clk;
assign pe_1_3_top =
  _guard128 ? top_1_3_out :
  32'd0;
assign pe_1_3_left =
  _guard141 ? left_1_3_out :
  32'd0;
assign pe_1_3_reset = reset;
assign pe_1_3_go = _guard154;
assign left_1_3_write_en = _guard157;
assign left_1_3_clk = clk;
assign left_1_3_reset = reset;
assign left_1_3_in = left_1_2_out;
assign l3_idx_write_en = _guard165;
assign l3_idx_clk = clk;
assign l3_idx_reset = reset;
assign l3_idx_in =
  _guard168 ? l3_add_out :
  _guard169 ? 3'd0 :
  'x;
assign index_lt_depth_plus_9_left = idx_add_out;
assign index_lt_depth_plus_9_right = depth_plus_9_out;
assign index_lt_min_depth_4_plus_2_left = idx_add_out;
assign index_lt_min_depth_4_plus_2_right = min_depth_4_plus_2_out;
assign index_lt_min_depth_4_plus_3_left = idx_add_out;
assign index_lt_min_depth_4_plus_3_right = min_depth_4_plus_3_out;
assign index_lt_depth_plus_6_left = idx_add_out;
assign index_lt_depth_plus_6_right = depth_plus_6_out;
assign index_ge_8_left = idx_add_out;
assign index_ge_8_right = 32'd8;
assign idx_between_depth_plus_6_depth_plus_7_reg_write_en = _guard182;
assign idx_between_depth_plus_6_depth_plus_7_reg_clk = clk;
assign idx_between_depth_plus_6_depth_plus_7_reg_reset = reset;
assign idx_between_depth_plus_6_depth_plus_7_reg_in =
  _guard183 ? idx_between_depth_plus_6_depth_plus_7_comb_out :
  _guard184 ? 1'd0 :
  'x;
assign t2_addr0 =
  _guard187 ? t2_idx_out :
  3'd0;
assign done = _guard188;
assign l0_addr0 =
  _guard191 ? l0_idx_out :
  3'd0;
assign out_mem_1_addr0 =
  _guard194 ? 32'd0 :
  _guard197 ? 32'd2 :
  _guard200 ? 32'd1 :
  _guard203 ? 32'd3 :
  32'd0;
assign out_mem_0_write_data =
  _guard206 ? pe_0_1_out :
  _guard209 ? pe_0_3_out :
  _guard212 ? pe_0_2_out :
  _guard215 ? pe_0_0_out :
  32'd0;
assign out_mem_3_write_data =
  _guard218 ? pe_3_2_out :
  _guard221 ? pe_3_0_out :
  _guard224 ? pe_3_1_out :
  _guard227 ? pe_3_3_out :
  32'd0;
assign l1_addr0 =
  _guard230 ? l1_idx_out :
  3'd0;
assign l3_addr0 =
  _guard233 ? l3_idx_out :
  3'd0;
assign out_mem_2_write_data =
  _guard236 ? pe_2_1_out :
  _guard239 ? pe_2_3_out :
  _guard242 ? pe_2_0_out :
  _guard245 ? pe_2_2_out :
  32'd0;
assign out_mem_1_write_data =
  _guard248 ? pe_1_2_out :
  _guard251 ? pe_1_3_out :
  _guard254 ? pe_1_0_out :
  _guard257 ? pe_1_1_out :
  32'd0;
assign out_mem_1_write_en = _guard282;
assign t0_addr0 =
  _guard285 ? t0_idx_out :
  3'd0;
assign t1_addr0 =
  _guard288 ? t1_idx_out :
  3'd0;
assign out_mem_0_write_en = _guard313;
assign out_mem_2_write_en = _guard338;
assign out_mem_3_write_en = _guard363;
assign l2_addr0 =
  _guard366 ? l2_idx_out :
  3'd0;
assign out_mem_0_addr0 =
  _guard369 ? 32'd0 :
  _guard372 ? 32'd2 :
  _guard375 ? 32'd1 :
  _guard378 ? 32'd3 :
  32'd0;
assign out_mem_3_addr0 =
  _guard381 ? 32'd0 :
  _guard384 ? 32'd2 :
  _guard387 ? 32'd1 :
  _guard390 ? 32'd3 :
  32'd0;
assign t3_addr0 =
  _guard393 ? t3_idx_out :
  3'd0;
assign out_mem_2_addr0 =
  _guard396 ? 32'd0 :
  _guard399 ? 32'd2 :
  _guard402 ? 32'd1 :
  _guard405 ? 32'd3 :
  32'd0;
assign cond_wire0_in =
  _guard406 ? idx_between_1_min_depth_4_plus_1_reg_out :
  _guard409 ? cond0_out :
  1'd0;
assign cond_wire4_in =
  _guard412 ? cond4_out :
  _guard413 ? idx_between_1_depth_plus_1_reg_out :
  1'd0;
assign cond6_write_en = _guard414;
assign cond6_clk = clk;
assign cond6_reset = reset;
assign cond6_in =
  _guard415 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond_wire13_in =
  _guard418 ? cond13_out :
  _guard419 ? idx_between_depth_plus_7_depth_plus_8_reg_out :
  1'd0;
assign cond_wire16_in =
  _guard422 ? cond16_out :
  _guard423 ? idx_between_4_depth_plus_4_reg_out :
  1'd0;
assign cond30_write_en = _guard424;
assign cond30_clk = clk;
assign cond30_reset = reset;
assign cond30_in =
  _guard425 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire32_in =
  _guard428 ? cond32_out :
  _guard429 ? idx_between_5_min_depth_4_plus_5_reg_out :
  1'd0;
assign cond_wire40_in =
  _guard432 ? cond40_out :
  _guard433 ? idx_between_depth_plus_7_depth_plus_8_reg_out :
  1'd0;
assign cond44_write_en = _guard434;
assign cond44_clk = clk;
assign cond44_reset = reset;
assign cond44_in =
  _guard435 ? idx_between_depth_plus_8_depth_plus_9_reg_out :
  1'd0;
assign cond45_write_en = _guard436;
assign cond45_clk = clk;
assign cond45_reset = reset;
assign cond45_in =
  _guard437 ? idx_between_5_min_depth_4_plus_5_reg_out :
  1'd0;
assign fsm_write_en = _guard440;
assign fsm_clk = clk;
assign fsm_reset = reset;
assign fsm_in =
  _guard443 ? adder_out :
  _guard450 ? 1'd0 :
  _guard453 ? adder0_out :
  1'd0;
assign adder_left =
  _guard454 ? fsm_out :
  1'd0;
assign adder_right = _guard455;
assign early_reset_static_par0_go_in = _guard456;
assign depth_plus_10_left = depth;
assign depth_plus_10_right = 32'd10;
assign depth_plus_4_left = depth;
assign depth_plus_4_right = 32'd4;
assign l0_idx_write_en = _guard465;
assign l0_idx_clk = clk;
assign l0_idx_reset = reset;
assign l0_idx_in =
  _guard468 ? l0_add_out :
  _guard469 ? 3'd0 :
  'x;
assign idx_between_3_min_depth_4_plus_3_comb_left = index_ge_3_out;
assign idx_between_3_min_depth_4_plus_3_comb_right = index_lt_min_depth_4_plus_3_out;
assign index_ge_depth_plus_9_left = idx_add_out;
assign index_ge_depth_plus_9_right = depth_plus_9_out;
assign idx_between_1_min_depth_4_plus_1_reg_write_en = _guard476;
assign idx_between_1_min_depth_4_plus_1_reg_clk = clk;
assign idx_between_1_min_depth_4_plus_1_reg_reset = reset;
assign idx_between_1_min_depth_4_plus_1_reg_in =
  _guard477 ? 1'd0 :
  _guard478 ? idx_between_1_min_depth_4_plus_1_comb_out :
  'x;
assign cond11_write_en = _guard479;
assign cond11_clk = clk;
assign cond11_reset = reset;
assign cond11_in =
  _guard480 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond15_write_en = _guard481;
assign cond15_clk = clk;
assign cond15_reset = reset;
assign cond15_in =
  _guard482 ? idx_between_4_min_depth_4_plus_4_reg_out :
  1'd0;
assign cond_wire27_in =
  _guard485 ? cond27_out :
  _guard486 ? idx_between_depth_plus_7_depth_plus_8_reg_out :
  1'd0;
assign cond43_write_en = _guard487;
assign cond43_clk = clk;
assign cond43_reset = reset;
assign cond43_in =
  _guard488 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire43_in =
  _guard491 ? cond43_out :
  _guard492 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire44_in =
  _guard493 ? idx_between_depth_plus_8_depth_plus_9_reg_out :
  _guard496 ? cond44_out :
  1'd0;
assign cond62_write_en = _guard497;
assign cond62_clk = clk;
assign cond62_reset = reset;
assign cond62_in =
  _guard498 ? idx_between_6_min_depth_4_plus_6_reg_out :
  1'd0;
assign cond_wire63_in =
  _guard501 ? cond63_out :
  _guard502 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire67_in =
  _guard503 ? idx_between_11_depth_plus_11_reg_out :
  _guard506 ? cond67_out :
  1'd0;
assign pe_0_1_mul_ready =
  _guard509 ? 1'd1 :
  _guard512 ? 1'd0 :
  1'd0;
assign pe_0_1_clk = clk;
assign pe_0_1_top =
  _guard525 ? top_0_1_out :
  32'd0;
assign pe_0_1_left =
  _guard538 ? left_0_1_out :
  32'd0;
assign pe_0_1_reset = reset;
assign pe_0_1_go = _guard551;
assign left_1_2_write_en = _guard554;
assign left_1_2_clk = clk;
assign left_1_2_reset = reset;
assign left_1_2_in = left_1_1_out;
assign left_2_2_write_en = _guard560;
assign left_2_2_clk = clk;
assign left_2_2_reset = reset;
assign left_2_2_in = left_2_1_out;
assign l3_add_left = 3'd1;
assign l3_add_right = l3_idx_out;
assign idx_between_11_depth_plus_11_comb_left = index_ge_11_out;
assign idx_between_11_depth_plus_11_comb_right = index_lt_depth_plus_11_out;
assign index_lt_min_depth_4_plus_7_left = idx_add_out;
assign index_lt_min_depth_4_plus_7_right = min_depth_4_plus_7_out;
assign index_ge_3_left = idx_add_out;
assign index_ge_3_right = 32'd3;
assign index_lt_depth_plus_4_left = idx_add_out;
assign index_lt_depth_plus_4_right = depth_plus_4_out;
assign idx_between_5_depth_plus_5_comb_left = index_ge_5_out;
assign idx_between_5_depth_plus_5_comb_right = index_lt_depth_plus_5_out;
assign cond_write_en = _guard580;
assign cond_clk = clk;
assign cond_reset = reset;
assign cond_in =
  _guard581 ? idx_between_0_depth_plus_0_reg_out :
  1'd0;
assign cond_wire26_in =
  _guard582 ? idx_between_7_depth_plus_7_reg_out :
  _guard585 ? cond26_out :
  1'd0;
assign cond35_write_en = _guard586;
assign cond35_clk = clk;
assign cond35_reset = reset;
assign cond35_in =
  _guard587 ? idx_between_depth_plus_9_depth_plus_10_reg_out :
  1'd0;
assign cond_wire35_in =
  _guard590 ? cond35_out :
  _guard591 ? idx_between_depth_plus_9_depth_plus_10_reg_out :
  1'd0;
assign cond_wire50_in =
  _guard594 ? cond50_out :
  _guard595 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire56_in =
  _guard598 ? cond56_out :
  _guard599 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond60_write_en = _guard600;
assign cond60_clk = clk;
assign cond60_reset = reset;
assign cond60_in =
  _guard601 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign depth_plus_5_left = depth;
assign depth_plus_5_right = 32'd5;
assign pe_1_0_mul_ready =
  _guard606 ? 1'd1 :
  _guard609 ? 1'd0 :
  1'd0;
assign pe_1_0_clk = clk;
assign pe_1_0_top =
  _guard622 ? top_1_0_out :
  32'd0;
assign pe_1_0_left =
  _guard635 ? left_1_0_out :
  32'd0;
assign pe_1_0_reset = reset;
assign pe_1_0_go = _guard648;
assign left_1_0_write_en = _guard651;
assign left_1_0_clk = clk;
assign left_1_0_reset = reset;
assign left_1_0_in = l1_read_data;
assign left_1_1_write_en = _guard657;
assign left_1_1_clk = clk;
assign left_1_1_reset = reset;
assign left_1_1_in = left_1_0_out;
assign top_1_2_write_en = _guard663;
assign top_1_2_clk = clk;
assign top_1_2_reset = reset;
assign top_1_2_in = top_0_2_out;
assign left_2_0_write_en = _guard669;
assign left_2_0_clk = clk;
assign left_2_0_reset = reset;
assign left_2_0_in = l2_read_data;
assign left_3_1_write_en = _guard675;
assign left_3_1_clk = clk;
assign left_3_1_reset = reset;
assign left_3_1_in = left_3_0_out;
assign pe_3_2_mul_ready =
  _guard681 ? 1'd1 :
  _guard684 ? 1'd0 :
  1'd0;
assign pe_3_2_clk = clk;
assign pe_3_2_top =
  _guard697 ? top_3_2_out :
  32'd0;
assign pe_3_2_left =
  _guard710 ? left_3_2_out :
  32'd0;
assign pe_3_2_reset = reset;
assign pe_3_2_go = _guard723;
assign t1_idx_write_en = _guard728;
assign t1_idx_clk = clk;
assign t1_idx_reset = reset;
assign t1_idx_in =
  _guard731 ? t1_add_out :
  _guard732 ? 3'd0 :
  'x;
assign idx_between_depth_plus_8_depth_plus_9_comb_left = index_ge_depth_plus_8_out;
assign idx_between_depth_plus_8_depth_plus_9_comb_right = index_lt_depth_plus_9_out;
assign idx_between_7_min_depth_4_plus_7_comb_left = index_ge_7_out;
assign idx_between_7_min_depth_4_plus_7_comb_right = index_lt_min_depth_4_plus_7_out;
assign idx_between_depth_plus_9_depth_plus_10_reg_write_en = _guard739;
assign idx_between_depth_plus_9_depth_plus_10_reg_clk = clk;
assign idx_between_depth_plus_9_depth_plus_10_reg_reset = reset;
assign idx_between_depth_plus_9_depth_plus_10_reg_in =
  _guard740 ? 1'd0 :
  _guard741 ? idx_between_depth_plus_9_depth_plus_10_comb_out :
  'x;
assign index_lt_depth_plus_10_left = idx_add_out;
assign index_lt_depth_plus_10_right = depth_plus_10_out;
assign idx_between_depth_plus_6_depth_plus_7_comb_left = index_ge_depth_plus_6_out;
assign idx_between_depth_plus_6_depth_plus_7_comb_right = index_lt_depth_plus_7_out;
assign cond18_write_en = _guard746;
assign cond18_clk = clk;
assign cond18_reset = reset;
assign cond18_in =
  _guard747 ? idx_between_depth_plus_8_depth_plus_9_reg_out :
  1'd0;
assign cond_wire24_in =
  _guard748 ? idx_between_3_min_depth_4_plus_3_reg_out :
  _guard751 ? cond24_out :
  1'd0;
assign cond_wire31_in =
  _guard752 ? idx_between_depth_plus_8_depth_plus_9_reg_out :
  _guard755 ? cond31_out :
  1'd0;
assign cond_wire46_in =
  _guard758 ? cond46_out :
  _guard759 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond_wire48_in =
  _guard760 ? idx_between_depth_plus_9_depth_plus_10_reg_out :
  _guard763 ? cond48_out :
  1'd0;
assign min_depth_4_plus_2_left = min_depth_4_out;
assign min_depth_4_plus_2_right = 32'd2;
assign depth_plus_1_left = depth;
assign depth_plus_1_right = 32'd1;
assign depth_plus_12_left = depth;
assign depth_plus_12_right = 32'd12;
assign left_0_0_write_en = _guard772;
assign left_0_0_clk = clk;
assign left_0_0_reset = reset;
assign left_0_0_in = l0_read_data;
assign pe_0_3_mul_ready =
  _guard778 ? 1'd1 :
  _guard781 ? 1'd0 :
  1'd0;
assign pe_0_3_clk = clk;
assign pe_0_3_top =
  _guard794 ? top_0_3_out :
  32'd0;
assign pe_0_3_left =
  _guard807 ? left_0_3_out :
  32'd0;
assign pe_0_3_reset = reset;
assign pe_0_3_go = _guard820;
assign top_1_3_write_en = _guard823;
assign top_1_3_clk = clk;
assign top_1_3_reset = reset;
assign top_1_3_in = top_0_3_out;
assign left_2_3_write_en = _guard829;
assign left_2_3_clk = clk;
assign left_2_3_reset = reset;
assign left_2_3_in = left_2_2_out;
assign pe_3_0_mul_ready =
  _guard835 ? 1'd1 :
  _guard838 ? 1'd0 :
  1'd0;
assign pe_3_0_clk = clk;
assign pe_3_0_top =
  _guard851 ? top_3_0_out :
  32'd0;
assign pe_3_0_left =
  _guard864 ? left_3_0_out :
  32'd0;
assign pe_3_0_reset = reset;
assign pe_3_0_go = _guard877;
assign top_3_2_write_en = _guard880;
assign top_3_2_clk = clk;
assign top_3_2_reset = reset;
assign top_3_2_in = top_2_2_out;
assign idx_between_7_min_depth_4_plus_7_reg_write_en = _guard886;
assign idx_between_7_min_depth_4_plus_7_reg_clk = clk;
assign idx_between_7_min_depth_4_plus_7_reg_reset = reset;
assign idx_between_7_min_depth_4_plus_7_reg_in =
  _guard887 ? idx_between_7_min_depth_4_plus_7_comb_out :
  _guard888 ? 1'd0 :
  'x;
assign idx_between_depth_plus_5_depth_plus_6_reg_write_en = _guard891;
assign idx_between_depth_plus_5_depth_plus_6_reg_clk = clk;
assign idx_between_depth_plus_5_depth_plus_6_reg_reset = reset;
assign idx_between_depth_plus_5_depth_plus_6_reg_in =
  _guard892 ? 1'd0 :
  _guard893 ? idx_between_depth_plus_5_depth_plus_6_comb_out :
  'x;
assign index_lt_depth_plus_8_left = idx_add_out;
assign index_lt_depth_plus_8_right = depth_plus_8_out;
assign idx_between_6_min_depth_4_plus_6_comb_left = index_ge_6_out;
assign idx_between_6_min_depth_4_plus_6_comb_right = index_lt_min_depth_4_plus_6_out;
assign cond_wire18_in =
  _guard898 ? idx_between_depth_plus_8_depth_plus_9_reg_out :
  _guard901 ? cond18_out :
  1'd0;
assign cond19_write_en = _guard902;
assign cond19_clk = clk;
assign cond19_reset = reset;
assign cond19_in =
  _guard903 ? idx_between_1_depth_plus_1_reg_out :
  1'd0;
assign cond_wire29_in =
  _guard906 ? cond29_out :
  _guard907 ? idx_between_4_depth_plus_4_reg_out :
  1'd0;
assign cond34_write_en = _guard908;
assign cond34_clk = clk;
assign cond34_reset = reset;
assign cond34_in =
  _guard909 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond40_write_en = _guard910;
assign cond40_clk = clk;
assign cond40_reset = reset;
assign cond40_in =
  _guard911 ? idx_between_depth_plus_7_depth_plus_8_reg_out :
  1'd0;
assign cond57_write_en = _guard912;
assign cond57_clk = clk;
assign cond57_reset = reset;
assign cond57_in =
  _guard913 ? idx_between_depth_plus_8_depth_plus_9_reg_out :
  1'd0;
assign cond_wire59_in =
  _guard914 ? idx_between_5_depth_plus_5_reg_out :
  _guard917 ? cond59_out :
  1'd0;
assign cond_wire61_in =
  _guard918 ? idx_between_depth_plus_9_depth_plus_10_reg_out :
  _guard921 ? cond61_out :
  1'd0;
assign wrapper_early_reset_static_par_go_in = _guard927;
assign depth_plus_7_left = depth;
assign depth_plus_7_right = 32'd7;
assign pe_0_2_mul_ready =
  _guard932 ? 1'd1 :
  _guard935 ? 1'd0 :
  1'd0;
assign pe_0_2_clk = clk;
assign pe_0_2_top =
  _guard948 ? top_0_2_out :
  32'd0;
assign pe_0_2_left =
  _guard961 ? left_0_2_out :
  32'd0;
assign pe_0_2_reset = reset;
assign pe_0_2_go = _guard974;
assign t0_idx_write_en = _guard979;
assign t0_idx_clk = clk;
assign t0_idx_reset = reset;
assign t0_idx_in =
  _guard982 ? t0_add_out :
  _guard983 ? 3'd0 :
  'x;
assign l1_idx_write_en = _guard988;
assign l1_idx_clk = clk;
assign l1_idx_reset = reset;
assign l1_idx_in =
  _guard991 ? l1_add_out :
  _guard992 ? 3'd0 :
  'x;
assign idx_add_left = idx_out;
assign idx_add_right = 32'd1;
assign idx_between_2_min_depth_4_plus_2_comb_left = index_ge_2_out;
assign idx_between_2_min_depth_4_plus_2_comb_right = index_lt_min_depth_4_plus_2_out;
assign index_ge_7_left = idx_add_out;
assign index_ge_7_right = 32'd7;
assign idx_between_6_min_depth_4_plus_6_reg_write_en = _guard1001;
assign idx_between_6_min_depth_4_plus_6_reg_clk = clk;
assign idx_between_6_min_depth_4_plus_6_reg_reset = reset;
assign idx_between_6_min_depth_4_plus_6_reg_in =
  _guard1002 ? idx_between_6_min_depth_4_plus_6_comb_out :
  _guard1003 ? 1'd0 :
  'x;
assign cond3_write_en = _guard1004;
assign cond3_clk = clk;
assign cond3_reset = reset;
assign cond3_in =
  _guard1005 ? idx_between_depth_plus_5_depth_plus_6_reg_out :
  1'd0;
assign cond13_write_en = _guard1006;
assign cond13_clk = clk;
assign cond13_reset = reset;
assign cond13_in =
  _guard1007 ? idx_between_depth_plus_7_depth_plus_8_reg_out :
  1'd0;
assign cond29_write_en = _guard1008;
assign cond29_clk = clk;
assign cond29_reset = reset;
assign cond29_in =
  _guard1009 ? idx_between_4_depth_plus_4_reg_out :
  1'd0;
assign cond41_write_en = _guard1010;
assign cond41_clk = clk;
assign cond41_reset = reset;
assign cond41_in =
  _guard1011 ? idx_between_4_min_depth_4_plus_4_reg_out :
  1'd0;
assign cond54_write_en = _guard1012;
assign cond54_clk = clk;
assign cond54_reset = reset;
assign cond54_in =
  _guard1013 ? idx_between_4_min_depth_4_plus_4_reg_out :
  1'd0;
assign cond64_write_en = _guard1014;
assign cond64_clk = clk;
assign cond64_reset = reset;
assign cond64_in =
  _guard1015 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond67_write_en = _guard1016;
assign cond67_clk = clk;
assign cond67_reset = reset;
assign cond67_in =
  _guard1017 ? idx_between_11_depth_plus_11_reg_out :
  1'd0;
assign cond68_write_en = _guard1018;
assign cond68_clk = clk;
assign cond68_reset = reset;
assign cond68_in =
  _guard1019 ? idx_between_depth_plus_11_depth_plus_12_reg_out :
  1'd0;
assign wrapper_early_reset_static_par_done_in = _guard1022;
assign early_reset_static_par0_done_in = ud0_out;
assign tdcc_go_in = go;
assign pe_2_1_mul_ready =
  _guard1025 ? 1'd1 :
  _guard1028 ? 1'd0 :
  1'd0;
assign pe_2_1_clk = clk;
assign pe_2_1_top =
  _guard1041 ? top_2_1_out :
  32'd0;
assign pe_2_1_left =
  _guard1054 ? left_2_1_out :
  32'd0;
assign pe_2_1_reset = reset;
assign pe_2_1_go = _guard1067;
assign pe_2_3_mul_ready =
  _guard1070 ? 1'd1 :
  _guard1073 ? 1'd0 :
  1'd0;
assign pe_2_3_clk = clk;
assign pe_2_3_top =
  _guard1086 ? top_2_3_out :
  32'd0;
assign pe_2_3_left =
  _guard1099 ? left_2_3_out :
  32'd0;
assign pe_2_3_reset = reset;
assign pe_2_3_go = _guard1112;
assign pe_3_1_mul_ready =
  _guard1115 ? 1'd1 :
  _guard1118 ? 1'd0 :
  1'd0;
assign pe_3_1_clk = clk;
assign pe_3_1_top =
  _guard1131 ? top_3_1_out :
  32'd0;
assign pe_3_1_left =
  _guard1144 ? left_3_1_out :
  32'd0;
assign pe_3_1_reset = reset;
assign pe_3_1_go = _guard1157;
assign lt_iter_limit_left =
  _guard1158 ? depth :
  _guard1159 ? idx_add_out :
  'x;
assign lt_iter_limit_right =
  _guard1160 ? 32'd4 :
  _guard1161 ? iter_limit_out :
  'x;
assign idx_between_7_depth_plus_7_comb_left = index_ge_7_out;
assign idx_between_7_depth_plus_7_comb_right = index_lt_depth_plus_7_out;
assign idx_between_6_depth_plus_6_comb_left = index_ge_6_out;
assign idx_between_6_depth_plus_6_comb_right = index_lt_depth_plus_6_out;
assign index_ge_depth_plus_7_left = idx_add_out;
assign index_ge_depth_plus_7_right = depth_plus_7_out;
assign cond17_write_en = _guard1168;
assign cond17_clk = clk;
assign cond17_reset = reset;
assign cond17_in =
  _guard1169 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire22_in =
  _guard1170 ? idx_between_6_depth_plus_6_reg_out :
  _guard1173 ? cond22_out :
  1'd0;
assign cond23_write_en = _guard1174;
assign cond23_clk = clk;
assign cond23_reset = reset;
assign cond23_in =
  _guard1175 ? idx_between_depth_plus_6_depth_plus_7_reg_out :
  1'd0;
assign cond25_write_en = _guard1176;
assign cond25_clk = clk;
assign cond25_reset = reset;
assign cond25_in =
  _guard1177 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond_wire33_in =
  _guard1180 ? cond33_out :
  _guard1181 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond52_write_en = _guard1182;
assign cond52_clk = clk;
assign cond52_reset = reset;
assign cond52_in =
  _guard1183 ? idx_between_depth_plus_10_depth_plus_11_reg_out :
  1'd0;
assign cond56_write_en = _guard1184;
assign cond56_clk = clk;
assign cond56_reset = reset;
assign cond56_in =
  _guard1185 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond58_write_en = _guard1186;
assign cond58_clk = clk;
assign cond58_reset = reset;
assign cond58_in =
  _guard1187 ? idx_between_5_min_depth_4_plus_5_reg_out :
  1'd0;
assign fsm0_write_en = _guard1200;
assign fsm0_clk = clk;
assign fsm0_reset = reset;
assign fsm0_in =
  _guard1205 ? 2'd1 :
  _guard1206 ? 2'd0 :
  _guard1211 ? 2'd2 :
  2'd0;
assign depth_plus_8_left =
  _guard1212 ? depth :
  _guard1213 ? 32'd12 :
  'x;
assign depth_plus_8_right =
  _guard1214 ? depth :
  _guard1215 ? 32'd8 :
  'x;
assign min_depth_4_plus_4_left = min_depth_4_out;
assign min_depth_4_plus_4_right = 32'd4;
assign depth_plus_0_left = depth;
assign depth_plus_0_right = 32'd0;
assign top_2_0_write_en = _guard1222;
assign top_2_0_clk = clk;
assign top_2_0_reset = reset;
assign top_2_0_in = top_1_0_out;
assign top_3_0_write_en = _guard1228;
assign top_3_0_clk = clk;
assign top_3_0_reset = reset;
assign top_3_0_in = top_2_0_out;
assign top_3_1_write_en = _guard1234;
assign top_3_1_clk = clk;
assign top_3_1_reset = reset;
assign top_3_1_in = top_2_1_out;
assign idx_write_en = _guard1240;
assign idx_clk = clk;
assign idx_reset = reset;
assign idx_in =
  _guard1241 ? 32'd0 :
  _guard1242 ? idx_add_out :
  'x;
assign idx_between_7_depth_plus_7_reg_write_en = _guard1245;
assign idx_between_7_depth_plus_7_reg_clk = clk;
assign idx_between_7_depth_plus_7_reg_reset = reset;
assign idx_between_7_depth_plus_7_reg_in =
  _guard1246 ? idx_between_7_depth_plus_7_comb_out :
  _guard1247 ? 1'd0 :
  'x;
assign index_lt_depth_plus_3_left = idx_add_out;
assign index_lt_depth_plus_3_right = depth_plus_3_out;
assign idx_between_depth_plus_10_depth_plus_11_reg_write_en = _guard1252;
assign idx_between_depth_plus_10_depth_plus_11_reg_clk = clk;
assign idx_between_depth_plus_10_depth_plus_11_reg_reset = reset;
assign idx_between_depth_plus_10_depth_plus_11_reg_in =
  _guard1253 ? 1'd0 :
  _guard1254 ? idx_between_depth_plus_10_depth_plus_11_comb_out :
  'x;
assign idx_between_4_depth_plus_4_comb_left = index_ge_4_out;
assign idx_between_4_depth_plus_4_comb_right = index_lt_depth_plus_4_out;
assign index_lt_min_depth_4_plus_5_left = idx_add_out;
assign index_lt_min_depth_4_plus_5_right = min_depth_4_plus_5_out;
assign index_lt_depth_plus_0_left = idx_add_out;
assign index_lt_depth_plus_0_right = depth_plus_0_out;
assign idx_between_9_depth_plus_9_reg_write_en = _guard1263;
assign idx_between_9_depth_plus_9_reg_clk = clk;
assign idx_between_9_depth_plus_9_reg_reset = reset;
assign idx_between_9_depth_plus_9_reg_in =
  _guard1264 ? 1'd0 :
  _guard1265 ? idx_between_9_depth_plus_9_comb_out :
  'x;
assign idx_between_1_depth_plus_1_comb_left = index_ge_1_out;
assign idx_between_1_depth_plus_1_comb_right = index_lt_depth_plus_1_out;
assign index_ge_depth_plus_11_left = idx_add_out;
assign index_ge_depth_plus_11_right = depth_plus_11_out;
assign idx_between_depth_plus_11_depth_plus_12_comb_left = index_ge_depth_plus_11_out;
assign idx_between_depth_plus_11_depth_plus_12_comb_right = index_lt_depth_plus_12_out;
assign cond7_write_en = _guard1272;
assign cond7_clk = clk;
assign cond7_reset = reset;
assign cond7_in =
  _guard1273 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire8_in =
  _guard1274 ? idx_between_depth_plus_6_depth_plus_7_reg_out :
  _guard1277 ? cond8_out :
  1'd0;
assign cond9_write_en = _guard1278;
assign cond9_clk = clk;
assign cond9_reset = reset;
assign cond9_in =
  _guard1279 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond14_write_en = _guard1280;
assign cond14_clk = clk;
assign cond14_reset = reset;
assign cond14_in =
  _guard1281 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond_wire20_in =
  _guard1284 ? cond20_out :
  _guard1285 ? idx_between_2_min_depth_4_plus_2_reg_out :
  1'd0;
assign cond27_write_en = _guard1286;
assign cond27_clk = clk;
assign cond27_reset = reset;
assign cond27_in =
  _guard1287 ? idx_between_depth_plus_7_depth_plus_8_reg_out :
  1'd0;
assign cond32_write_en = _guard1288;
assign cond32_clk = clk;
assign cond32_reset = reset;
assign cond32_in =
  _guard1289 ? idx_between_5_min_depth_4_plus_5_reg_out :
  1'd0;
assign cond_wire37_in =
  _guard1290 ? idx_between_3_min_depth_4_plus_3_reg_out :
  _guard1293 ? cond37_out :
  1'd0;
assign cond50_write_en = _guard1294;
assign cond50_clk = clk;
assign cond50_reset = reset;
assign cond50_in =
  _guard1295 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire60_in =
  _guard1298 ? cond60_out :
  _guard1299 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond_wire64_in =
  _guard1302 ? cond64_out :
  _guard1303 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign min_depth_4_write_en = _guard1304;
assign min_depth_4_clk = clk;
assign min_depth_4_reset = reset;
assign min_depth_4_in =
  _guard1307 ? depth :
  _guard1311 ? 32'd4 :
  'x;
assign min_depth_4_plus_6_left = min_depth_4_out;
assign min_depth_4_plus_6_right = 32'd6;
assign top_0_1_write_en = _guard1316;
assign top_0_1_clk = clk;
assign top_0_1_reset = reset;
assign top_0_1_in = t1_read_data;
assign left_0_2_write_en = _guard1322;
assign left_0_2_clk = clk;
assign left_0_2_reset = reset;
assign left_0_2_in = left_0_1_out;
assign top_2_3_write_en = _guard1328;
assign top_2_3_clk = clk;
assign top_2_3_reset = reset;
assign top_2_3_in = top_1_3_out;
assign left_3_0_write_en = _guard1334;
assign left_3_0_clk = clk;
assign left_3_0_reset = reset;
assign left_3_0_in = l3_read_data;
assign idx_between_3_min_depth_4_plus_3_reg_write_en = _guard1340;
assign idx_between_3_min_depth_4_plus_3_reg_clk = clk;
assign idx_between_3_min_depth_4_plus_3_reg_reset = reset;
assign idx_between_3_min_depth_4_plus_3_reg_in =
  _guard1341 ? idx_between_3_min_depth_4_plus_3_comb_out :
  _guard1342 ? 1'd0 :
  'x;
assign index_ge_4_left = idx_add_out;
assign index_ge_4_right = 32'd4;
assign idx_between_5_min_depth_4_plus_5_reg_write_en = _guard1347;
assign idx_between_5_min_depth_4_plus_5_reg_clk = clk;
assign idx_between_5_min_depth_4_plus_5_reg_reset = reset;
assign idx_between_5_min_depth_4_plus_5_reg_in =
  _guard1348 ? 1'd0 :
  _guard1349 ? idx_between_5_min_depth_4_plus_5_comb_out :
  'x;
assign index_ge_1_left = idx_add_out;
assign index_ge_1_right = 32'd1;
assign cond4_write_en = _guard1352;
assign cond4_clk = clk;
assign cond4_reset = reset;
assign cond4_in =
  _guard1353 ? idx_between_1_depth_plus_1_reg_out :
  1'd0;
assign cond5_write_en = _guard1354;
assign cond5_clk = clk;
assign cond5_reset = reset;
assign cond5_in =
  _guard1355 ? idx_between_2_min_depth_4_plus_2_reg_out :
  1'd0;
assign cond_wire6_in =
  _guard1358 ? cond6_out :
  _guard1359 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond20_write_en = _guard1360;
assign cond20_clk = clk;
assign cond20_reset = reset;
assign cond20_in =
  _guard1361 ? idx_between_2_min_depth_4_plus_2_reg_out :
  1'd0;
assign cond_wire36_in =
  _guard1364 ? cond36_out :
  _guard1365 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond46_write_en = _guard1366;
assign cond46_clk = clk;
assign cond46_reset = reset;
assign cond46_in =
  _guard1367 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond_wire62_in =
  _guard1370 ? cond62_out :
  _guard1371 ? idx_between_6_min_depth_4_plus_6_reg_out :
  1'd0;
assign cond63_write_en = _guard1372;
assign cond63_clk = clk;
assign cond63_reset = reset;
assign cond63_in =
  _guard1373 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire66_in =
  _guard1374 ? idx_between_7_min_depth_4_plus_7_reg_out :
  _guard1377 ? cond66_out :
  1'd0;
assign adder0_left =
  _guard1378 ? fsm_out :
  1'd0;
assign adder0_right = _guard1379;
assign early_reset_static_par_done_in = ud_out;
assign depth_plus_3_left = depth;
assign depth_plus_3_right = 32'd3;
assign top_0_2_write_en = _guard1384;
assign top_0_2_clk = clk;
assign top_0_2_reset = reset;
assign top_0_2_in = t2_read_data;
assign top_1_1_write_en = _guard1390;
assign top_1_1_clk = clk;
assign top_1_1_reset = reset;
assign top_1_1_in = top_0_1_out;
assign left_3_2_write_en = _guard1396;
assign left_3_2_clk = clk;
assign left_3_2_reset = reset;
assign left_3_2_in = left_3_1_out;
assign t0_add_left = 3'd1;
assign t0_add_right = t0_idx_out;
assign l0_add_left = 3'd1;
assign l0_add_right = l0_idx_out;
assign index_ge_11_left = idx_add_out;
assign index_ge_11_right = 32'd11;
assign index_ge_9_left = idx_add_out;
assign index_ge_9_right = 32'd9;
assign idx_between_1_min_depth_4_plus_1_comb_left = index_ge_1_out;
assign idx_between_1_min_depth_4_plus_1_comb_right = index_lt_min_depth_4_plus_1_out;
assign idx_between_depth_plus_7_depth_plus_8_comb_left = index_ge_depth_plus_7_out;
assign idx_between_depth_plus_7_depth_plus_8_comb_right = index_lt_depth_plus_8_out;
assign cond_wire2_in =
  _guard1422 ? cond2_out :
  _guard1423 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond_wire9_in =
  _guard1426 ? cond9_out :
  _guard1427 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond10_write_en = _guard1428;
assign cond10_clk = clk;
assign cond10_reset = reset;
assign cond10_in =
  _guard1429 ? idx_between_3_min_depth_4_plus_3_reg_out :
  1'd0;
assign cond_wire11_in =
  _guard1432 ? cond11_out :
  _guard1433 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond21_write_en = _guard1434;
assign cond21_clk = clk;
assign cond21_reset = reset;
assign cond21_in =
  _guard1435 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond24_write_en = _guard1436;
assign cond24_clk = clk;
assign cond24_reset = reset;
assign cond24_in =
  _guard1437 ? idx_between_3_min_depth_4_plus_3_reg_out :
  1'd0;
assign cond31_write_en = _guard1438;
assign cond31_clk = clk;
assign cond31_reset = reset;
assign cond31_in =
  _guard1439 ? idx_between_depth_plus_8_depth_plus_9_reg_out :
  1'd0;
assign cond36_write_en = _guard1440;
assign cond36_clk = clk;
assign cond36_reset = reset;
assign cond36_in =
  _guard1441 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond_wire41_in =
  _guard1444 ? cond41_out :
  _guard1445 ? idx_between_4_min_depth_4_plus_4_reg_out :
  1'd0;
assign cond_wire45_in =
  _guard1448 ? cond45_out :
  _guard1449 ? idx_between_5_min_depth_4_plus_5_reg_out :
  1'd0;
assign cond51_write_en = _guard1450;
assign cond51_clk = clk;
assign cond51_reset = reset;
assign cond51_in =
  _guard1451 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond_wire57_in =
  _guard1452 ? idx_between_depth_plus_8_depth_plus_9_reg_out :
  _guard1455 ? cond57_out :
  1'd0;
assign cond_wire58_in =
  _guard1458 ? cond58_out :
  _guard1459 ? idx_between_5_min_depth_4_plus_5_reg_out :
  1'd0;
assign cond61_write_en = _guard1460;
assign cond61_clk = clk;
assign cond61_reset = reset;
assign cond61_in =
  _guard1461 ? idx_between_depth_plus_9_depth_plus_10_reg_out :
  1'd0;
assign signal_reg_write_en = _guard1471;
assign signal_reg_clk = clk;
assign signal_reg_reset = reset;
assign signal_reg_in =
  _guard1477 ? 1'd1 :
  _guard1480 ? 1'd0 :
  1'd0;
assign depth_plus_9_left = depth;
assign depth_plus_9_right = 32'd9;
assign depth_plus_6_left = depth;
assign depth_plus_6_right = 32'd6;
assign pe_2_0_mul_ready =
  _guard1487 ? 1'd1 :
  _guard1490 ? 1'd0 :
  1'd0;
assign pe_2_0_clk = clk;
assign pe_2_0_top =
  _guard1503 ? top_2_0_out :
  32'd0;
assign pe_2_0_left =
  _guard1516 ? left_2_0_out :
  32'd0;
assign pe_2_0_reset = reset;
assign pe_2_0_go = _guard1529;
assign left_2_1_write_en = _guard1532;
assign left_2_1_clk = clk;
assign left_2_1_reset = reset;
assign left_2_1_in = left_2_0_out;
assign top_2_2_write_en = _guard1538;
assign top_2_2_clk = clk;
assign top_2_2_reset = reset;
assign top_2_2_in = top_1_2_out;
assign t1_add_left = 3'd1;
assign t1_add_right = t1_idx_out;
assign t3_idx_write_en = _guard1552;
assign t3_idx_clk = clk;
assign t3_idx_reset = reset;
assign t3_idx_in =
  _guard1555 ? t3_add_out :
  _guard1556 ? 3'd0 :
  'x;
assign index_ge_2_left = idx_add_out;
assign index_ge_2_right = 32'd2;
assign index_lt_depth_plus_11_left = idx_add_out;
assign index_lt_depth_plus_11_right = depth_plus_11_out;
assign index_lt_depth_plus_7_left = idx_add_out;
assign index_lt_depth_plus_7_right = depth_plus_7_out;
assign idx_between_6_depth_plus_6_reg_write_en = _guard1565;
assign idx_between_6_depth_plus_6_reg_clk = clk;
assign idx_between_6_depth_plus_6_reg_reset = reset;
assign idx_between_6_depth_plus_6_reg_in =
  _guard1566 ? idx_between_6_depth_plus_6_comb_out :
  _guard1567 ? 1'd0 :
  'x;
assign idx_between_4_min_depth_4_plus_4_comb_left = index_ge_4_out;
assign idx_between_4_min_depth_4_plus_4_comb_right = index_lt_min_depth_4_plus_4_out;
assign idx_between_5_min_depth_4_plus_5_comb_left = index_ge_5_out;
assign idx_between_5_min_depth_4_plus_5_comb_right = index_lt_min_depth_4_plus_5_out;
assign idx_between_0_depth_plus_0_reg_write_en = _guard1574;
assign idx_between_0_depth_plus_0_reg_clk = clk;
assign idx_between_0_depth_plus_0_reg_reset = reset;
assign idx_between_0_depth_plus_0_reg_in =
  _guard1575 ? 1'd1 :
  _guard1576 ? index_lt_depth_plus_0_out :
  'x;
assign idx_between_10_depth_plus_10_comb_left = index_ge_10_out;
assign idx_between_10_depth_plus_10_comb_right = index_lt_depth_plus_10_out;
assign idx_between_depth_plus_7_depth_plus_8_reg_write_en = _guard1581;
assign idx_between_depth_plus_7_depth_plus_8_reg_clk = clk;
assign idx_between_depth_plus_7_depth_plus_8_reg_reset = reset;
assign idx_between_depth_plus_7_depth_plus_8_reg_in =
  _guard1582 ? 1'd0 :
  _guard1583 ? idx_between_depth_plus_7_depth_plus_8_comb_out :
  'x;
assign cond_wire_in =
  _guard1586 ? cond_out :
  _guard1587 ? idx_between_0_depth_plus_0_reg_out :
  1'd0;
assign cond_wire15_in =
  _guard1590 ? cond15_out :
  _guard1591 ? idx_between_4_min_depth_4_plus_4_reg_out :
  1'd0;
assign cond16_write_en = _guard1592;
assign cond16_clk = clk;
assign cond16_reset = reset;
assign cond16_in =
  _guard1593 ? idx_between_4_depth_plus_4_reg_out :
  1'd0;
assign cond37_write_en = _guard1594;
assign cond37_clk = clk;
assign cond37_reset = reset;
assign cond37_in =
  _guard1595 ? idx_between_3_min_depth_4_plus_3_reg_out :
  1'd0;
assign cond_wire49_in =
  _guard1596 ? idx_between_6_min_depth_4_plus_6_reg_out :
  _guard1599 ? cond49_out :
  1'd0;
assign cond_wire55_in =
  _guard1600 ? idx_between_4_depth_plus_4_reg_out :
  _guard1603 ? cond55_out :
  1'd0;
assign depth_plus_2_left = depth;
assign depth_plus_2_right = 32'd2;
assign pe_0_0_mul_ready =
  _guard1608 ? 1'd1 :
  _guard1611 ? 1'd0 :
  1'd0;
assign pe_0_0_clk = clk;
assign pe_0_0_top =
  _guard1624 ? top_0_0_out :
  32'd0;
assign pe_0_0_left =
  _guard1637 ? left_0_0_out :
  32'd0;
assign pe_0_0_reset = reset;
assign pe_0_0_go = _guard1650;
assign pe_3_3_mul_ready =
  _guard1653 ? 1'd1 :
  _guard1656 ? 1'd0 :
  1'd0;
assign pe_3_3_clk = clk;
assign pe_3_3_top =
  _guard1669 ? top_3_3_out :
  32'd0;
assign pe_3_3_left =
  _guard1682 ? left_3_3_out :
  32'd0;
assign pe_3_3_reset = reset;
assign pe_3_3_go = _guard1695;
assign top_3_3_write_en = _guard1698;
assign top_3_3_clk = clk;
assign top_3_3_reset = reset;
assign top_3_3_in = top_2_3_out;
assign t2_add_left = 3'd1;
assign t2_add_right = t2_idx_out;
assign idx_between_2_min_depth_4_plus_2_reg_write_en = _guard1710;
assign idx_between_2_min_depth_4_plus_2_reg_clk = clk;
assign idx_between_2_min_depth_4_plus_2_reg_reset = reset;
assign idx_between_2_min_depth_4_plus_2_reg_in =
  _guard1711 ? idx_between_2_min_depth_4_plus_2_comb_out :
  _guard1712 ? 1'd0 :
  'x;
assign idx_between_2_depth_plus_2_reg_write_en = _guard1715;
assign idx_between_2_depth_plus_2_reg_clk = clk;
assign idx_between_2_depth_plus_2_reg_reset = reset;
assign idx_between_2_depth_plus_2_reg_in =
  _guard1716 ? 1'd0 :
  _guard1717 ? idx_between_2_depth_plus_2_comb_out :
  'x;
assign idx_between_2_depth_plus_2_comb_left = index_ge_2_out;
assign idx_between_2_depth_plus_2_comb_right = index_lt_depth_plus_2_out;
assign idx_between_3_depth_plus_3_reg_write_en = _guard1722;
assign idx_between_3_depth_plus_3_reg_clk = clk;
assign idx_between_3_depth_plus_3_reg_reset = reset;
assign idx_between_3_depth_plus_3_reg_in =
  _guard1723 ? 1'd0 :
  _guard1724 ? idx_between_3_depth_plus_3_comb_out :
  'x;
assign idx_between_depth_plus_9_depth_plus_10_comb_left = index_ge_depth_plus_9_out;
assign idx_between_depth_plus_9_depth_plus_10_comb_right = index_lt_depth_plus_10_out;
assign idx_between_8_depth_plus_8_reg_write_en = _guard1729;
assign idx_between_8_depth_plus_8_reg_clk = clk;
assign idx_between_8_depth_plus_8_reg_reset = reset;
assign idx_between_8_depth_plus_8_reg_in =
  _guard1730 ? 1'd0 :
  _guard1731 ? idx_between_8_depth_plus_8_comb_out :
  'x;
assign index_ge_depth_plus_10_left = idx_add_out;
assign index_ge_depth_plus_10_right = depth_plus_10_out;
assign index_ge_depth_plus_6_left = idx_add_out;
assign index_ge_depth_plus_6_right = depth_plus_6_out;
assign idx_between_4_depth_plus_4_reg_write_en = _guard1738;
assign idx_between_4_depth_plus_4_reg_clk = clk;
assign idx_between_4_depth_plus_4_reg_reset = reset;
assign idx_between_4_depth_plus_4_reg_in =
  _guard1739 ? idx_between_4_depth_plus_4_comb_out :
  _guard1740 ? 1'd0 :
  'x;
assign index_lt_min_depth_4_plus_4_left = idx_add_out;
assign index_lt_min_depth_4_plus_4_right = min_depth_4_plus_4_out;
assign index_ge_5_left = idx_add_out;
assign index_ge_5_right = 32'd5;
assign index_lt_depth_plus_12_left = idx_add_out;
assign index_lt_depth_plus_12_right = depth_plus_12_out;
assign idx_between_10_depth_plus_10_reg_write_en = _guard1749;
assign idx_between_10_depth_plus_10_reg_clk = clk;
assign idx_between_10_depth_plus_10_reg_reset = reset;
assign idx_between_10_depth_plus_10_reg_in =
  _guard1750 ? 1'd0 :
  _guard1751 ? idx_between_10_depth_plus_10_comb_out :
  'x;
assign index_ge_10_left = idx_add_out;
assign index_ge_10_right = 32'd10;
assign index_lt_min_depth_4_plus_6_left = idx_add_out;
assign index_lt_min_depth_4_plus_6_right = min_depth_4_plus_6_out;
assign cond0_write_en = _guard1756;
assign cond0_clk = clk;
assign cond0_reset = reset;
assign cond0_in =
  _guard1757 ? idx_between_1_min_depth_4_plus_1_reg_out :
  1'd0;
assign cond_wire7_in =
  _guard1760 ? cond7_out :
  _guard1761 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond_wire10_in =
  _guard1762 ? idx_between_3_min_depth_4_plus_3_reg_out :
  _guard1765 ? cond10_out :
  1'd0;
assign cond_wire12_in =
  _guard1766 ? idx_between_7_depth_plus_7_reg_out :
  _guard1769 ? cond12_out :
  1'd0;
assign cond_wire17_in =
  _guard1772 ? cond17_out :
  _guard1773 ? idx_between_8_depth_plus_8_reg_out :
  1'd0;
assign cond_wire19_in =
  _guard1776 ? cond19_out :
  _guard1777 ? idx_between_1_depth_plus_1_reg_out :
  1'd0;
assign cond_wire23_in =
  _guard1778 ? idx_between_depth_plus_6_depth_plus_7_reg_out :
  _guard1781 ? cond23_out :
  1'd0;
assign cond_wire25_in =
  _guard1784 ? cond25_out :
  _guard1785 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond33_write_en = _guard1786;
assign cond33_clk = clk;
assign cond33_reset = reset;
assign cond33_in =
  _guard1787 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond_wire42_in =
  _guard1788 ? idx_between_4_depth_plus_4_reg_out :
  _guard1791 ? cond42_out :
  1'd0;
assign cond47_write_en = _guard1792;
assign cond47_clk = clk;
assign cond47_reset = reset;
assign cond47_in =
  _guard1793 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond48_write_en = _guard1794;
assign cond48_clk = clk;
assign cond48_reset = reset;
assign cond48_in =
  _guard1795 ? idx_between_depth_plus_9_depth_plus_10_reg_out :
  1'd0;
assign cond66_write_en = _guard1796;
assign cond66_clk = clk;
assign cond66_reset = reset;
assign cond66_in =
  _guard1797 ? idx_between_7_min_depth_4_plus_7_reg_out :
  1'd0;
assign tdcc_done_in = _guard1798;
assign top_0_3_write_en = _guard1801;
assign top_0_3_clk = clk;
assign top_0_3_reset = reset;
assign top_0_3_in = t3_read_data;
assign top_2_1_write_en = _guard1807;
assign top_2_1_clk = clk;
assign top_2_1_reset = reset;
assign top_2_1_in = top_1_1_out;
assign left_3_3_write_en = _guard1813;
assign left_3_3_clk = clk;
assign left_3_3_reset = reset;
assign left_3_3_in = left_3_2_out;
assign t2_idx_write_en = _guard1821;
assign t2_idx_clk = clk;
assign t2_idx_reset = reset;
assign t2_idx_in =
  _guard1824 ? t2_add_out :
  _guard1825 ? 3'd0 :
  'x;
assign l2_idx_write_en = _guard1830;
assign l2_idx_clk = clk;
assign l2_idx_reset = reset;
assign l2_idx_in =
  _guard1831 ? 3'd0 :
  _guard1834 ? l2_add_out :
  'x;
assign index_ge_depth_plus_5_left = idx_add_out;
assign index_ge_depth_plus_5_right = depth_plus_5_out;
assign index_ge_6_left = idx_add_out;
assign index_ge_6_right = 32'd6;
assign index_lt_depth_plus_5_left = idx_add_out;
assign index_lt_depth_plus_5_right = depth_plus_5_out;
assign idx_between_1_depth_plus_1_reg_write_en = _guard1843;
assign idx_between_1_depth_plus_1_reg_clk = clk;
assign idx_between_1_depth_plus_1_reg_reset = reset;
assign idx_between_1_depth_plus_1_reg_in =
  _guard1844 ? idx_between_1_depth_plus_1_comb_out :
  _guard1845 ? 1'd0 :
  'x;
assign cond1_write_en = _guard1846;
assign cond1_clk = clk;
assign cond1_reset = reset;
assign cond1_in =
  _guard1847 ? idx_between_1_depth_plus_1_reg_out :
  1'd0;
assign cond2_write_en = _guard1848;
assign cond2_clk = clk;
assign cond2_reset = reset;
assign cond2_in =
  _guard1849 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign cond_wire5_in =
  _guard1852 ? cond5_out :
  _guard1853 ? idx_between_2_min_depth_4_plus_2_reg_out :
  1'd0;
assign cond22_write_en = _guard1854;
assign cond22_clk = clk;
assign cond22_reset = reset;
assign cond22_in =
  _guard1855 ? idx_between_6_depth_plus_6_reg_out :
  1'd0;
assign cond26_write_en = _guard1856;
assign cond26_clk = clk;
assign cond26_reset = reset;
assign cond26_in =
  _guard1857 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond_wire34_in =
  _guard1860 ? cond34_out :
  _guard1861 ? idx_between_9_depth_plus_9_reg_out :
  1'd0;
assign cond39_write_en = _guard1862;
assign cond39_clk = clk;
assign cond39_reset = reset;
assign cond39_in =
  _guard1863 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond49_write_en = _guard1864;
assign cond49_clk = clk;
assign cond49_reset = reset;
assign cond49_in =
  _guard1865 ? idx_between_6_min_depth_4_plus_6_reg_out :
  1'd0;
assign cond_wire52_in =
  _guard1868 ? cond52_out :
  _guard1869 ? idx_between_depth_plus_10_depth_plus_11_reg_out :
  1'd0;
assign cond_wire68_in =
  _guard1872 ? cond68_out :
  _guard1873 ? idx_between_depth_plus_11_depth_plus_12_reg_out :
  1'd0;
assign early_reset_static_par_go_in = _guard1874;
assign iter_limit_write_en = _guard1875;
assign iter_limit_clk = clk;
assign iter_limit_reset = reset;
assign iter_limit_in = depth_plus_8_out;
assign depth_plus_11_left = depth;
assign depth_plus_11_right = 32'd11;
assign min_depth_4_plus_7_left = min_depth_4_out;
assign min_depth_4_plus_7_right = 32'd7;
assign min_depth_4_plus_3_left = min_depth_4_out;
assign min_depth_4_plus_3_right = 32'd3;
assign min_depth_4_plus_1_left = min_depth_4_out;
assign min_depth_4_plus_1_right = 32'd1;
assign top_0_0_write_en = _guard1887;
assign top_0_0_clk = clk;
assign top_0_0_reset = reset;
assign top_0_0_in = t0_read_data;
assign pe_1_1_mul_ready =
  _guard1893 ? 1'd1 :
  _guard1896 ? 1'd0 :
  1'd0;
assign pe_1_1_clk = clk;
assign pe_1_1_top =
  _guard1909 ? top_1_1_out :
  32'd0;
assign pe_1_1_left =
  _guard1922 ? left_1_1_out :
  32'd0;
assign pe_1_1_reset = reset;
assign pe_1_1_go = _guard1935;
assign index_lt_depth_plus_2_left = idx_add_out;
assign index_lt_depth_plus_2_right = depth_plus_2_out;
assign idx_between_depth_plus_5_depth_plus_6_comb_left = index_ge_depth_plus_5_out;
assign idx_between_depth_plus_5_depth_plus_6_comb_right = index_lt_depth_plus_6_out;
assign idx_between_8_depth_plus_8_comb_left = index_ge_8_out;
assign idx_between_8_depth_plus_8_comb_right = index_lt_depth_plus_8_out;
assign idx_between_depth_plus_10_depth_plus_11_comb_left = index_ge_depth_plus_10_out;
assign idx_between_depth_plus_10_depth_plus_11_comb_right = index_lt_depth_plus_11_out;
assign idx_between_4_min_depth_4_plus_4_reg_write_en = _guard1946;
assign idx_between_4_min_depth_4_plus_4_reg_clk = clk;
assign idx_between_4_min_depth_4_plus_4_reg_reset = reset;
assign idx_between_4_min_depth_4_plus_4_reg_in =
  _guard1947 ? 1'd0 :
  _guard1948 ? idx_between_4_min_depth_4_plus_4_comb_out :
  'x;
assign index_lt_min_depth_4_plus_1_left = idx_add_out;
assign index_lt_min_depth_4_plus_1_right = min_depth_4_plus_1_out;
assign cond_wire1_in =
  _guard1951 ? idx_between_1_depth_plus_1_reg_out :
  _guard1954 ? cond1_out :
  1'd0;
assign cond8_write_en = _guard1955;
assign cond8_clk = clk;
assign cond8_reset = reset;
assign cond8_in =
  _guard1956 ? idx_between_depth_plus_6_depth_plus_7_reg_out :
  1'd0;
assign cond12_write_en = _guard1957;
assign cond12_clk = clk;
assign cond12_reset = reset;
assign cond12_in =
  _guard1958 ? idx_between_7_depth_plus_7_reg_out :
  1'd0;
assign cond28_write_en = _guard1959;
assign cond28_clk = clk;
assign cond28_reset = reset;
assign cond28_in =
  _guard1960 ? idx_between_4_min_depth_4_plus_4_reg_out :
  1'd0;
assign cond_wire28_in =
  _guard1961 ? idx_between_4_min_depth_4_plus_4_reg_out :
  _guard1964 ? cond28_out :
  1'd0;
assign cond_wire53_in =
  _guard1967 ? cond53_out :
  _guard1968 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond55_write_en = _guard1969;
assign cond55_clk = clk;
assign cond55_reset = reset;
assign cond55_in =
  _guard1970 ? idx_between_4_depth_plus_4_reg_out :
  1'd0;
assign cond_wire65_in =
  _guard1973 ? cond65_out :
  _guard1974 ? idx_between_depth_plus_10_depth_plus_11_reg_out :
  1'd0;
assign left_0_1_write_en = _guard1977;
assign left_0_1_clk = clk;
assign left_0_1_reset = reset;
assign left_0_1_in = left_0_0_out;
assign pe_2_2_mul_ready =
  _guard1983 ? 1'd1 :
  _guard1986 ? 1'd0 :
  1'd0;
assign pe_2_2_clk = clk;
assign pe_2_2_top =
  _guard1999 ? top_2_2_out :
  32'd0;
assign pe_2_2_left =
  _guard2012 ? left_2_2_out :
  32'd0;
assign pe_2_2_reset = reset;
assign pe_2_2_go = _guard2025;
assign l2_add_left = 3'd1;
assign l2_add_right = l2_idx_out;
assign cond_reg_write_en = _guard2034;
assign cond_reg_clk = clk;
assign cond_reg_reset = reset;
assign cond_reg_in =
  _guard2035 ? 1'd1 :
  _guard2036 ? lt_iter_limit_out :
  'x;
assign index_ge_depth_plus_8_left = idx_add_out;
assign index_ge_depth_plus_8_right = depth_plus_8_out;
assign idx_between_3_depth_plus_3_comb_left = index_ge_3_out;
assign idx_between_3_depth_plus_3_comb_right = index_lt_depth_plus_3_out;
assign idx_between_5_depth_plus_5_reg_write_en = _guard2043;
assign idx_between_5_depth_plus_5_reg_clk = clk;
assign idx_between_5_depth_plus_5_reg_reset = reset;
assign idx_between_5_depth_plus_5_reg_in =
  _guard2044 ? idx_between_5_depth_plus_5_comb_out :
  _guard2045 ? 1'd0 :
  'x;
assign idx_between_9_depth_plus_9_comb_left = index_ge_9_out;
assign idx_between_9_depth_plus_9_comb_right = index_lt_depth_plus_9_out;
assign index_lt_depth_plus_1_left = idx_add_out;
assign index_lt_depth_plus_1_right = depth_plus_1_out;
assign idx_between_depth_plus_11_depth_plus_12_reg_write_en = _guard2052;
assign idx_between_depth_plus_11_depth_plus_12_reg_clk = clk;
assign idx_between_depth_plus_11_depth_plus_12_reg_reset = reset;
assign idx_between_depth_plus_11_depth_plus_12_reg_in =
  _guard2053 ? idx_between_depth_plus_11_depth_plus_12_comb_out :
  _guard2054 ? 1'd0 :
  'x;
assign cond_wire14_in =
  _guard2057 ? cond14_out :
  _guard2058 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond_wire21_in =
  _guard2061 ? cond21_out :
  _guard2062 ? idx_between_2_depth_plus_2_reg_out :
  1'd0;
assign cond38_write_en = _guard2063;
assign cond38_clk = clk;
assign cond38_reset = reset;
assign cond38_in =
  _guard2064 ? idx_between_3_depth_plus_3_reg_out :
  1'd0;
assign cond42_write_en = _guard2065;
assign cond42_clk = clk;
assign cond42_reset = reset;
assign cond42_in =
  _guard2066 ? idx_between_4_depth_plus_4_reg_out :
  1'd0;
assign cond_wire51_in =
  _guard2069 ? cond51_out :
  _guard2070 ? idx_between_10_depth_plus_10_reg_out :
  1'd0;
assign cond59_write_en = _guard2071;
assign cond59_clk = clk;
assign cond59_reset = reset;
assign cond59_in =
  _guard2072 ? idx_between_5_depth_plus_5_reg_out :
  1'd0;
assign while_wrapper_early_reset_static_par0_go_in = _guard2078;
assign while_wrapper_early_reset_static_par0_done_in = _guard2082;
// COMPONENT END: systolic_array_comp
endmodule
module main(
  input logic go,
  input logic clk,
  input logic reset,
  output logic done,
  output logic [2:0] t0_addr0,
  output logic [31:0] t0_write_data,
  output logic t0_write_en,
  output logic t0_clk,
  output logic t0_reset,
  input logic [31:0] t0_read_data,
  input logic t0_done,
  output logic [2:0] t1_addr0,
  output logic [31:0] t1_write_data,
  output logic t1_write_en,
  output logic t1_clk,
  output logic t1_reset,
  input logic [31:0] t1_read_data,
  input logic t1_done,
  output logic [2:0] t2_addr0,
  output logic [31:0] t2_write_data,
  output logic t2_write_en,
  output logic t2_clk,
  output logic t2_reset,
  input logic [31:0] t2_read_data,
  input logic t2_done,
  output logic [2:0] t3_addr0,
  output logic [31:0] t3_write_data,
  output logic t3_write_en,
  output logic t3_clk,
  output logic t3_reset,
  input logic [31:0] t3_read_data,
  input logic t3_done,
  output logic [2:0] l0_addr0,
  output logic [31:0] l0_write_data,
  output logic l0_write_en,
  output logic l0_clk,
  output logic l0_reset,
  input logic [31:0] l0_read_data,
  input logic l0_done,
  output logic [2:0] l1_addr0,
  output logic [31:0] l1_write_data,
  output logic l1_write_en,
  output logic l1_clk,
  output logic l1_reset,
  input logic [31:0] l1_read_data,
  input logic l1_done,
  output logic [2:0] l2_addr0,
  output logic [31:0] l2_write_data,
  output logic l2_write_en,
  output logic l2_clk,
  output logic l2_reset,
  input logic [31:0] l2_read_data,
  input logic l2_done,
  output logic [2:0] l3_addr0,
  output logic [31:0] l3_write_data,
  output logic l3_write_en,
  output logic l3_clk,
  output logic l3_reset,
  input logic [31:0] l3_read_data,
  input logic l3_done,
  output logic [31:0] out_mem_0_addr0,
  output logic [31:0] out_mem_0_write_data,
  output logic out_mem_0_write_en,
  output logic out_mem_0_clk,
  output logic out_mem_0_reset,
  input logic [31:0] out_mem_0_read_data,
  input logic out_mem_0_done,
  output logic [31:0] out_mem_1_addr0,
  output logic [31:0] out_mem_1_write_data,
  output logic out_mem_1_write_en,
  output logic out_mem_1_clk,
  output logic out_mem_1_reset,
  input logic [31:0] out_mem_1_read_data,
  input logic out_mem_1_done,
  output logic [31:0] out_mem_2_addr0,
  output logic [31:0] out_mem_2_write_data,
  output logic out_mem_2_write_en,
  output logic out_mem_2_clk,
  output logic out_mem_2_reset,
  input logic [31:0] out_mem_2_read_data,
  input logic out_mem_2_done,
  output logic [31:0] out_mem_3_addr0,
  output logic [31:0] out_mem_3_write_data,
  output logic out_mem_3_write_en,
  output logic out_mem_3_clk,
  output logic out_mem_3_reset,
  input logic [31:0] out_mem_3_read_data,
  input logic out_mem_3_done
);
// COMPONENT START: main
logic [31:0] systolic_array_depth;
logic [31:0] systolic_array_t0_read_data;
logic [31:0] systolic_array_t1_read_data;
logic [31:0] systolic_array_t2_read_data;
logic [31:0] systolic_array_t3_read_data;
logic [31:0] systolic_array_l0_read_data;
logic [31:0] systolic_array_l1_read_data;
logic [31:0] systolic_array_l2_read_data;
logic [31:0] systolic_array_l3_read_data;
logic [2:0] systolic_array_t0_addr0;
logic [2:0] systolic_array_t1_addr0;
logic [2:0] systolic_array_t2_addr0;
logic [2:0] systolic_array_t3_addr0;
logic [2:0] systolic_array_l0_addr0;
logic [2:0] systolic_array_l1_addr0;
logic [2:0] systolic_array_l2_addr0;
logic [2:0] systolic_array_l3_addr0;
logic [31:0] systolic_array_out_mem_0_addr0;
logic [31:0] systolic_array_out_mem_0_write_data;
logic systolic_array_out_mem_0_write_en;
logic [31:0] systolic_array_out_mem_1_addr0;
logic [31:0] systolic_array_out_mem_1_write_data;
logic systolic_array_out_mem_1_write_en;
logic [31:0] systolic_array_out_mem_2_addr0;
logic [31:0] systolic_array_out_mem_2_write_data;
logic systolic_array_out_mem_2_write_en;
logic [31:0] systolic_array_out_mem_3_addr0;
logic [31:0] systolic_array_out_mem_3_write_data;
logic systolic_array_out_mem_3_write_en;
logic systolic_array_go;
logic systolic_array_clk;
logic systolic_array_reset;
logic systolic_array_done;
logic invoke0_go_in;
logic invoke0_go_out;
logic invoke0_done_in;
logic invoke0_done_out;
systolic_array_comp systolic_array (
    .clk(systolic_array_clk),
    .depth(systolic_array_depth),
    .done(systolic_array_done),
    .go(systolic_array_go),
    .l0_addr0(systolic_array_l0_addr0),
    .l0_read_data(systolic_array_l0_read_data),
    .l1_addr0(systolic_array_l1_addr0),
    .l1_read_data(systolic_array_l1_read_data),
    .l2_addr0(systolic_array_l2_addr0),
    .l2_read_data(systolic_array_l2_read_data),
    .l3_addr0(systolic_array_l3_addr0),
    .l3_read_data(systolic_array_l3_read_data),
    .out_mem_0_addr0(systolic_array_out_mem_0_addr0),
    .out_mem_0_write_data(systolic_array_out_mem_0_write_data),
    .out_mem_0_write_en(systolic_array_out_mem_0_write_en),
    .out_mem_1_addr0(systolic_array_out_mem_1_addr0),
    .out_mem_1_write_data(systolic_array_out_mem_1_write_data),
    .out_mem_1_write_en(systolic_array_out_mem_1_write_en),
    .out_mem_2_addr0(systolic_array_out_mem_2_addr0),
    .out_mem_2_write_data(systolic_array_out_mem_2_write_data),
    .out_mem_2_write_en(systolic_array_out_mem_2_write_en),
    .out_mem_3_addr0(systolic_array_out_mem_3_addr0),
    .out_mem_3_write_data(systolic_array_out_mem_3_write_data),
    .out_mem_3_write_en(systolic_array_out_mem_3_write_en),
    .reset(systolic_array_reset),
    .t0_addr0(systolic_array_t0_addr0),
    .t0_read_data(systolic_array_t0_read_data),
    .t1_addr0(systolic_array_t1_addr0),
    .t1_read_data(systolic_array_t1_read_data),
    .t2_addr0(systolic_array_t2_addr0),
    .t2_read_data(systolic_array_t2_read_data),
    .t3_addr0(systolic_array_t3_addr0),
    .t3_read_data(systolic_array_t3_read_data)
);
std_wire # (
    .WIDTH(1)
) invoke0_go (
    .in(invoke0_go_in),
    .out(invoke0_go_out)
);
std_wire # (
    .WIDTH(1)
) invoke0_done (
    .in(invoke0_done_in),
    .out(invoke0_done_out)
);
wire _guard0 = 1;
wire _guard1 = invoke0_go_out;
wire _guard2 = invoke0_done_out;
wire _guard3 = invoke0_go_out;
wire _guard4 = invoke0_go_out;
wire _guard5 = invoke0_go_out;
wire _guard6 = invoke0_go_out;
wire _guard7 = invoke0_go_out;
wire _guard8 = invoke0_go_out;
wire _guard9 = invoke0_go_out;
wire _guard10 = invoke0_go_out;
wire _guard11 = invoke0_go_out;
wire _guard12 = invoke0_go_out;
wire _guard13 = invoke0_go_out;
wire _guard14 = invoke0_go_out;
wire _guard15 = invoke0_go_out;
wire _guard16 = invoke0_go_out;
wire _guard17 = invoke0_go_out;
wire _guard18 = invoke0_go_out;
wire _guard19 = invoke0_go_out;
wire _guard20 = invoke0_go_out;
wire _guard21 = invoke0_go_out;
wire _guard22 = invoke0_go_out;
wire _guard23 = invoke0_go_out;
wire _guard24 = invoke0_go_out;
wire _guard25 = invoke0_go_out;
wire _guard26 = invoke0_go_out;
wire _guard27 = invoke0_go_out;
wire _guard28 = invoke0_go_out;
wire _guard29 = invoke0_go_out;
wire _guard30 = invoke0_go_out;
wire _guard31 = invoke0_go_out;
assign t2_addr0 =
  _guard1 ? systolic_array_t2_addr0 :
  3'd0;
assign done = _guard2;
assign t3_reset = reset;
assign t0_reset = reset;
assign out_mem_2_reset = reset;
assign l0_addr0 =
  _guard3 ? systolic_array_l0_addr0 :
  3'd0;
assign out_mem_1_addr0 =
  _guard4 ? systolic_array_out_mem_1_addr0 :
  32'd0;
assign t2_clk = clk;
assign l3_clk = clk;
assign out_mem_1_clk = clk;
assign out_mem_3_reset = reset;
assign out_mem_0_write_data =
  _guard5 ? systolic_array_out_mem_0_write_data :
  32'd0;
assign out_mem_3_write_data =
  _guard6 ? systolic_array_out_mem_3_write_data :
  32'd0;
assign t0_clk = clk;
assign out_mem_1_reset = reset;
assign l1_addr0 =
  _guard7 ? systolic_array_l1_addr0 :
  3'd0;
assign l0_reset = reset;
assign out_mem_0_clk = clk;
assign t1_reset = reset;
assign out_mem_3_clk = clk;
assign l3_addr0 =
  _guard8 ? systolic_array_l3_addr0 :
  3'd0;
assign out_mem_2_write_data =
  _guard9 ? systolic_array_out_mem_2_write_data :
  32'd0;
assign out_mem_1_write_data =
  _guard10 ? systolic_array_out_mem_1_write_data :
  32'd0;
assign out_mem_1_write_en =
  _guard11 ? systolic_array_out_mem_1_write_en :
  1'd0;
assign out_mem_0_reset = reset;
assign t0_addr0 =
  _guard12 ? systolic_array_t0_addr0 :
  3'd0;
assign t1_addr0 =
  _guard13 ? systolic_array_t1_addr0 :
  3'd0;
assign out_mem_0_write_en =
  _guard14 ? systolic_array_out_mem_0_write_en :
  1'd0;
assign out_mem_2_write_en =
  _guard15 ? systolic_array_out_mem_2_write_en :
  1'd0;
assign t1_clk = clk;
assign l1_reset = reset;
assign l2_clk = clk;
assign l2_reset = reset;
assign out_mem_2_clk = clk;
assign out_mem_3_write_en =
  _guard16 ? systolic_array_out_mem_3_write_en :
  1'd0;
assign t3_clk = clk;
assign l2_addr0 =
  _guard17 ? systolic_array_l2_addr0 :
  3'd0;
assign out_mem_0_addr0 =
  _guard18 ? systolic_array_out_mem_0_addr0 :
  32'd0;
assign out_mem_3_addr0 =
  _guard19 ? systolic_array_out_mem_3_addr0 :
  32'd0;
assign l0_clk = clk;
assign l1_clk = clk;
assign l3_reset = reset;
assign t3_addr0 =
  _guard20 ? systolic_array_t3_addr0 :
  3'd0;
assign out_mem_2_addr0 =
  _guard21 ? systolic_array_out_mem_2_addr0 :
  32'd0;
assign t2_reset = reset;
assign invoke0_go_in = go;
assign invoke0_done_in = systolic_array_done;
assign systolic_array_l1_read_data =
  _guard22 ? l1_read_data :
  32'd0;
assign systolic_array_l2_read_data =
  _guard23 ? l2_read_data :
  32'd0;
assign systolic_array_l3_read_data =
  _guard24 ? l3_read_data :
  32'd0;
assign systolic_array_depth =
  _guard25 ? 32'd4 :
  32'd0;
assign systolic_array_clk = clk;
assign systolic_array_t3_read_data =
  _guard26 ? t3_read_data :
  32'd0;
assign systolic_array_l0_read_data =
  _guard27 ? l0_read_data :
  32'd0;
assign systolic_array_reset = reset;
assign systolic_array_go = _guard28;
assign systolic_array_t1_read_data =
  _guard29 ? t1_read_data :
  32'd0;
assign systolic_array_t0_read_data =
  _guard30 ? t0_read_data :
  32'd0;
assign systolic_array_t2_read_data =
  _guard31 ? t2_read_data :
  32'd0;
// COMPONENT END: main
endmodule

