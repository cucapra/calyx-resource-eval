
/// This is mostly used for testing the static guarantees currently.
/// A realistic implementation would probably take four cycles.
module pipelined_mult (
    input wire clk,
    input wire reset,
    // inputs
    input wire [31:0] left,
    input wire [31:0] right,
    // The input has been committed
    output wire [31:0] out
);

logic [31:0] lt, rt, buff0, buff1, buff2, tmp_prod;

assign out = buff2;
assign tmp_prod = lt * rt;

always_ff @(posedge clk) begin
    if (reset) begin
        lt <= 0;
        rt <= 0;
        buff0 <= 0;
        buff1 <= 0;
        buff2 <= 0;
    end else begin
        lt <= left;
        rt <= right;
        buff0 <= tmp_prod;
        buff1 <= buff0;
        buff2 <= buff1;
    end
end

endmodule

module bb_pipelined_mult(
	               input wire [31:0] left,
	               input wire [31:0] right,
	               output wire [31:0] out,
	               input wire clk
	               );
`ifdef __ICARUS__
   reg [31:0] reg0;
   reg [31:0] reg1;
   reg [31:0] reg2;
   reg [31:0] reg3;
   always @( posedge clk ) begin
      reg0 <= left * right;
      reg1 <= reg0;
      reg2 <= reg1;
      reg3 <= reg2;
   end
   assign out = reg3;
`elsif VERILATOR
   reg [31:0] reg0;
   reg [31:0] reg1;
   reg [31:0] reg2;
   reg [31:0] reg3;
   always @( posedge clk ) begin
      reg0 <= left * right;
      reg1 <= reg0;
      reg2 <= reg1;
      reg3 <= reg2;
   end
   assign out = reg3;
`else
   // mul_uint32 is a black box module generated by Xilinx's IP Core generator.
   // Generation commands are in the synth.tcl file.
   mul_uint32 mul_uint32 (
                   .A(left),
                   .B(right),
                   .P(out),
                   .CLK(clk)
                   );
`endif
endmodule
/* verilator lint_off MULTITOP */
/// =================== Unsigned, Fixed Point =========================
module std_fp_add #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  assign out = left + right;
endmodule

module std_fp_sub #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module std_fp_mult_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16,
    parameter SIGNED = 0
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    input  logic             go,
    input  logic             clk,
    input  logic             reset,
    output logic [WIDTH-1:0] out,
    output logic             done
);
  logic [WIDTH-1:0]          rtmp;
  logic [WIDTH-1:0]          ltmp;
  logic [(WIDTH << 1) - 1:0] out_tmp;
  // Buffer used to walk through the 3 cycles of the pipeline.
  logic done_buf[1:0];

  assign done = done_buf[1];

  assign out = out_tmp[(WIDTH << 1) - INT_WIDTH - 1 : WIDTH - INT_WIDTH];

  // If the done buffer is completely empty and go is high then execution
  // just started.
  logic start;
  assign start = go;

  // Start sending the done signal.
  always_ff @(posedge clk) begin
    if (start)
      done_buf[0] <= 1;
    else
      done_buf[0] <= 0;
  end

  // Push the done signal through the pipeline.
  always_ff @(posedge clk) begin
    if (go) begin
      done_buf[1] <= done_buf[0];
    end else begin
      done_buf[1] <= 0;
    end
  end

  // Register the inputs
  always_ff @(posedge clk) begin
    if (reset) begin
      rtmp <= 0;
      ltmp <= 0;
    end else if (go) begin
      if (SIGNED) begin
        rtmp <= $signed(right);
        ltmp <= $signed(left);
      end else begin
        rtmp <= right;
        ltmp <= left;
      end
    end else begin
      rtmp <= 0;
      ltmp <= 0;
    end

  end

  // Compute the output and save it into out_tmp
  always_ff @(posedge clk) begin
    if (reset) begin
      out_tmp <= 0;
    end else if (go) begin
      if (SIGNED) begin
        // In the first cycle, this performs an invalid computation because
        // ltmp and rtmp only get their actual values in cycle 1
        out_tmp <= $signed(
          { {WIDTH{ltmp[WIDTH-1]}}, ltmp} *
          { {WIDTH{rtmp[WIDTH-1]}}, rtmp}
        );
      end else begin
        out_tmp <= ltmp * rtmp;
      end
    end else begin
      out_tmp <= out_tmp;
    end
  end
endmodule

/* verilator lint_off WIDTH */
module std_fp_div_pipe #(
  parameter WIDTH = 32,
  parameter INT_WIDTH = 16,
  parameter FRAC_WIDTH = 16
) (
    input  logic             go,
    input  logic             clk,
    input  logic             reset,
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out_remainder,
    output logic [WIDTH-1:0] out_quotient,
    output logic             done
);
    localparam ITERATIONS = WIDTH + FRAC_WIDTH;

    logic [WIDTH-1:0] quotient, quotient_next;
    logic [WIDTH:0] acc, acc_next;
    logic [$clog2(ITERATIONS)-1:0] idx;
    logic start, running, finished, dividend_is_zero;

    assign start = go && !running;
    assign dividend_is_zero = start && left == 0;
    assign finished = idx == ITERATIONS - 1 && running;

    always_ff @(posedge clk) begin
      if (reset || finished || dividend_is_zero)
        running <= 0;
      else if (start)
        running <= 1;
      else
        running <= running;
    end

    always_comb begin
      if (acc >= {1'b0, right}) begin
        acc_next = acc - right;
        {acc_next, quotient_next} = {acc_next[WIDTH-1:0], quotient, 1'b1};
      end else begin
        {acc_next, quotient_next} = {acc, quotient} << 1;
      end
    end

    // `done` signaling
    always_ff @(posedge clk) begin
      if (dividend_is_zero || finished)
        done <= 1;
      else
        done <= 0;
    end

    always_ff @(posedge clk) begin
      if (running)
        idx <= idx + 1;
      else
        idx <= 0;
    end

    always_ff @(posedge clk) begin
      if (reset) begin
        out_quotient <= 0;
        out_remainder <= 0;
      end else if (start) begin
        out_quotient <= 0;
        out_remainder <= left;
      end else if (go == 0) begin
        out_quotient <= out_quotient;
        out_remainder <= out_remainder;
      end else if (dividend_is_zero) begin
        out_quotient <= 0;
        out_remainder <= 0;
      end else if (finished) begin
        out_quotient <= quotient_next;
        out_remainder <= out_remainder;
      end else begin
        out_quotient <= out_quotient;
        if (right <= out_remainder)
          out_remainder <= out_remainder - right;
        else
          out_remainder <= out_remainder;
      end
    end

    always_ff @(posedge clk) begin
      if (reset) begin
        acc <= 0;
        quotient <= 0;
      end else if (start) begin
        {acc, quotient} <= {{WIDTH{1'b0}}, left, 1'b0};
      end else begin
        acc <= acc_next;
        quotient <= quotient_next;
      end
    end
endmodule

module std_fp_gt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    output logic             out
);
  assign out = left > right;
endmodule

/// =================== Signed, Fixed Point =========================
module std_fp_sadd #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left + right);
endmodule

module std_fp_ssub #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);

  assign out = $signed(left - right);
endmodule

module std_fp_smult_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  [WIDTH-1:0]              left,
    input  [WIDTH-1:0]              right,
    input  logic                    reset,
    input  logic                    go,
    input  logic                    clk,
    output logic [WIDTH-1:0]        out,
    output logic                    done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(INT_WIDTH),
    .FRAC_WIDTH(FRAC_WIDTH),
    .SIGNED(1)
  ) comp (
    .clk(clk),
    .done(done),
    .reset(reset),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

module std_fp_sdiv_pipe #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input                     clk,
    input                     go,
    input                     reset,
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out_quotient,
    output signed [WIDTH-1:0] out_remainder,
    output logic              done
);

  logic signed [WIDTH-1:0] left_abs, right_abs, comp_out_q, comp_out_r, right_save, out_rem_intermediate;

  // Registers to figure out how to transform outputs.
  logic different_signs, left_sign, right_sign;

  // Latch the value of control registers so that their available after
  // go signal becomes low.
  always_ff @(posedge clk) begin
    if (go) begin
      right_save <= right_abs;
      left_sign <= left[WIDTH-1];
      right_sign <= right[WIDTH-1];
    end else begin
      left_sign <= left_sign;
      right_save <= right_save;
      right_sign <= right_sign;
    end
  end

  assign right_abs = right[WIDTH-1] ? -right : right;
  assign left_abs = left[WIDTH-1] ? -left : left;

  assign different_signs = left_sign ^ right_sign;
  assign out_quotient = different_signs ? -comp_out_q : comp_out_q;

  // Remainder is computed as:
  //  t0 = |left| % |right|
  //  t1 = if left * right < 0 and t0 != 0 then |right| - t0 else t0
  //  rem = if right < 0 then -t1 else t1
  assign out_rem_intermediate = different_signs & |comp_out_r ? $signed(right_save - comp_out_r) : comp_out_r;
  assign out_remainder = right_sign ? -out_rem_intermediate : out_rem_intermediate;

  std_fp_div_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(INT_WIDTH),
    .FRAC_WIDTH(FRAC_WIDTH)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left_abs),
    .right(right_abs),
    .out_quotient(comp_out_q),
    .out_remainder(comp_out_r)
  );
endmodule

module std_fp_sgt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
    input  logic signed [WIDTH-1:0] left,
    input  logic signed [WIDTH-1:0] right,
    output logic signed             out
);
  assign out = $signed(left > right);
endmodule

module std_fp_slt #(
    parameter WIDTH = 32,
    parameter INT_WIDTH = 16,
    parameter FRAC_WIDTH = 16
) (
   input logic signed [WIDTH-1:0] left,
   input logic signed [WIDTH-1:0] right,
   output logic signed            out
);
  assign out = $signed(left < right);
endmodule

/// =================== Unsigned, Bitnum =========================
module std_mult_pipe #(
    parameter WIDTH = 32
) (
    input  logic [WIDTH-1:0] left,
    input  logic [WIDTH-1:0] right,
    input  logic             reset,
    input  logic             go,
    input  logic             clk,
    output logic [WIDTH-1:0] out,
    output logic             done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(WIDTH),
    .FRAC_WIDTH(0),
    .SIGNED(0)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

module std_div_pipe #(
    parameter WIDTH = 32
) (
    input                    reset,
    input                    clk,
    input                    go,
    input        [WIDTH-1:0] left,
    input        [WIDTH-1:0] right,
    output logic [WIDTH-1:0] out_remainder,
    output logic [WIDTH-1:0] out_quotient,
    output logic             done
);

  logic [WIDTH-1:0] dividend;
  logic [(WIDTH-1)*2:0] divisor;
  logic [WIDTH-1:0] quotient;
  logic [WIDTH-1:0] quotient_msk;
  logic start, running, finished, dividend_is_zero;

  assign start = go && !running;
  assign finished = quotient_msk == 0 && running;
  assign dividend_is_zero = start && left == 0;

  always_ff @(posedge clk) begin
    // Early return if the divisor is zero.
    if (finished || dividend_is_zero)
      done <= 1;
    else
      done <= 0;
  end

  always_ff @(posedge clk) begin
    if (reset || finished || dividend_is_zero)
      running <= 0;
    else if (start)
      running <= 1;
    else
      running <= running;
  end

  // Outputs
  always_ff @(posedge clk) begin
    if (dividend_is_zero || start) begin
      out_quotient <= 0;
      out_remainder <= 0;
    end else if (finished) begin
      out_quotient <= quotient;
      out_remainder <= dividend;
    end else begin
      // Otherwise, explicitly latch the values.
      out_quotient <= out_quotient;
      out_remainder <= out_remainder;
    end
  end

  // Calculate the quotient mask.
  always_ff @(posedge clk) begin
    if (start)
      quotient_msk <= 1 << WIDTH - 1;
    else if (running)
      quotient_msk <= quotient_msk >> 1;
    else
      quotient_msk <= quotient_msk;
  end

  // Calculate the quotient.
  always_ff @(posedge clk) begin
    if (start)
      quotient <= 0;
    else if (divisor <= dividend)
      quotient <= quotient | quotient_msk;
    else
      quotient <= quotient;
  end

  // Calculate the dividend.
  always_ff @(posedge clk) begin
    if (start)
      dividend <= left;
    else if (divisor <= dividend)
      dividend <= dividend - divisor;
    else
      dividend <= dividend;
  end

  always_ff @(posedge clk) begin
    if (start) begin
      divisor <= right << WIDTH - 1;
    end else if (finished) begin
      divisor <= 0;
    end else begin
      divisor <= divisor >> 1;
    end
  end

  // Simulation self test against unsynthesizable implementation.
  `ifdef VERILATOR
    logic [WIDTH-1:0] l, r;
    always_ff @(posedge clk) begin
      if (go) begin
        l <= left;
        r <= right;
      end else begin
        l <= l;
        r <= r;
      end
    end

    always @(posedge clk) begin
      if (done && $unsigned(out_remainder) != $unsigned(l % r))
        $error(
          "\nstd_div_pipe (Remainder): Computed and golden outputs do not match!\n",
          "left: %0d", $unsigned(l),
          "  right: %0d\n", $unsigned(r),
          "expected: %0d", $unsigned(l % r),
          "  computed: %0d", $unsigned(out_remainder)
        );

      if (done && $unsigned(out_quotient) != $unsigned(l / r))
        $error(
          "\nstd_div_pipe (Quotient): Computed and golden outputs do not match!\n",
          "left: %0d", $unsigned(l),
          "  right: %0d\n", $unsigned(r),
          "expected: %0d", $unsigned(l / r),
          "  computed: %0d", $unsigned(out_quotient)
        );
    end
  `endif
endmodule

/// =================== Signed, Bitnum =========================
module std_sadd #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left + right);
endmodule

module std_ssub #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = $signed(left - right);
endmodule

module std_smult_pipe #(
    parameter WIDTH = 32
) (
    input  logic                    reset,
    input  logic                    go,
    input  logic                    clk,
    input  signed       [WIDTH-1:0] left,
    input  signed       [WIDTH-1:0] right,
    output logic signed [WIDTH-1:0] out,
    output logic                    done
);
  std_fp_mult_pipe #(
    .WIDTH(WIDTH),
    .INT_WIDTH(WIDTH),
    .FRAC_WIDTH(0),
    .SIGNED(1)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left),
    .right(right),
    .out(out)
  );
endmodule

/* verilator lint_off WIDTH */
module std_sdiv_pipe #(
    parameter WIDTH = 32
) (
    input                           reset,
    input                           clk,
    input                           go,
    input  logic signed [WIDTH-1:0] left,
    input  logic signed [WIDTH-1:0] right,
    output logic signed [WIDTH-1:0] out_quotient,
    output logic signed [WIDTH-1:0] out_remainder,
    output logic                    done
);

  logic signed [WIDTH-1:0] left_abs, right_abs, comp_out_q, comp_out_r, right_save, out_rem_intermediate;

  // Registers to figure out how to transform outputs.
  logic different_signs, left_sign, right_sign;

  // Latch the value of control registers so that their available after
  // go signal becomes low.
  always_ff @(posedge clk) begin
    if (go) begin
      right_save <= right_abs;
      left_sign <= left[WIDTH-1];
      right_sign <= right[WIDTH-1];
    end else begin
      left_sign <= left_sign;
      right_save <= right_save;
      right_sign <= right_sign;
    end
  end

  assign right_abs = right[WIDTH-1] ? -right : right;
  assign left_abs = left[WIDTH-1] ? -left : left;

  assign different_signs = left_sign ^ right_sign;
  assign out_quotient = different_signs ? -comp_out_q : comp_out_q;

  // Remainder is computed as:
  //  t0 = |left| % |right|
  //  t1 = if left * right < 0 and t0 != 0 then |right| - t0 else t0
  //  rem = if right < 0 then -t1 else t1
  assign out_rem_intermediate = different_signs & |comp_out_r ? $signed(right_save - comp_out_r) : comp_out_r;
  assign out_remainder = right_sign ? -out_rem_intermediate : out_rem_intermediate;

  std_div_pipe #(
    .WIDTH(WIDTH)
  ) comp (
    .reset(reset),
    .clk(clk),
    .done(done),
    .go(go),
    .left(left_abs),
    .right(right_abs),
    .out_quotient(comp_out_q),
    .out_remainder(comp_out_r)
  );

  // Simulation self test against unsynthesizable implementation.
  `ifdef VERILATOR
    logic signed [WIDTH-1:0] l, r;
    always_ff @(posedge clk) begin
      if (go) begin
        l <= left;
        r <= right;
      end else begin
        l <= l;
        r <= r;
      end
    end

    always @(posedge clk) begin
      if (done && out_quotient != $signed(l / r))
        $error(
          "\nstd_sdiv_pipe (Quotient): Computed and golden outputs do not match!\n",
          "left: %0d", l,
          "  right: %0d\n", r,
          "expected: %0d", $signed(l / r),
          "  computed: %0d", $signed(out_quotient),
        );
      if (done && out_remainder != $signed(((l % r) + r) % r))
        $error(
          "\nstd_sdiv_pipe (Remainder): Computed and golden outputs do not match!\n",
          "left: %0d", l,
          "  right: %0d\n", r,
          "expected: %0d", $signed(((l % r) + r) % r),
          "  computed: %0d", $signed(out_remainder),
        );
    end
  `endif
endmodule

module std_sgt #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left > right);
endmodule

module std_slt #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left < right);
endmodule

module std_seq #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left == right);
endmodule

module std_sneq #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left != right);
endmodule

module std_sge #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left >= right);
endmodule

module std_sle #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed             out
);
  assign out = $signed(left <= right);
endmodule

module std_slsh #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = left <<< right;
endmodule

module std_srsh #(
    parameter WIDTH = 32
) (
    input  signed [WIDTH-1:0] left,
    input  signed [WIDTH-1:0] right,
    output signed [WIDTH-1:0] out
);
  assign out = left >>> right;
endmodule

/**
 * Core primitives for Calyx.
 * Implements core primitives used by the compiler.
 *
 * Conventions:
 * - All parameter names must be SNAKE_CASE and all caps.
 * - Port names must be snake_case, no caps.
 */
`default_nettype none

module std_slice #(
    parameter IN_WIDTH  = 32,
    parameter OUT_WIDTH = 32
) (
   input wire                   logic [ IN_WIDTH-1:0] in,
   output logic [OUT_WIDTH-1:0] out
);
  assign out = in[OUT_WIDTH-1:0];

  `ifdef VERILATOR
    always_comb begin
      if (IN_WIDTH < OUT_WIDTH)
        $error(
          "std_slice: Input width less than output width\n",
          "IN_WIDTH: %0d", IN_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_pad #(
    parameter IN_WIDTH  = 32,
    parameter OUT_WIDTH = 32
) (
   input wire logic [IN_WIDTH-1:0]  in,
   output logic     [OUT_WIDTH-1:0] out
);
  localparam EXTEND = OUT_WIDTH - IN_WIDTH;
  assign out = { {EXTEND {1'b0}}, in};

  `ifdef VERILATOR
    always_comb begin
      if (IN_WIDTH > OUT_WIDTH)
        $error(
          "std_pad: Output width less than input width\n",
          "IN_WIDTH: %0d", IN_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_cat #(
  parameter LEFT_WIDTH  = 32,
  parameter RIGHT_WIDTH = 32,
  parameter OUT_WIDTH = 64
) (
  input wire logic [LEFT_WIDTH-1:0] left,
  input wire logic [RIGHT_WIDTH-1:0] right,
  output logic [OUT_WIDTH-1:0] out
);
  assign out = {left, right};

  `ifdef VERILATOR
    always_comb begin
      if (LEFT_WIDTH + RIGHT_WIDTH != OUT_WIDTH)
        $error(
          "std_cat: Output width must equal sum of input widths\n",
          "LEFT_WIDTH: %0d", LEFT_WIDTH,
          "RIGHT_WIDTH: %0d", RIGHT_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_not #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] in,
   output logic [WIDTH-1:0] out
);
  assign out = ~in;
endmodule

module std_and #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left & right;
endmodule

module std_or #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left | right;
endmodule

module std_xor #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left ^ right;
endmodule

module std_sub #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module std_gt #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left > right;
endmodule

module std_lt #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left < right;
endmodule

module std_eq #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left == right;
endmodule

module std_neq #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left != right;
endmodule

module std_ge #(
    parameter WIDTH = 32
) (
    input wire   logic [WIDTH-1:0] left,
    input wire   logic [WIDTH-1:0] right,
    output logic out
);
  assign out = left >= right;
endmodule

module std_le #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left <= right;
endmodule

module std_lsh #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left << right;
endmodule

module std_rsh #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left >> right;
endmodule

/// this primitive is intended to be used
/// for lowering purposes (not in source programs)
module std_mux #(
    parameter WIDTH = 32
) (
   input wire               logic cond,
   input wire               logic [WIDTH-1:0] tru,
   input wire               logic [WIDTH-1:0] fal,
   output logic [WIDTH-1:0] out
);
  assign out = cond ? tru : fal;
endmodule

module std_mem_d1 #(
    parameter WIDTH = 32,
    parameter SIZE = 16,
    parameter IDX_SIZE = 4
) (
   input wire                logic [IDX_SIZE-1:0] addr0,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  logic [WIDTH-1:0] mem[SIZE-1:0];

  /* verilator lint_off WIDTH */
  assign read_data = mem[addr0];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= SIZE)
        $error(
          "std_mem_d1: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "SIZE: %0d", SIZE
        );
    end
  `endif
endmodule

module std_mem_d2 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0];

  assign read_data = mem[addr0][addr1];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d2: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d2: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
    end
  `endif
endmodule

module std_mem_d3 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D2_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4,
    parameter D2_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [D2_IDX_SIZE-1:0] addr2,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0][D2_SIZE-1:0];

  assign read_data = mem[addr0][addr1][addr2];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1][addr2] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
      if (addr2 >= D2_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr2: %0d\n", addr2,
          "D2_SIZE: %0d", D2_SIZE
        );
    end
  `endif
endmodule

module std_mem_d4 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D2_SIZE = 16,
    parameter D3_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4,
    parameter D2_IDX_SIZE = 4,
    parameter D3_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [D2_IDX_SIZE-1:0] addr2,
   input wire                logic [D3_IDX_SIZE-1:0] addr3,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   input wire                logic reset,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0][D2_SIZE-1:0][D3_SIZE-1:0];

  assign read_data = mem[addr0][addr1][addr2][addr3];

  always_ff @(posedge clk) begin
    if (reset)
      done <= '0;
    else if (write_en)
      done <= '1;
    else
      done <= '0;
  end

  always_ff @(posedge clk) begin
    if (!reset && write_en)
      mem[addr0][addr1][addr2][addr3] <= write_data;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
      if (addr2 >= D2_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr2: %0d\n", addr2,
          "D2_SIZE: %0d", D2_SIZE
        );
      if (addr3 >= D3_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr3: %0d\n", addr3,
          "D3_SIZE: %0d", D3_SIZE
        );
    end
  `endif
endmodule

`default_nettype wire

module undef #(
    parameter WIDTH = 32
) (
   output logic [WIDTH-1:0] out
);
assign out = 'x;
endmodule

module std_const #(
    parameter WIDTH = 32,
    parameter VALUE = 32
) (
   output logic [WIDTH-1:0] out
);
assign out = VALUE;
endmodule

module std_wire #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] in,
   output logic [WIDTH-1:0] out
);
assign out = in;
endmodule

module std_add #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] left,
   input logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
assign out = left + right;
endmodule

module std_reg #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] in,
   input logic write_en,
   input logic clk,
   input logic reset,
   output logic [WIDTH-1:0] out,
   output logic done
);
always_ff @(posedge clk) begin
    if (reset) begin
       out <= 0;
       done <= 0;
    end else if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module mac_pe(
  input logic [31:0] top,
  input logic [31:0] left,
  input logic mul_ready,
  output logic [31:0] out,
  input logic go,
  input logic clk,
  input logic reset,
  output logic done
);
// COMPONENT START: mac_pe
logic [31:0] acc_in;
logic acc_write_en;
logic acc_clk;
logic acc_reset;
logic [31:0] acc_out;
logic acc_done;
logic [31:0] add_left;
logic [31:0] add_right;
logic [31:0] add_out;
logic mul_clk;
logic [31:0] mul_left;
logic [31:0] mul_right;
logic [31:0] mul_out;
logic fsm_in;
logic fsm_write_en;
logic fsm_clk;
logic fsm_reset;
logic fsm_out;
logic fsm_done;
logic ud_out;
logic adder_left;
logic adder_right;
logic adder_out;
logic signal_reg_in;
logic signal_reg_write_en;
logic signal_reg_clk;
logic signal_reg_reset;
logic signal_reg_out;
logic signal_reg_done;
logic early_reset_static_par_go_in;
logic early_reset_static_par_go_out;
logic early_reset_static_par_done_in;
logic early_reset_static_par_done_out;
logic wrapper_early_reset_static_par_go_in;
logic wrapper_early_reset_static_par_go_out;
logic wrapper_early_reset_static_par_done_in;
logic wrapper_early_reset_static_par_done_out;
std_reg # (
    .WIDTH(32)
) acc (
    .clk(acc_clk),
    .done(acc_done),
    .in(acc_in),
    .out(acc_out),
    .reset(acc_reset),
    .write_en(acc_write_en)
);
std_add # (
    .WIDTH(32)
) add (
    .left(add_left),
    .out(add_out),
    .right(add_right)
);
bb_pipelined_mult mul (
    .clk(mul_clk),
    .left(mul_left),
    .out(mul_out),
    .right(mul_right)
);
std_reg # (
    .WIDTH(1)
) fsm (
    .clk(fsm_clk),
    .done(fsm_done),
    .in(fsm_in),
    .out(fsm_out),
    .reset(fsm_reset),
    .write_en(fsm_write_en)
);
undef # (
    .WIDTH(1)
) ud (
    .out(ud_out)
);
std_add # (
    .WIDTH(1)
) adder (
    .left(adder_left),
    .out(adder_out),
    .right(adder_right)
);
std_reg # (
    .WIDTH(1)
) signal_reg (
    .clk(signal_reg_clk),
    .done(signal_reg_done),
    .in(signal_reg_in),
    .out(signal_reg_out),
    .reset(signal_reg_reset),
    .write_en(signal_reg_write_en)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_go (
    .in(early_reset_static_par_go_in),
    .out(early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par_done (
    .in(early_reset_static_par_done_in),
    .out(early_reset_static_par_done_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_go (
    .in(wrapper_early_reset_static_par_go_in),
    .out(wrapper_early_reset_static_par_go_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_par_done (
    .in(wrapper_early_reset_static_par_done_in),
    .out(wrapper_early_reset_static_par_done_out)
);
wire _guard0 = 1;
wire _guard1 = early_reset_static_par_go_out;
wire _guard2 = early_reset_static_par_go_out;
wire _guard3 = wrapper_early_reset_static_par_done_out;
wire _guard4 = early_reset_static_par_go_out;
wire _guard5 = fsm_out != 1'd0;
wire _guard6 = early_reset_static_par_go_out;
wire _guard7 = _guard5 & _guard6;
wire _guard8 = fsm_out == 1'd0;
wire _guard9 = early_reset_static_par_go_out;
wire _guard10 = _guard8 & _guard9;
wire _guard11 = early_reset_static_par_go_out;
wire _guard12 = early_reset_static_par_go_out;
wire _guard13 = fsm_out == 1'd0;
wire _guard14 = signal_reg_out;
wire _guard15 = _guard13 & _guard14;
wire _guard16 = fsm_out == 1'd0;
wire _guard17 = signal_reg_out;
wire _guard18 = _guard16 & _guard17;
wire _guard19 = fsm_out == 1'd0;
wire _guard20 = signal_reg_out;
wire _guard21 = ~_guard20;
wire _guard22 = _guard19 & _guard21;
wire _guard23 = wrapper_early_reset_static_par_go_out;
wire _guard24 = _guard22 & _guard23;
wire _guard25 = _guard18 | _guard24;
wire _guard26 = fsm_out == 1'd0;
wire _guard27 = signal_reg_out;
wire _guard28 = ~_guard27;
wire _guard29 = _guard26 & _guard28;
wire _guard30 = wrapper_early_reset_static_par_go_out;
wire _guard31 = _guard29 & _guard30;
wire _guard32 = fsm_out == 1'd0;
wire _guard33 = signal_reg_out;
wire _guard34 = _guard32 & _guard33;
wire _guard35 = early_reset_static_par_go_out;
wire _guard36 = early_reset_static_par_go_out;
wire _guard37 = early_reset_static_par_go_out;
wire _guard38 = early_reset_static_par_go_out;
wire _guard39 = wrapper_early_reset_static_par_go_out;
assign acc_write_en =
  _guard1 ? mul_ready :
  1'd0;
assign acc_clk = clk;
assign acc_reset = reset;
assign acc_in = add_out;
assign done = _guard3;
assign out = acc_out;
assign fsm_write_en = _guard4;
assign fsm_clk = clk;
assign fsm_reset = reset;
assign fsm_in =
  _guard7 ? adder_out :
  _guard10 ? 1'd0 :
  1'd0;
assign adder_left =
  _guard11 ? fsm_out :
  1'd0;
assign adder_right = _guard12;
assign wrapper_early_reset_static_par_go_in = go;
assign wrapper_early_reset_static_par_done_in = _guard15;
assign early_reset_static_par_done_in = ud_out;
assign signal_reg_write_en = _guard25;
assign signal_reg_clk = clk;
assign signal_reg_reset = reset;
assign signal_reg_in =
  _guard31 ? 1'd1 :
  _guard34 ? 1'd0 :
  1'd0;
assign add_left = acc_out;
assign add_right = mul_out;
assign mul_clk = clk;
assign mul_left =
  _guard37 ? top :
  32'd0;
assign mul_right =
  _guard38 ? left :
  32'd0;
assign early_reset_static_par_go_in = _guard39;
// COMPONENT END: mac_pe
endmodule
module main(
  input logic go,
  input logic clk,
  input logic reset,
  output logic done,
  output logic [2:0] t0_addr0,
  output logic [31:0] t0_write_data,
  output logic t0_write_en,
  output logic t0_clk,
  output logic t0_reset,
  input logic [31:0] t0_read_data,
  input logic t0_done,
  output logic [2:0] t1_addr0,
  output logic [31:0] t1_write_data,
  output logic t1_write_en,
  output logic t1_clk,
  output logic t1_reset,
  input logic [31:0] t1_read_data,
  input logic t1_done,
  output logic [2:0] t2_addr0,
  output logic [31:0] t2_write_data,
  output logic t2_write_en,
  output logic t2_clk,
  output logic t2_reset,
  input logic [31:0] t2_read_data,
  input logic t2_done,
  output logic [2:0] t3_addr0,
  output logic [31:0] t3_write_data,
  output logic t3_write_en,
  output logic t3_clk,
  output logic t3_reset,
  input logic [31:0] t3_read_data,
  input logic t3_done,
  output logic [2:0] l0_addr0,
  output logic [31:0] l0_write_data,
  output logic l0_write_en,
  output logic l0_clk,
  output logic l0_reset,
  input logic [31:0] l0_read_data,
  input logic l0_done,
  output logic [2:0] l1_addr0,
  output logic [31:0] l1_write_data,
  output logic l1_write_en,
  output logic l1_clk,
  output logic l1_reset,
  input logic [31:0] l1_read_data,
  input logic l1_done,
  output logic [2:0] l2_addr0,
  output logic [31:0] l2_write_data,
  output logic l2_write_en,
  output logic l2_clk,
  output logic l2_reset,
  input logic [31:0] l2_read_data,
  input logic l2_done,
  output logic [2:0] l3_addr0,
  output logic [31:0] l3_write_data,
  output logic l3_write_en,
  output logic l3_clk,
  output logic l3_reset,
  input logic [31:0] l3_read_data,
  input logic l3_done,
  output logic [2:0] out_mem_0_addr0,
  output logic [31:0] out_mem_0_write_data,
  output logic out_mem_0_write_en,
  output logic out_mem_0_clk,
  output logic out_mem_0_reset,
  input logic [31:0] out_mem_0_read_data,
  input logic out_mem_0_done,
  output logic [2:0] out_mem_1_addr0,
  output logic [31:0] out_mem_1_write_data,
  output logic out_mem_1_write_en,
  output logic out_mem_1_clk,
  output logic out_mem_1_reset,
  input logic [31:0] out_mem_1_read_data,
  input logic out_mem_1_done,
  output logic [2:0] out_mem_2_addr0,
  output logic [31:0] out_mem_2_write_data,
  output logic out_mem_2_write_en,
  output logic out_mem_2_clk,
  output logic out_mem_2_reset,
  input logic [31:0] out_mem_2_read_data,
  input logic out_mem_2_done,
  output logic [2:0] out_mem_3_addr0,
  output logic [31:0] out_mem_3_write_data,
  output logic out_mem_3_write_en,
  output logic out_mem_3_clk,
  output logic out_mem_3_reset,
  input logic [31:0] out_mem_3_read_data,
  input logic out_mem_3_done
);
// COMPONENT START: main
logic [31:0] pe_0_0_top;
logic [31:0] pe_0_0_left;
logic pe_0_0_mul_ready;
logic [31:0] pe_0_0_out;
logic pe_0_0_go;
logic pe_0_0_clk;
logic pe_0_0_reset;
logic pe_0_0_done;
logic [31:0] top_0_0_in;
logic top_0_0_write_en;
logic top_0_0_clk;
logic top_0_0_reset;
logic [31:0] top_0_0_out;
logic top_0_0_done;
logic [31:0] left_0_0_in;
logic left_0_0_write_en;
logic left_0_0_clk;
logic left_0_0_reset;
logic [31:0] left_0_0_out;
logic left_0_0_done;
logic [31:0] pe_0_1_top;
logic [31:0] pe_0_1_left;
logic pe_0_1_mul_ready;
logic [31:0] pe_0_1_out;
logic pe_0_1_go;
logic pe_0_1_clk;
logic pe_0_1_reset;
logic pe_0_1_done;
logic [31:0] top_0_1_in;
logic top_0_1_write_en;
logic top_0_1_clk;
logic top_0_1_reset;
logic [31:0] top_0_1_out;
logic top_0_1_done;
logic [31:0] left_0_1_in;
logic left_0_1_write_en;
logic left_0_1_clk;
logic left_0_1_reset;
logic [31:0] left_0_1_out;
logic left_0_1_done;
logic [31:0] pe_0_2_top;
logic [31:0] pe_0_2_left;
logic pe_0_2_mul_ready;
logic [31:0] pe_0_2_out;
logic pe_0_2_go;
logic pe_0_2_clk;
logic pe_0_2_reset;
logic pe_0_2_done;
logic [31:0] top_0_2_in;
logic top_0_2_write_en;
logic top_0_2_clk;
logic top_0_2_reset;
logic [31:0] top_0_2_out;
logic top_0_2_done;
logic [31:0] left_0_2_in;
logic left_0_2_write_en;
logic left_0_2_clk;
logic left_0_2_reset;
logic [31:0] left_0_2_out;
logic left_0_2_done;
logic [31:0] pe_0_3_top;
logic [31:0] pe_0_3_left;
logic pe_0_3_mul_ready;
logic [31:0] pe_0_3_out;
logic pe_0_3_go;
logic pe_0_3_clk;
logic pe_0_3_reset;
logic pe_0_3_done;
logic [31:0] top_0_3_in;
logic top_0_3_write_en;
logic top_0_3_clk;
logic top_0_3_reset;
logic [31:0] top_0_3_out;
logic top_0_3_done;
logic [31:0] left_0_3_in;
logic left_0_3_write_en;
logic left_0_3_clk;
logic left_0_3_reset;
logic [31:0] left_0_3_out;
logic left_0_3_done;
logic [31:0] pe_1_0_top;
logic [31:0] pe_1_0_left;
logic pe_1_0_mul_ready;
logic [31:0] pe_1_0_out;
logic pe_1_0_go;
logic pe_1_0_clk;
logic pe_1_0_reset;
logic pe_1_0_done;
logic [31:0] top_1_0_in;
logic top_1_0_write_en;
logic top_1_0_clk;
logic top_1_0_reset;
logic [31:0] top_1_0_out;
logic top_1_0_done;
logic [31:0] left_1_0_in;
logic left_1_0_write_en;
logic left_1_0_clk;
logic left_1_0_reset;
logic [31:0] left_1_0_out;
logic left_1_0_done;
logic [31:0] pe_1_1_top;
logic [31:0] pe_1_1_left;
logic pe_1_1_mul_ready;
logic [31:0] pe_1_1_out;
logic pe_1_1_go;
logic pe_1_1_clk;
logic pe_1_1_reset;
logic pe_1_1_done;
logic [31:0] top_1_1_in;
logic top_1_1_write_en;
logic top_1_1_clk;
logic top_1_1_reset;
logic [31:0] top_1_1_out;
logic top_1_1_done;
logic [31:0] left_1_1_in;
logic left_1_1_write_en;
logic left_1_1_clk;
logic left_1_1_reset;
logic [31:0] left_1_1_out;
logic left_1_1_done;
logic [31:0] pe_1_2_top;
logic [31:0] pe_1_2_left;
logic pe_1_2_mul_ready;
logic [31:0] pe_1_2_out;
logic pe_1_2_go;
logic pe_1_2_clk;
logic pe_1_2_reset;
logic pe_1_2_done;
logic [31:0] top_1_2_in;
logic top_1_2_write_en;
logic top_1_2_clk;
logic top_1_2_reset;
logic [31:0] top_1_2_out;
logic top_1_2_done;
logic [31:0] left_1_2_in;
logic left_1_2_write_en;
logic left_1_2_clk;
logic left_1_2_reset;
logic [31:0] left_1_2_out;
logic left_1_2_done;
logic [31:0] pe_1_3_top;
logic [31:0] pe_1_3_left;
logic pe_1_3_mul_ready;
logic [31:0] pe_1_3_out;
logic pe_1_3_go;
logic pe_1_3_clk;
logic pe_1_3_reset;
logic pe_1_3_done;
logic [31:0] top_1_3_in;
logic top_1_3_write_en;
logic top_1_3_clk;
logic top_1_3_reset;
logic [31:0] top_1_3_out;
logic top_1_3_done;
logic [31:0] left_1_3_in;
logic left_1_3_write_en;
logic left_1_3_clk;
logic left_1_3_reset;
logic [31:0] left_1_3_out;
logic left_1_3_done;
logic [31:0] pe_2_0_top;
logic [31:0] pe_2_0_left;
logic pe_2_0_mul_ready;
logic [31:0] pe_2_0_out;
logic pe_2_0_go;
logic pe_2_0_clk;
logic pe_2_0_reset;
logic pe_2_0_done;
logic [31:0] top_2_0_in;
logic top_2_0_write_en;
logic top_2_0_clk;
logic top_2_0_reset;
logic [31:0] top_2_0_out;
logic top_2_0_done;
logic [31:0] left_2_0_in;
logic left_2_0_write_en;
logic left_2_0_clk;
logic left_2_0_reset;
logic [31:0] left_2_0_out;
logic left_2_0_done;
logic [31:0] pe_2_1_top;
logic [31:0] pe_2_1_left;
logic pe_2_1_mul_ready;
logic [31:0] pe_2_1_out;
logic pe_2_1_go;
logic pe_2_1_clk;
logic pe_2_1_reset;
logic pe_2_1_done;
logic [31:0] top_2_1_in;
logic top_2_1_write_en;
logic top_2_1_clk;
logic top_2_1_reset;
logic [31:0] top_2_1_out;
logic top_2_1_done;
logic [31:0] left_2_1_in;
logic left_2_1_write_en;
logic left_2_1_clk;
logic left_2_1_reset;
logic [31:0] left_2_1_out;
logic left_2_1_done;
logic [31:0] pe_2_2_top;
logic [31:0] pe_2_2_left;
logic pe_2_2_mul_ready;
logic [31:0] pe_2_2_out;
logic pe_2_2_go;
logic pe_2_2_clk;
logic pe_2_2_reset;
logic pe_2_2_done;
logic [31:0] top_2_2_in;
logic top_2_2_write_en;
logic top_2_2_clk;
logic top_2_2_reset;
logic [31:0] top_2_2_out;
logic top_2_2_done;
logic [31:0] left_2_2_in;
logic left_2_2_write_en;
logic left_2_2_clk;
logic left_2_2_reset;
logic [31:0] left_2_2_out;
logic left_2_2_done;
logic [31:0] pe_2_3_top;
logic [31:0] pe_2_3_left;
logic pe_2_3_mul_ready;
logic [31:0] pe_2_3_out;
logic pe_2_3_go;
logic pe_2_3_clk;
logic pe_2_3_reset;
logic pe_2_3_done;
logic [31:0] top_2_3_in;
logic top_2_3_write_en;
logic top_2_3_clk;
logic top_2_3_reset;
logic [31:0] top_2_3_out;
logic top_2_3_done;
logic [31:0] left_2_3_in;
logic left_2_3_write_en;
logic left_2_3_clk;
logic left_2_3_reset;
logic [31:0] left_2_3_out;
logic left_2_3_done;
logic [31:0] pe_3_0_top;
logic [31:0] pe_3_0_left;
logic pe_3_0_mul_ready;
logic [31:0] pe_3_0_out;
logic pe_3_0_go;
logic pe_3_0_clk;
logic pe_3_0_reset;
logic pe_3_0_done;
logic [31:0] top_3_0_in;
logic top_3_0_write_en;
logic top_3_0_clk;
logic top_3_0_reset;
logic [31:0] top_3_0_out;
logic top_3_0_done;
logic [31:0] left_3_0_in;
logic left_3_0_write_en;
logic left_3_0_clk;
logic left_3_0_reset;
logic [31:0] left_3_0_out;
logic left_3_0_done;
logic [31:0] pe_3_1_top;
logic [31:0] pe_3_1_left;
logic pe_3_1_mul_ready;
logic [31:0] pe_3_1_out;
logic pe_3_1_go;
logic pe_3_1_clk;
logic pe_3_1_reset;
logic pe_3_1_done;
logic [31:0] top_3_1_in;
logic top_3_1_write_en;
logic top_3_1_clk;
logic top_3_1_reset;
logic [31:0] top_3_1_out;
logic top_3_1_done;
logic [31:0] left_3_1_in;
logic left_3_1_write_en;
logic left_3_1_clk;
logic left_3_1_reset;
logic [31:0] left_3_1_out;
logic left_3_1_done;
logic [31:0] pe_3_2_top;
logic [31:0] pe_3_2_left;
logic pe_3_2_mul_ready;
logic [31:0] pe_3_2_out;
logic pe_3_2_go;
logic pe_3_2_clk;
logic pe_3_2_reset;
logic pe_3_2_done;
logic [31:0] top_3_2_in;
logic top_3_2_write_en;
logic top_3_2_clk;
logic top_3_2_reset;
logic [31:0] top_3_2_out;
logic top_3_2_done;
logic [31:0] left_3_2_in;
logic left_3_2_write_en;
logic left_3_2_clk;
logic left_3_2_reset;
logic [31:0] left_3_2_out;
logic left_3_2_done;
logic [31:0] pe_3_3_top;
logic [31:0] pe_3_3_left;
logic pe_3_3_mul_ready;
logic [31:0] pe_3_3_out;
logic pe_3_3_go;
logic pe_3_3_clk;
logic pe_3_3_reset;
logic pe_3_3_done;
logic [31:0] top_3_3_in;
logic top_3_3_write_en;
logic top_3_3_clk;
logic top_3_3_reset;
logic [31:0] top_3_3_out;
logic top_3_3_done;
logic [31:0] left_3_3_in;
logic left_3_3_write_en;
logic left_3_3_clk;
logic left_3_3_reset;
logic [31:0] left_3_3_out;
logic left_3_3_done;
logic [2:0] t0_idx_in;
logic t0_idx_write_en;
logic t0_idx_clk;
logic t0_idx_reset;
logic [2:0] t0_idx_out;
logic t0_idx_done;
logic [2:0] t0_add_left;
logic [2:0] t0_add_right;
logic [2:0] t0_add_out;
logic [2:0] t1_idx_in;
logic t1_idx_write_en;
logic t1_idx_clk;
logic t1_idx_reset;
logic [2:0] t1_idx_out;
logic t1_idx_done;
logic [2:0] t1_add_left;
logic [2:0] t1_add_right;
logic [2:0] t1_add_out;
logic [2:0] t2_idx_in;
logic t2_idx_write_en;
logic t2_idx_clk;
logic t2_idx_reset;
logic [2:0] t2_idx_out;
logic t2_idx_done;
logic [2:0] t2_add_left;
logic [2:0] t2_add_right;
logic [2:0] t2_add_out;
logic [2:0] t3_idx_in;
logic t3_idx_write_en;
logic t3_idx_clk;
logic t3_idx_reset;
logic [2:0] t3_idx_out;
logic t3_idx_done;
logic [2:0] t3_add_left;
logic [2:0] t3_add_right;
logic [2:0] t3_add_out;
logic [2:0] l0_idx_in;
logic l0_idx_write_en;
logic l0_idx_clk;
logic l0_idx_reset;
logic [2:0] l0_idx_out;
logic l0_idx_done;
logic [2:0] l0_add_left;
logic [2:0] l0_add_right;
logic [2:0] l0_add_out;
logic [2:0] l1_idx_in;
logic l1_idx_write_en;
logic l1_idx_clk;
logic l1_idx_reset;
logic [2:0] l1_idx_out;
logic l1_idx_done;
logic [2:0] l1_add_left;
logic [2:0] l1_add_right;
logic [2:0] l1_add_out;
logic [2:0] l2_idx_in;
logic l2_idx_write_en;
logic l2_idx_clk;
logic l2_idx_reset;
logic [2:0] l2_idx_out;
logic l2_idx_done;
logic [2:0] l2_add_left;
logic [2:0] l2_add_right;
logic [2:0] l2_add_out;
logic [2:0] l3_idx_in;
logic l3_idx_write_en;
logic l3_idx_clk;
logic l3_idx_reset;
logic [2:0] l3_idx_out;
logic l3_idx_done;
logic [2:0] l3_add_left;
logic [2:0] l3_add_right;
logic [2:0] l3_add_out;
logic [4:0] idx_in;
logic idx_write_en;
logic idx_clk;
logic idx_reset;
logic [4:0] idx_out;
logic idx_done;
logic [4:0] idx_add_left;
logic [4:0] idx_add_right;
logic [4:0] idx_add_out;
logic idx_between_3_7_reg_in;
logic idx_between_3_7_reg_write_en;
logic idx_between_3_7_reg_clk;
logic idx_between_3_7_reg_reset;
logic idx_between_3_7_reg_out;
logic idx_between_3_7_reg_done;
logic [4:0] index_lt_7_left;
logic [4:0] index_lt_7_right;
logic index_lt_7_out;
logic [4:0] index_ge_3_left;
logic [4:0] index_ge_3_right;
logic index_ge_3_out;
logic idx_between_3_7_comb_left;
logic idx_between_3_7_comb_right;
logic idx_between_3_7_comb_out;
logic idx_between_12_13_reg_in;
logic idx_between_12_13_reg_write_en;
logic idx_between_12_13_reg_clk;
logic idx_between_12_13_reg_reset;
logic idx_between_12_13_reg_out;
logic idx_between_12_13_reg_done;
logic [4:0] index_lt_13_left;
logic [4:0] index_lt_13_right;
logic index_lt_13_out;
logic [4:0] index_ge_12_left;
logic [4:0] index_ge_12_right;
logic index_ge_12_out;
logic idx_between_12_13_comb_left;
logic idx_between_12_13_comb_right;
logic idx_between_12_13_comb_out;
logic idx_between_8_12_reg_in;
logic idx_between_8_12_reg_write_en;
logic idx_between_8_12_reg_clk;
logic idx_between_8_12_reg_reset;
logic idx_between_8_12_reg_out;
logic idx_between_8_12_reg_done;
logic [4:0] index_lt_12_left;
logic [4:0] index_lt_12_right;
logic index_lt_12_out;
logic [4:0] index_ge_8_left;
logic [4:0] index_ge_8_right;
logic index_ge_8_out;
logic idx_between_8_12_comb_left;
logic idx_between_8_12_comb_right;
logic idx_between_8_12_comb_out;
logic idx_between_13_14_reg_in;
logic idx_between_13_14_reg_write_en;
logic idx_between_13_14_reg_clk;
logic idx_between_13_14_reg_reset;
logic idx_between_13_14_reg_out;
logic idx_between_13_14_reg_done;
logic [4:0] index_lt_14_left;
logic [4:0] index_lt_14_right;
logic index_lt_14_out;
logic [4:0] index_ge_13_left;
logic [4:0] index_ge_13_right;
logic index_ge_13_out;
logic idx_between_13_14_comb_left;
logic idx_between_13_14_comb_right;
logic idx_between_13_14_comb_out;
logic idx_between_4_8_reg_in;
logic idx_between_4_8_reg_write_en;
logic idx_between_4_8_reg_clk;
logic idx_between_4_8_reg_reset;
logic idx_between_4_8_reg_out;
logic idx_between_4_8_reg_done;
logic [4:0] index_lt_8_left;
logic [4:0] index_lt_8_right;
logic index_lt_8_out;
logic [4:0] index_ge_4_left;
logic [4:0] index_ge_4_right;
logic index_ge_4_out;
logic idx_between_4_8_comb_left;
logic idx_between_4_8_comb_right;
logic idx_between_4_8_comb_out;
logic idx_between_5_9_reg_in;
logic idx_between_5_9_reg_write_en;
logic idx_between_5_9_reg_clk;
logic idx_between_5_9_reg_reset;
logic idx_between_5_9_reg_out;
logic idx_between_5_9_reg_done;
logic [4:0] index_lt_9_left;
logic [4:0] index_lt_9_right;
logic index_lt_9_out;
logic [4:0] index_ge_5_left;
logic [4:0] index_ge_5_right;
logic index_ge_5_out;
logic idx_between_5_9_comb_left;
logic idx_between_5_9_comb_right;
logic idx_between_5_9_comb_out;
logic idx_between_14_15_reg_in;
logic idx_between_14_15_reg_write_en;
logic idx_between_14_15_reg_clk;
logic idx_between_14_15_reg_reset;
logic idx_between_14_15_reg_out;
logic idx_between_14_15_reg_done;
logic [4:0] index_lt_15_left;
logic [4:0] index_lt_15_right;
logic index_lt_15_out;
logic [4:0] index_ge_14_left;
logic [4:0] index_ge_14_right;
logic index_ge_14_out;
logic idx_between_14_15_comb_left;
logic idx_between_14_15_comb_right;
logic idx_between_14_15_comb_out;
logic idx_between_9_10_reg_in;
logic idx_between_9_10_reg_write_en;
logic idx_between_9_10_reg_clk;
logic idx_between_9_10_reg_reset;
logic idx_between_9_10_reg_out;
logic idx_between_9_10_reg_done;
logic [4:0] index_lt_10_left;
logic [4:0] index_lt_10_right;
logic index_lt_10_out;
logic [4:0] index_ge_9_left;
logic [4:0] index_ge_9_right;
logic index_ge_9_out;
logic idx_between_9_10_comb_left;
logic idx_between_9_10_comb_right;
logic idx_between_9_10_comb_out;
logic idx_between_10_11_reg_in;
logic idx_between_10_11_reg_write_en;
logic idx_between_10_11_reg_clk;
logic idx_between_10_11_reg_reset;
logic idx_between_10_11_reg_out;
logic idx_between_10_11_reg_done;
logic [4:0] index_lt_11_left;
logic [4:0] index_lt_11_right;
logic index_lt_11_out;
logic [4:0] index_ge_10_left;
logic [4:0] index_ge_10_right;
logic index_ge_10_out;
logic idx_between_10_11_comb_left;
logic idx_between_10_11_comb_right;
logic idx_between_10_11_comb_out;
logic idx_between_0_4_reg_in;
logic idx_between_0_4_reg_write_en;
logic idx_between_0_4_reg_clk;
logic idx_between_0_4_reg_reset;
logic idx_between_0_4_reg_out;
logic idx_between_0_4_reg_done;
logic [4:0] index_lt_4_left;
logic [4:0] index_lt_4_right;
logic index_lt_4_out;
logic idx_between_9_13_reg_in;
logic idx_between_9_13_reg_write_en;
logic idx_between_9_13_reg_clk;
logic idx_between_9_13_reg_reset;
logic idx_between_9_13_reg_out;
logic idx_between_9_13_reg_done;
logic idx_between_9_13_comb_left;
logic idx_between_9_13_comb_right;
logic idx_between_9_13_comb_out;
logic idx_between_1_5_reg_in;
logic idx_between_1_5_reg_write_en;
logic idx_between_1_5_reg_clk;
logic idx_between_1_5_reg_reset;
logic idx_between_1_5_reg_out;
logic idx_between_1_5_reg_done;
logic [4:0] index_lt_5_left;
logic [4:0] index_lt_5_right;
logic index_lt_5_out;
logic [4:0] index_ge_1_left;
logic [4:0] index_ge_1_right;
logic index_ge_1_out;
logic idx_between_1_5_comb_left;
logic idx_between_1_5_comb_right;
logic idx_between_1_5_comb_out;
logic idx_between_10_14_reg_in;
logic idx_between_10_14_reg_write_en;
logic idx_between_10_14_reg_clk;
logic idx_between_10_14_reg_reset;
logic idx_between_10_14_reg_out;
logic idx_between_10_14_reg_done;
logic idx_between_10_14_comb_left;
logic idx_between_10_14_comb_right;
logic idx_between_10_14_comb_out;
logic idx_between_15_16_reg_in;
logic idx_between_15_16_reg_write_en;
logic idx_between_15_16_reg_clk;
logic idx_between_15_16_reg_reset;
logic idx_between_15_16_reg_out;
logic idx_between_15_16_reg_done;
logic [4:0] index_lt_16_left;
logic [4:0] index_lt_16_right;
logic index_lt_16_out;
logic [4:0] index_ge_15_left;
logic [4:0] index_ge_15_right;
logic index_ge_15_out;
logic idx_between_15_16_comb_left;
logic idx_between_15_16_comb_right;
logic idx_between_15_16_comb_out;
logic idx_between_6_10_reg_in;
logic idx_between_6_10_reg_write_en;
logic idx_between_6_10_reg_clk;
logic idx_between_6_10_reg_reset;
logic idx_between_6_10_reg_out;
logic idx_between_6_10_reg_done;
logic [4:0] index_ge_6_left;
logic [4:0] index_ge_6_right;
logic index_ge_6_out;
logic idx_between_6_10_comb_left;
logic idx_between_6_10_comb_right;
logic idx_between_6_10_comb_out;
logic idx_between_11_12_reg_in;
logic idx_between_11_12_reg_write_en;
logic idx_between_11_12_reg_clk;
logic idx_between_11_12_reg_reset;
logic idx_between_11_12_reg_out;
logic idx_between_11_12_reg_done;
logic [4:0] index_ge_11_left;
logic [4:0] index_ge_11_right;
logic index_ge_11_out;
logic idx_between_11_12_comb_left;
logic idx_between_11_12_comb_right;
logic idx_between_11_12_comb_out;
logic idx_between_2_6_reg_in;
logic idx_between_2_6_reg_write_en;
logic idx_between_2_6_reg_clk;
logic idx_between_2_6_reg_reset;
logic idx_between_2_6_reg_out;
logic idx_between_2_6_reg_done;
logic [4:0] index_lt_6_left;
logic [4:0] index_lt_6_right;
logic index_lt_6_out;
logic [4:0] index_ge_2_left;
logic [4:0] index_ge_2_right;
logic index_ge_2_out;
logic idx_between_2_6_comb_left;
logic idx_between_2_6_comb_right;
logic idx_between_2_6_comb_out;
logic idx_between_11_15_reg_in;
logic idx_between_11_15_reg_write_en;
logic idx_between_11_15_reg_clk;
logic idx_between_11_15_reg_reset;
logic idx_between_11_15_reg_out;
logic idx_between_11_15_reg_done;
logic idx_between_11_15_comb_left;
logic idx_between_11_15_comb_right;
logic idx_between_11_15_comb_out;
logic idx_between_7_11_reg_in;
logic idx_between_7_11_reg_write_en;
logic idx_between_7_11_reg_clk;
logic idx_between_7_11_reg_reset;
logic idx_between_7_11_reg_out;
logic idx_between_7_11_reg_done;
logic [4:0] index_ge_7_left;
logic [4:0] index_ge_7_right;
logic index_ge_7_out;
logic idx_between_7_11_comb_left;
logic idx_between_7_11_comb_right;
logic idx_between_7_11_comb_out;
logic cond_in;
logic cond_write_en;
logic cond_clk;
logic cond_reset;
logic cond_out;
logic cond_done;
logic cond_wire_in;
logic cond_wire_out;
logic cond0_in;
logic cond0_write_en;
logic cond0_clk;
logic cond0_reset;
logic cond0_out;
logic cond0_done;
logic cond_wire0_in;
logic cond_wire0_out;
logic cond1_in;
logic cond1_write_en;
logic cond1_clk;
logic cond1_reset;
logic cond1_out;
logic cond1_done;
logic cond_wire1_in;
logic cond_wire1_out;
logic cond2_in;
logic cond2_write_en;
logic cond2_clk;
logic cond2_reset;
logic cond2_out;
logic cond2_done;
logic cond_wire2_in;
logic cond_wire2_out;
logic cond3_in;
logic cond3_write_en;
logic cond3_clk;
logic cond3_reset;
logic cond3_out;
logic cond3_done;
logic cond_wire3_in;
logic cond_wire3_out;
logic cond4_in;
logic cond4_write_en;
logic cond4_clk;
logic cond4_reset;
logic cond4_out;
logic cond4_done;
logic cond_wire4_in;
logic cond_wire4_out;
logic cond5_in;
logic cond5_write_en;
logic cond5_clk;
logic cond5_reset;
logic cond5_out;
logic cond5_done;
logic cond_wire5_in;
logic cond_wire5_out;
logic cond6_in;
logic cond6_write_en;
logic cond6_clk;
logic cond6_reset;
logic cond6_out;
logic cond6_done;
logic cond_wire6_in;
logic cond_wire6_out;
logic cond7_in;
logic cond7_write_en;
logic cond7_clk;
logic cond7_reset;
logic cond7_out;
logic cond7_done;
logic cond_wire7_in;
logic cond_wire7_out;
logic cond8_in;
logic cond8_write_en;
logic cond8_clk;
logic cond8_reset;
logic cond8_out;
logic cond8_done;
logic cond_wire8_in;
logic cond_wire8_out;
logic cond9_in;
logic cond9_write_en;
logic cond9_clk;
logic cond9_reset;
logic cond9_out;
logic cond9_done;
logic cond_wire9_in;
logic cond_wire9_out;
logic cond10_in;
logic cond10_write_en;
logic cond10_clk;
logic cond10_reset;
logic cond10_out;
logic cond10_done;
logic cond_wire10_in;
logic cond_wire10_out;
logic cond11_in;
logic cond11_write_en;
logic cond11_clk;
logic cond11_reset;
logic cond11_out;
logic cond11_done;
logic cond_wire11_in;
logic cond_wire11_out;
logic cond12_in;
logic cond12_write_en;
logic cond12_clk;
logic cond12_reset;
logic cond12_out;
logic cond12_done;
logic cond_wire12_in;
logic cond_wire12_out;
logic cond13_in;
logic cond13_write_en;
logic cond13_clk;
logic cond13_reset;
logic cond13_out;
logic cond13_done;
logic cond_wire13_in;
logic cond_wire13_out;
logic cond14_in;
logic cond14_write_en;
logic cond14_clk;
logic cond14_reset;
logic cond14_out;
logic cond14_done;
logic cond_wire14_in;
logic cond_wire14_out;
logic cond15_in;
logic cond15_write_en;
logic cond15_clk;
logic cond15_reset;
logic cond15_out;
logic cond15_done;
logic cond_wire15_in;
logic cond_wire15_out;
logic cond16_in;
logic cond16_write_en;
logic cond16_clk;
logic cond16_reset;
logic cond16_out;
logic cond16_done;
logic cond_wire16_in;
logic cond_wire16_out;
logic cond17_in;
logic cond17_write_en;
logic cond17_clk;
logic cond17_reset;
logic cond17_out;
logic cond17_done;
logic cond_wire17_in;
logic cond_wire17_out;
logic cond18_in;
logic cond18_write_en;
logic cond18_clk;
logic cond18_reset;
logic cond18_out;
logic cond18_done;
logic cond_wire18_in;
logic cond_wire18_out;
logic cond19_in;
logic cond19_write_en;
logic cond19_clk;
logic cond19_reset;
logic cond19_out;
logic cond19_done;
logic cond_wire19_in;
logic cond_wire19_out;
logic cond20_in;
logic cond20_write_en;
logic cond20_clk;
logic cond20_reset;
logic cond20_out;
logic cond20_done;
logic cond_wire20_in;
logic cond_wire20_out;
logic cond21_in;
logic cond21_write_en;
logic cond21_clk;
logic cond21_reset;
logic cond21_out;
logic cond21_done;
logic cond_wire21_in;
logic cond_wire21_out;
logic cond22_in;
logic cond22_write_en;
logic cond22_clk;
logic cond22_reset;
logic cond22_out;
logic cond22_done;
logic cond_wire22_in;
logic cond_wire22_out;
logic cond23_in;
logic cond23_write_en;
logic cond23_clk;
logic cond23_reset;
logic cond23_out;
logic cond23_done;
logic cond_wire23_in;
logic cond_wire23_out;
logic cond24_in;
logic cond24_write_en;
logic cond24_clk;
logic cond24_reset;
logic cond24_out;
logic cond24_done;
logic cond_wire24_in;
logic cond_wire24_out;
logic cond25_in;
logic cond25_write_en;
logic cond25_clk;
logic cond25_reset;
logic cond25_out;
logic cond25_done;
logic cond_wire25_in;
logic cond_wire25_out;
logic cond26_in;
logic cond26_write_en;
logic cond26_clk;
logic cond26_reset;
logic cond26_out;
logic cond26_done;
logic cond_wire26_in;
logic cond_wire26_out;
logic cond27_in;
logic cond27_write_en;
logic cond27_clk;
logic cond27_reset;
logic cond27_out;
logic cond27_done;
logic cond_wire27_in;
logic cond_wire27_out;
logic cond28_in;
logic cond28_write_en;
logic cond28_clk;
logic cond28_reset;
logic cond28_out;
logic cond28_done;
logic cond_wire28_in;
logic cond_wire28_out;
logic cond29_in;
logic cond29_write_en;
logic cond29_clk;
logic cond29_reset;
logic cond29_out;
logic cond29_done;
logic cond_wire29_in;
logic cond_wire29_out;
logic cond30_in;
logic cond30_write_en;
logic cond30_clk;
logic cond30_reset;
logic cond30_out;
logic cond30_done;
logic cond_wire30_in;
logic cond_wire30_out;
logic cond31_in;
logic cond31_write_en;
logic cond31_clk;
logic cond31_reset;
logic cond31_out;
logic cond31_done;
logic cond_wire31_in;
logic cond_wire31_out;
logic cond32_in;
logic cond32_write_en;
logic cond32_clk;
logic cond32_reset;
logic cond32_out;
logic cond32_done;
logic cond_wire32_in;
logic cond_wire32_out;
logic cond33_in;
logic cond33_write_en;
logic cond33_clk;
logic cond33_reset;
logic cond33_out;
logic cond33_done;
logic cond_wire33_in;
logic cond_wire33_out;
logic cond34_in;
logic cond34_write_en;
logic cond34_clk;
logic cond34_reset;
logic cond34_out;
logic cond34_done;
logic cond_wire34_in;
logic cond_wire34_out;
logic cond35_in;
logic cond35_write_en;
logic cond35_clk;
logic cond35_reset;
logic cond35_out;
logic cond35_done;
logic cond_wire35_in;
logic cond_wire35_out;
logic cond36_in;
logic cond36_write_en;
logic cond36_clk;
logic cond36_reset;
logic cond36_out;
logic cond36_done;
logic cond_wire36_in;
logic cond_wire36_out;
logic cond37_in;
logic cond37_write_en;
logic cond37_clk;
logic cond37_reset;
logic cond37_out;
logic cond37_done;
logic cond_wire37_in;
logic cond_wire37_out;
logic cond38_in;
logic cond38_write_en;
logic cond38_clk;
logic cond38_reset;
logic cond38_out;
logic cond38_done;
logic cond_wire38_in;
logic cond_wire38_out;
logic cond39_in;
logic cond39_write_en;
logic cond39_clk;
logic cond39_reset;
logic cond39_out;
logic cond39_done;
logic cond_wire39_in;
logic cond_wire39_out;
logic cond40_in;
logic cond40_write_en;
logic cond40_clk;
logic cond40_reset;
logic cond40_out;
logic cond40_done;
logic cond_wire40_in;
logic cond_wire40_out;
logic cond41_in;
logic cond41_write_en;
logic cond41_clk;
logic cond41_reset;
logic cond41_out;
logic cond41_done;
logic cond_wire41_in;
logic cond_wire41_out;
logic cond42_in;
logic cond42_write_en;
logic cond42_clk;
logic cond42_reset;
logic cond42_out;
logic cond42_done;
logic cond_wire42_in;
logic cond_wire42_out;
logic cond43_in;
logic cond43_write_en;
logic cond43_clk;
logic cond43_reset;
logic cond43_out;
logic cond43_done;
logic cond_wire43_in;
logic cond_wire43_out;
logic cond44_in;
logic cond44_write_en;
logic cond44_clk;
logic cond44_reset;
logic cond44_out;
logic cond44_done;
logic cond_wire44_in;
logic cond_wire44_out;
logic cond45_in;
logic cond45_write_en;
logic cond45_clk;
logic cond45_reset;
logic cond45_out;
logic cond45_done;
logic cond_wire45_in;
logic cond_wire45_out;
logic cond46_in;
logic cond46_write_en;
logic cond46_clk;
logic cond46_reset;
logic cond46_out;
logic cond46_done;
logic cond_wire46_in;
logic cond_wire46_out;
logic cond47_in;
logic cond47_write_en;
logic cond47_clk;
logic cond47_reset;
logic cond47_out;
logic cond47_done;
logic cond_wire47_in;
logic cond_wire47_out;
logic cond48_in;
logic cond48_write_en;
logic cond48_clk;
logic cond48_reset;
logic cond48_out;
logic cond48_done;
logic cond_wire48_in;
logic cond_wire48_out;
logic cond49_in;
logic cond49_write_en;
logic cond49_clk;
logic cond49_reset;
logic cond49_out;
logic cond49_done;
logic cond_wire49_in;
logic cond_wire49_out;
logic cond50_in;
logic cond50_write_en;
logic cond50_clk;
logic cond50_reset;
logic cond50_out;
logic cond50_done;
logic cond_wire50_in;
logic cond_wire50_out;
logic cond51_in;
logic cond51_write_en;
logic cond51_clk;
logic cond51_reset;
logic cond51_out;
logic cond51_done;
logic cond_wire51_in;
logic cond_wire51_out;
logic cond52_in;
logic cond52_write_en;
logic cond52_clk;
logic cond52_reset;
logic cond52_out;
logic cond52_done;
logic cond_wire52_in;
logic cond_wire52_out;
logic cond53_in;
logic cond53_write_en;
logic cond53_clk;
logic cond53_reset;
logic cond53_out;
logic cond53_done;
logic cond_wire53_in;
logic cond_wire53_out;
logic cond54_in;
logic cond54_write_en;
logic cond54_clk;
logic cond54_reset;
logic cond54_out;
logic cond54_done;
logic cond_wire54_in;
logic cond_wire54_out;
logic cond55_in;
logic cond55_write_en;
logic cond55_clk;
logic cond55_reset;
logic cond55_out;
logic cond55_done;
logic cond_wire55_in;
logic cond_wire55_out;
logic cond56_in;
logic cond56_write_en;
logic cond56_clk;
logic cond56_reset;
logic cond56_out;
logic cond56_done;
logic cond_wire56_in;
logic cond_wire56_out;
logic cond57_in;
logic cond57_write_en;
logic cond57_clk;
logic cond57_reset;
logic cond57_out;
logic cond57_done;
logic cond_wire57_in;
logic cond_wire57_out;
logic cond58_in;
logic cond58_write_en;
logic cond58_clk;
logic cond58_reset;
logic cond58_out;
logic cond58_done;
logic cond_wire58_in;
logic cond_wire58_out;
logic cond59_in;
logic cond59_write_en;
logic cond59_clk;
logic cond59_reset;
logic cond59_out;
logic cond59_done;
logic cond_wire59_in;
logic cond_wire59_out;
logic cond60_in;
logic cond60_write_en;
logic cond60_clk;
logic cond60_reset;
logic cond60_out;
logic cond60_done;
logic cond_wire60_in;
logic cond_wire60_out;
logic cond61_in;
logic cond61_write_en;
logic cond61_clk;
logic cond61_reset;
logic cond61_out;
logic cond61_done;
logic cond_wire61_in;
logic cond_wire61_out;
logic cond62_in;
logic cond62_write_en;
logic cond62_clk;
logic cond62_reset;
logic cond62_out;
logic cond62_done;
logic cond_wire62_in;
logic cond_wire62_out;
logic cond63_in;
logic cond63_write_en;
logic cond63_clk;
logic cond63_reset;
logic cond63_out;
logic cond63_done;
logic cond_wire63_in;
logic cond_wire63_out;
logic cond64_in;
logic cond64_write_en;
logic cond64_clk;
logic cond64_reset;
logic cond64_out;
logic cond64_done;
logic cond_wire64_in;
logic cond_wire64_out;
logic cond65_in;
logic cond65_write_en;
logic cond65_clk;
logic cond65_reset;
logic cond65_out;
logic cond65_done;
logic cond_wire65_in;
logic cond_wire65_out;
logic cond66_in;
logic cond66_write_en;
logic cond66_clk;
logic cond66_reset;
logic cond66_out;
logic cond66_done;
logic cond_wire66_in;
logic cond_wire66_out;
logic cond67_in;
logic cond67_write_en;
logic cond67_clk;
logic cond67_reset;
logic cond67_out;
logic cond67_done;
logic cond_wire67_in;
logic cond_wire67_out;
logic cond68_in;
logic cond68_write_en;
logic cond68_clk;
logic cond68_reset;
logic cond68_out;
logic cond68_done;
logic cond_wire68_in;
logic cond_wire68_out;
logic fsm_in;
logic fsm_write_en;
logic fsm_clk;
logic fsm_reset;
logic fsm_out;
logic fsm_done;
logic [4:0] fsm0_in;
logic fsm0_write_en;
logic fsm0_clk;
logic fsm0_reset;
logic [4:0] fsm0_out;
logic fsm0_done;
logic ud_out;
logic [4:0] adder_left;
logic [4:0] adder_right;
logic [4:0] adder_out;
logic ud0_out;
logic adder0_left;
logic adder0_right;
logic adder0_out;
logic signal_reg_in;
logic signal_reg_write_en;
logic signal_reg_clk;
logic signal_reg_reset;
logic signal_reg_out;
logic signal_reg_done;
logic early_reset_static_seq_go_in;
logic early_reset_static_seq_go_out;
logic early_reset_static_seq_done_in;
logic early_reset_static_seq_done_out;
logic early_reset_static_par0_go_in;
logic early_reset_static_par0_go_out;
logic early_reset_static_par0_done_in;
logic early_reset_static_par0_done_out;
logic wrapper_early_reset_static_seq_go_in;
logic wrapper_early_reset_static_seq_go_out;
logic wrapper_early_reset_static_seq_done_in;
logic wrapper_early_reset_static_seq_done_out;
mac_pe pe_0_0 (
    .clk(pe_0_0_clk),
    .done(pe_0_0_done),
    .go(pe_0_0_go),
    .left(pe_0_0_left),
    .mul_ready(pe_0_0_mul_ready),
    .out(pe_0_0_out),
    .reset(pe_0_0_reset),
    .top(pe_0_0_top)
);
std_reg # (
    .WIDTH(32)
) top_0_0 (
    .clk(top_0_0_clk),
    .done(top_0_0_done),
    .in(top_0_0_in),
    .out(top_0_0_out),
    .reset(top_0_0_reset),
    .write_en(top_0_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_0 (
    .clk(left_0_0_clk),
    .done(left_0_0_done),
    .in(left_0_0_in),
    .out(left_0_0_out),
    .reset(left_0_0_reset),
    .write_en(left_0_0_write_en)
);
mac_pe pe_0_1 (
    .clk(pe_0_1_clk),
    .done(pe_0_1_done),
    .go(pe_0_1_go),
    .left(pe_0_1_left),
    .mul_ready(pe_0_1_mul_ready),
    .out(pe_0_1_out),
    .reset(pe_0_1_reset),
    .top(pe_0_1_top)
);
std_reg # (
    .WIDTH(32)
) top_0_1 (
    .clk(top_0_1_clk),
    .done(top_0_1_done),
    .in(top_0_1_in),
    .out(top_0_1_out),
    .reset(top_0_1_reset),
    .write_en(top_0_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_1 (
    .clk(left_0_1_clk),
    .done(left_0_1_done),
    .in(left_0_1_in),
    .out(left_0_1_out),
    .reset(left_0_1_reset),
    .write_en(left_0_1_write_en)
);
mac_pe pe_0_2 (
    .clk(pe_0_2_clk),
    .done(pe_0_2_done),
    .go(pe_0_2_go),
    .left(pe_0_2_left),
    .mul_ready(pe_0_2_mul_ready),
    .out(pe_0_2_out),
    .reset(pe_0_2_reset),
    .top(pe_0_2_top)
);
std_reg # (
    .WIDTH(32)
) top_0_2 (
    .clk(top_0_2_clk),
    .done(top_0_2_done),
    .in(top_0_2_in),
    .out(top_0_2_out),
    .reset(top_0_2_reset),
    .write_en(top_0_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_2 (
    .clk(left_0_2_clk),
    .done(left_0_2_done),
    .in(left_0_2_in),
    .out(left_0_2_out),
    .reset(left_0_2_reset),
    .write_en(left_0_2_write_en)
);
mac_pe pe_0_3 (
    .clk(pe_0_3_clk),
    .done(pe_0_3_done),
    .go(pe_0_3_go),
    .left(pe_0_3_left),
    .mul_ready(pe_0_3_mul_ready),
    .out(pe_0_3_out),
    .reset(pe_0_3_reset),
    .top(pe_0_3_top)
);
std_reg # (
    .WIDTH(32)
) top_0_3 (
    .clk(top_0_3_clk),
    .done(top_0_3_done),
    .in(top_0_3_in),
    .out(top_0_3_out),
    .reset(top_0_3_reset),
    .write_en(top_0_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_0_3 (
    .clk(left_0_3_clk),
    .done(left_0_3_done),
    .in(left_0_3_in),
    .out(left_0_3_out),
    .reset(left_0_3_reset),
    .write_en(left_0_3_write_en)
);
mac_pe pe_1_0 (
    .clk(pe_1_0_clk),
    .done(pe_1_0_done),
    .go(pe_1_0_go),
    .left(pe_1_0_left),
    .mul_ready(pe_1_0_mul_ready),
    .out(pe_1_0_out),
    .reset(pe_1_0_reset),
    .top(pe_1_0_top)
);
std_reg # (
    .WIDTH(32)
) top_1_0 (
    .clk(top_1_0_clk),
    .done(top_1_0_done),
    .in(top_1_0_in),
    .out(top_1_0_out),
    .reset(top_1_0_reset),
    .write_en(top_1_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_0 (
    .clk(left_1_0_clk),
    .done(left_1_0_done),
    .in(left_1_0_in),
    .out(left_1_0_out),
    .reset(left_1_0_reset),
    .write_en(left_1_0_write_en)
);
mac_pe pe_1_1 (
    .clk(pe_1_1_clk),
    .done(pe_1_1_done),
    .go(pe_1_1_go),
    .left(pe_1_1_left),
    .mul_ready(pe_1_1_mul_ready),
    .out(pe_1_1_out),
    .reset(pe_1_1_reset),
    .top(pe_1_1_top)
);
std_reg # (
    .WIDTH(32)
) top_1_1 (
    .clk(top_1_1_clk),
    .done(top_1_1_done),
    .in(top_1_1_in),
    .out(top_1_1_out),
    .reset(top_1_1_reset),
    .write_en(top_1_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_1 (
    .clk(left_1_1_clk),
    .done(left_1_1_done),
    .in(left_1_1_in),
    .out(left_1_1_out),
    .reset(left_1_1_reset),
    .write_en(left_1_1_write_en)
);
mac_pe pe_1_2 (
    .clk(pe_1_2_clk),
    .done(pe_1_2_done),
    .go(pe_1_2_go),
    .left(pe_1_2_left),
    .mul_ready(pe_1_2_mul_ready),
    .out(pe_1_2_out),
    .reset(pe_1_2_reset),
    .top(pe_1_2_top)
);
std_reg # (
    .WIDTH(32)
) top_1_2 (
    .clk(top_1_2_clk),
    .done(top_1_2_done),
    .in(top_1_2_in),
    .out(top_1_2_out),
    .reset(top_1_2_reset),
    .write_en(top_1_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_2 (
    .clk(left_1_2_clk),
    .done(left_1_2_done),
    .in(left_1_2_in),
    .out(left_1_2_out),
    .reset(left_1_2_reset),
    .write_en(left_1_2_write_en)
);
mac_pe pe_1_3 (
    .clk(pe_1_3_clk),
    .done(pe_1_3_done),
    .go(pe_1_3_go),
    .left(pe_1_3_left),
    .mul_ready(pe_1_3_mul_ready),
    .out(pe_1_3_out),
    .reset(pe_1_3_reset),
    .top(pe_1_3_top)
);
std_reg # (
    .WIDTH(32)
) top_1_3 (
    .clk(top_1_3_clk),
    .done(top_1_3_done),
    .in(top_1_3_in),
    .out(top_1_3_out),
    .reset(top_1_3_reset),
    .write_en(top_1_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_1_3 (
    .clk(left_1_3_clk),
    .done(left_1_3_done),
    .in(left_1_3_in),
    .out(left_1_3_out),
    .reset(left_1_3_reset),
    .write_en(left_1_3_write_en)
);
mac_pe pe_2_0 (
    .clk(pe_2_0_clk),
    .done(pe_2_0_done),
    .go(pe_2_0_go),
    .left(pe_2_0_left),
    .mul_ready(pe_2_0_mul_ready),
    .out(pe_2_0_out),
    .reset(pe_2_0_reset),
    .top(pe_2_0_top)
);
std_reg # (
    .WIDTH(32)
) top_2_0 (
    .clk(top_2_0_clk),
    .done(top_2_0_done),
    .in(top_2_0_in),
    .out(top_2_0_out),
    .reset(top_2_0_reset),
    .write_en(top_2_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_0 (
    .clk(left_2_0_clk),
    .done(left_2_0_done),
    .in(left_2_0_in),
    .out(left_2_0_out),
    .reset(left_2_0_reset),
    .write_en(left_2_0_write_en)
);
mac_pe pe_2_1 (
    .clk(pe_2_1_clk),
    .done(pe_2_1_done),
    .go(pe_2_1_go),
    .left(pe_2_1_left),
    .mul_ready(pe_2_1_mul_ready),
    .out(pe_2_1_out),
    .reset(pe_2_1_reset),
    .top(pe_2_1_top)
);
std_reg # (
    .WIDTH(32)
) top_2_1 (
    .clk(top_2_1_clk),
    .done(top_2_1_done),
    .in(top_2_1_in),
    .out(top_2_1_out),
    .reset(top_2_1_reset),
    .write_en(top_2_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_1 (
    .clk(left_2_1_clk),
    .done(left_2_1_done),
    .in(left_2_1_in),
    .out(left_2_1_out),
    .reset(left_2_1_reset),
    .write_en(left_2_1_write_en)
);
mac_pe pe_2_2 (
    .clk(pe_2_2_clk),
    .done(pe_2_2_done),
    .go(pe_2_2_go),
    .left(pe_2_2_left),
    .mul_ready(pe_2_2_mul_ready),
    .out(pe_2_2_out),
    .reset(pe_2_2_reset),
    .top(pe_2_2_top)
);
std_reg # (
    .WIDTH(32)
) top_2_2 (
    .clk(top_2_2_clk),
    .done(top_2_2_done),
    .in(top_2_2_in),
    .out(top_2_2_out),
    .reset(top_2_2_reset),
    .write_en(top_2_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_2 (
    .clk(left_2_2_clk),
    .done(left_2_2_done),
    .in(left_2_2_in),
    .out(left_2_2_out),
    .reset(left_2_2_reset),
    .write_en(left_2_2_write_en)
);
mac_pe pe_2_3 (
    .clk(pe_2_3_clk),
    .done(pe_2_3_done),
    .go(pe_2_3_go),
    .left(pe_2_3_left),
    .mul_ready(pe_2_3_mul_ready),
    .out(pe_2_3_out),
    .reset(pe_2_3_reset),
    .top(pe_2_3_top)
);
std_reg # (
    .WIDTH(32)
) top_2_3 (
    .clk(top_2_3_clk),
    .done(top_2_3_done),
    .in(top_2_3_in),
    .out(top_2_3_out),
    .reset(top_2_3_reset),
    .write_en(top_2_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_2_3 (
    .clk(left_2_3_clk),
    .done(left_2_3_done),
    .in(left_2_3_in),
    .out(left_2_3_out),
    .reset(left_2_3_reset),
    .write_en(left_2_3_write_en)
);
mac_pe pe_3_0 (
    .clk(pe_3_0_clk),
    .done(pe_3_0_done),
    .go(pe_3_0_go),
    .left(pe_3_0_left),
    .mul_ready(pe_3_0_mul_ready),
    .out(pe_3_0_out),
    .reset(pe_3_0_reset),
    .top(pe_3_0_top)
);
std_reg # (
    .WIDTH(32)
) top_3_0 (
    .clk(top_3_0_clk),
    .done(top_3_0_done),
    .in(top_3_0_in),
    .out(top_3_0_out),
    .reset(top_3_0_reset),
    .write_en(top_3_0_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_0 (
    .clk(left_3_0_clk),
    .done(left_3_0_done),
    .in(left_3_0_in),
    .out(left_3_0_out),
    .reset(left_3_0_reset),
    .write_en(left_3_0_write_en)
);
mac_pe pe_3_1 (
    .clk(pe_3_1_clk),
    .done(pe_3_1_done),
    .go(pe_3_1_go),
    .left(pe_3_1_left),
    .mul_ready(pe_3_1_mul_ready),
    .out(pe_3_1_out),
    .reset(pe_3_1_reset),
    .top(pe_3_1_top)
);
std_reg # (
    .WIDTH(32)
) top_3_1 (
    .clk(top_3_1_clk),
    .done(top_3_1_done),
    .in(top_3_1_in),
    .out(top_3_1_out),
    .reset(top_3_1_reset),
    .write_en(top_3_1_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_1 (
    .clk(left_3_1_clk),
    .done(left_3_1_done),
    .in(left_3_1_in),
    .out(left_3_1_out),
    .reset(left_3_1_reset),
    .write_en(left_3_1_write_en)
);
mac_pe pe_3_2 (
    .clk(pe_3_2_clk),
    .done(pe_3_2_done),
    .go(pe_3_2_go),
    .left(pe_3_2_left),
    .mul_ready(pe_3_2_mul_ready),
    .out(pe_3_2_out),
    .reset(pe_3_2_reset),
    .top(pe_3_2_top)
);
std_reg # (
    .WIDTH(32)
) top_3_2 (
    .clk(top_3_2_clk),
    .done(top_3_2_done),
    .in(top_3_2_in),
    .out(top_3_2_out),
    .reset(top_3_2_reset),
    .write_en(top_3_2_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_2 (
    .clk(left_3_2_clk),
    .done(left_3_2_done),
    .in(left_3_2_in),
    .out(left_3_2_out),
    .reset(left_3_2_reset),
    .write_en(left_3_2_write_en)
);
mac_pe pe_3_3 (
    .clk(pe_3_3_clk),
    .done(pe_3_3_done),
    .go(pe_3_3_go),
    .left(pe_3_3_left),
    .mul_ready(pe_3_3_mul_ready),
    .out(pe_3_3_out),
    .reset(pe_3_3_reset),
    .top(pe_3_3_top)
);
std_reg # (
    .WIDTH(32)
) top_3_3 (
    .clk(top_3_3_clk),
    .done(top_3_3_done),
    .in(top_3_3_in),
    .out(top_3_3_out),
    .reset(top_3_3_reset),
    .write_en(top_3_3_write_en)
);
std_reg # (
    .WIDTH(32)
) left_3_3 (
    .clk(left_3_3_clk),
    .done(left_3_3_done),
    .in(left_3_3_in),
    .out(left_3_3_out),
    .reset(left_3_3_reset),
    .write_en(left_3_3_write_en)
);
std_reg # (
    .WIDTH(3)
) t0_idx (
    .clk(t0_idx_clk),
    .done(t0_idx_done),
    .in(t0_idx_in),
    .out(t0_idx_out),
    .reset(t0_idx_reset),
    .write_en(t0_idx_write_en)
);
std_add # (
    .WIDTH(3)
) t0_add (
    .left(t0_add_left),
    .out(t0_add_out),
    .right(t0_add_right)
);
std_reg # (
    .WIDTH(3)
) t1_idx (
    .clk(t1_idx_clk),
    .done(t1_idx_done),
    .in(t1_idx_in),
    .out(t1_idx_out),
    .reset(t1_idx_reset),
    .write_en(t1_idx_write_en)
);
std_add # (
    .WIDTH(3)
) t1_add (
    .left(t1_add_left),
    .out(t1_add_out),
    .right(t1_add_right)
);
std_reg # (
    .WIDTH(3)
) t2_idx (
    .clk(t2_idx_clk),
    .done(t2_idx_done),
    .in(t2_idx_in),
    .out(t2_idx_out),
    .reset(t2_idx_reset),
    .write_en(t2_idx_write_en)
);
std_add # (
    .WIDTH(3)
) t2_add (
    .left(t2_add_left),
    .out(t2_add_out),
    .right(t2_add_right)
);
std_reg # (
    .WIDTH(3)
) t3_idx (
    .clk(t3_idx_clk),
    .done(t3_idx_done),
    .in(t3_idx_in),
    .out(t3_idx_out),
    .reset(t3_idx_reset),
    .write_en(t3_idx_write_en)
);
std_add # (
    .WIDTH(3)
) t3_add (
    .left(t3_add_left),
    .out(t3_add_out),
    .right(t3_add_right)
);
std_reg # (
    .WIDTH(3)
) l0_idx (
    .clk(l0_idx_clk),
    .done(l0_idx_done),
    .in(l0_idx_in),
    .out(l0_idx_out),
    .reset(l0_idx_reset),
    .write_en(l0_idx_write_en)
);
std_add # (
    .WIDTH(3)
) l0_add (
    .left(l0_add_left),
    .out(l0_add_out),
    .right(l0_add_right)
);
std_reg # (
    .WIDTH(3)
) l1_idx (
    .clk(l1_idx_clk),
    .done(l1_idx_done),
    .in(l1_idx_in),
    .out(l1_idx_out),
    .reset(l1_idx_reset),
    .write_en(l1_idx_write_en)
);
std_add # (
    .WIDTH(3)
) l1_add (
    .left(l1_add_left),
    .out(l1_add_out),
    .right(l1_add_right)
);
std_reg # (
    .WIDTH(3)
) l2_idx (
    .clk(l2_idx_clk),
    .done(l2_idx_done),
    .in(l2_idx_in),
    .out(l2_idx_out),
    .reset(l2_idx_reset),
    .write_en(l2_idx_write_en)
);
std_add # (
    .WIDTH(3)
) l2_add (
    .left(l2_add_left),
    .out(l2_add_out),
    .right(l2_add_right)
);
std_reg # (
    .WIDTH(3)
) l3_idx (
    .clk(l3_idx_clk),
    .done(l3_idx_done),
    .in(l3_idx_in),
    .out(l3_idx_out),
    .reset(l3_idx_reset),
    .write_en(l3_idx_write_en)
);
std_add # (
    .WIDTH(3)
) l3_add (
    .left(l3_add_left),
    .out(l3_add_out),
    .right(l3_add_right)
);
std_reg # (
    .WIDTH(5)
) idx (
    .clk(idx_clk),
    .done(idx_done),
    .in(idx_in),
    .out(idx_out),
    .reset(idx_reset),
    .write_en(idx_write_en)
);
std_add # (
    .WIDTH(5)
) idx_add (
    .left(idx_add_left),
    .out(idx_add_out),
    .right(idx_add_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_3_7_reg (
    .clk(idx_between_3_7_reg_clk),
    .done(idx_between_3_7_reg_done),
    .in(idx_between_3_7_reg_in),
    .out(idx_between_3_7_reg_out),
    .reset(idx_between_3_7_reg_reset),
    .write_en(idx_between_3_7_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_7 (
    .left(index_lt_7_left),
    .out(index_lt_7_out),
    .right(index_lt_7_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_3 (
    .left(index_ge_3_left),
    .out(index_ge_3_out),
    .right(index_ge_3_right)
);
std_and # (
    .WIDTH(1)
) idx_between_3_7_comb (
    .left(idx_between_3_7_comb_left),
    .out(idx_between_3_7_comb_out),
    .right(idx_between_3_7_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_12_13_reg (
    .clk(idx_between_12_13_reg_clk),
    .done(idx_between_12_13_reg_done),
    .in(idx_between_12_13_reg_in),
    .out(idx_between_12_13_reg_out),
    .reset(idx_between_12_13_reg_reset),
    .write_en(idx_between_12_13_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_13 (
    .left(index_lt_13_left),
    .out(index_lt_13_out),
    .right(index_lt_13_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_12 (
    .left(index_ge_12_left),
    .out(index_ge_12_out),
    .right(index_ge_12_right)
);
std_and # (
    .WIDTH(1)
) idx_between_12_13_comb (
    .left(idx_between_12_13_comb_left),
    .out(idx_between_12_13_comb_out),
    .right(idx_between_12_13_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_8_12_reg (
    .clk(idx_between_8_12_reg_clk),
    .done(idx_between_8_12_reg_done),
    .in(idx_between_8_12_reg_in),
    .out(idx_between_8_12_reg_out),
    .reset(idx_between_8_12_reg_reset),
    .write_en(idx_between_8_12_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_12 (
    .left(index_lt_12_left),
    .out(index_lt_12_out),
    .right(index_lt_12_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_8 (
    .left(index_ge_8_left),
    .out(index_ge_8_out),
    .right(index_ge_8_right)
);
std_and # (
    .WIDTH(1)
) idx_between_8_12_comb (
    .left(idx_between_8_12_comb_left),
    .out(idx_between_8_12_comb_out),
    .right(idx_between_8_12_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_13_14_reg (
    .clk(idx_between_13_14_reg_clk),
    .done(idx_between_13_14_reg_done),
    .in(idx_between_13_14_reg_in),
    .out(idx_between_13_14_reg_out),
    .reset(idx_between_13_14_reg_reset),
    .write_en(idx_between_13_14_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_14 (
    .left(index_lt_14_left),
    .out(index_lt_14_out),
    .right(index_lt_14_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_13 (
    .left(index_ge_13_left),
    .out(index_ge_13_out),
    .right(index_ge_13_right)
);
std_and # (
    .WIDTH(1)
) idx_between_13_14_comb (
    .left(idx_between_13_14_comb_left),
    .out(idx_between_13_14_comb_out),
    .right(idx_between_13_14_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_4_8_reg (
    .clk(idx_between_4_8_reg_clk),
    .done(idx_between_4_8_reg_done),
    .in(idx_between_4_8_reg_in),
    .out(idx_between_4_8_reg_out),
    .reset(idx_between_4_8_reg_reset),
    .write_en(idx_between_4_8_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_8 (
    .left(index_lt_8_left),
    .out(index_lt_8_out),
    .right(index_lt_8_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_4 (
    .left(index_ge_4_left),
    .out(index_ge_4_out),
    .right(index_ge_4_right)
);
std_and # (
    .WIDTH(1)
) idx_between_4_8_comb (
    .left(idx_between_4_8_comb_left),
    .out(idx_between_4_8_comb_out),
    .right(idx_between_4_8_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_5_9_reg (
    .clk(idx_between_5_9_reg_clk),
    .done(idx_between_5_9_reg_done),
    .in(idx_between_5_9_reg_in),
    .out(idx_between_5_9_reg_out),
    .reset(idx_between_5_9_reg_reset),
    .write_en(idx_between_5_9_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_9 (
    .left(index_lt_9_left),
    .out(index_lt_9_out),
    .right(index_lt_9_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_5 (
    .left(index_ge_5_left),
    .out(index_ge_5_out),
    .right(index_ge_5_right)
);
std_and # (
    .WIDTH(1)
) idx_between_5_9_comb (
    .left(idx_between_5_9_comb_left),
    .out(idx_between_5_9_comb_out),
    .right(idx_between_5_9_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_14_15_reg (
    .clk(idx_between_14_15_reg_clk),
    .done(idx_between_14_15_reg_done),
    .in(idx_between_14_15_reg_in),
    .out(idx_between_14_15_reg_out),
    .reset(idx_between_14_15_reg_reset),
    .write_en(idx_between_14_15_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_15 (
    .left(index_lt_15_left),
    .out(index_lt_15_out),
    .right(index_lt_15_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_14 (
    .left(index_ge_14_left),
    .out(index_ge_14_out),
    .right(index_ge_14_right)
);
std_and # (
    .WIDTH(1)
) idx_between_14_15_comb (
    .left(idx_between_14_15_comb_left),
    .out(idx_between_14_15_comb_out),
    .right(idx_between_14_15_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_9_10_reg (
    .clk(idx_between_9_10_reg_clk),
    .done(idx_between_9_10_reg_done),
    .in(idx_between_9_10_reg_in),
    .out(idx_between_9_10_reg_out),
    .reset(idx_between_9_10_reg_reset),
    .write_en(idx_between_9_10_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_10 (
    .left(index_lt_10_left),
    .out(index_lt_10_out),
    .right(index_lt_10_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_9 (
    .left(index_ge_9_left),
    .out(index_ge_9_out),
    .right(index_ge_9_right)
);
std_and # (
    .WIDTH(1)
) idx_between_9_10_comb (
    .left(idx_between_9_10_comb_left),
    .out(idx_between_9_10_comb_out),
    .right(idx_between_9_10_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_10_11_reg (
    .clk(idx_between_10_11_reg_clk),
    .done(idx_between_10_11_reg_done),
    .in(idx_between_10_11_reg_in),
    .out(idx_between_10_11_reg_out),
    .reset(idx_between_10_11_reg_reset),
    .write_en(idx_between_10_11_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_11 (
    .left(index_lt_11_left),
    .out(index_lt_11_out),
    .right(index_lt_11_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_10 (
    .left(index_ge_10_left),
    .out(index_ge_10_out),
    .right(index_ge_10_right)
);
std_and # (
    .WIDTH(1)
) idx_between_10_11_comb (
    .left(idx_between_10_11_comb_left),
    .out(idx_between_10_11_comb_out),
    .right(idx_between_10_11_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_0_4_reg (
    .clk(idx_between_0_4_reg_clk),
    .done(idx_between_0_4_reg_done),
    .in(idx_between_0_4_reg_in),
    .out(idx_between_0_4_reg_out),
    .reset(idx_between_0_4_reg_reset),
    .write_en(idx_between_0_4_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_4 (
    .left(index_lt_4_left),
    .out(index_lt_4_out),
    .right(index_lt_4_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_9_13_reg (
    .clk(idx_between_9_13_reg_clk),
    .done(idx_between_9_13_reg_done),
    .in(idx_between_9_13_reg_in),
    .out(idx_between_9_13_reg_out),
    .reset(idx_between_9_13_reg_reset),
    .write_en(idx_between_9_13_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_9_13_comb (
    .left(idx_between_9_13_comb_left),
    .out(idx_between_9_13_comb_out),
    .right(idx_between_9_13_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_1_5_reg (
    .clk(idx_between_1_5_reg_clk),
    .done(idx_between_1_5_reg_done),
    .in(idx_between_1_5_reg_in),
    .out(idx_between_1_5_reg_out),
    .reset(idx_between_1_5_reg_reset),
    .write_en(idx_between_1_5_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_5 (
    .left(index_lt_5_left),
    .out(index_lt_5_out),
    .right(index_lt_5_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_1 (
    .left(index_ge_1_left),
    .out(index_ge_1_out),
    .right(index_ge_1_right)
);
std_and # (
    .WIDTH(1)
) idx_between_1_5_comb (
    .left(idx_between_1_5_comb_left),
    .out(idx_between_1_5_comb_out),
    .right(idx_between_1_5_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_10_14_reg (
    .clk(idx_between_10_14_reg_clk),
    .done(idx_between_10_14_reg_done),
    .in(idx_between_10_14_reg_in),
    .out(idx_between_10_14_reg_out),
    .reset(idx_between_10_14_reg_reset),
    .write_en(idx_between_10_14_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_10_14_comb (
    .left(idx_between_10_14_comb_left),
    .out(idx_between_10_14_comb_out),
    .right(idx_between_10_14_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_15_16_reg (
    .clk(idx_between_15_16_reg_clk),
    .done(idx_between_15_16_reg_done),
    .in(idx_between_15_16_reg_in),
    .out(idx_between_15_16_reg_out),
    .reset(idx_between_15_16_reg_reset),
    .write_en(idx_between_15_16_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_16 (
    .left(index_lt_16_left),
    .out(index_lt_16_out),
    .right(index_lt_16_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_15 (
    .left(index_ge_15_left),
    .out(index_ge_15_out),
    .right(index_ge_15_right)
);
std_and # (
    .WIDTH(1)
) idx_between_15_16_comb (
    .left(idx_between_15_16_comb_left),
    .out(idx_between_15_16_comb_out),
    .right(idx_between_15_16_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_6_10_reg (
    .clk(idx_between_6_10_reg_clk),
    .done(idx_between_6_10_reg_done),
    .in(idx_between_6_10_reg_in),
    .out(idx_between_6_10_reg_out),
    .reset(idx_between_6_10_reg_reset),
    .write_en(idx_between_6_10_reg_write_en)
);
std_ge # (
    .WIDTH(5)
) index_ge_6 (
    .left(index_ge_6_left),
    .out(index_ge_6_out),
    .right(index_ge_6_right)
);
std_and # (
    .WIDTH(1)
) idx_between_6_10_comb (
    .left(idx_between_6_10_comb_left),
    .out(idx_between_6_10_comb_out),
    .right(idx_between_6_10_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_11_12_reg (
    .clk(idx_between_11_12_reg_clk),
    .done(idx_between_11_12_reg_done),
    .in(idx_between_11_12_reg_in),
    .out(idx_between_11_12_reg_out),
    .reset(idx_between_11_12_reg_reset),
    .write_en(idx_between_11_12_reg_write_en)
);
std_ge # (
    .WIDTH(5)
) index_ge_11 (
    .left(index_ge_11_left),
    .out(index_ge_11_out),
    .right(index_ge_11_right)
);
std_and # (
    .WIDTH(1)
) idx_between_11_12_comb (
    .left(idx_between_11_12_comb_left),
    .out(idx_between_11_12_comb_out),
    .right(idx_between_11_12_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_2_6_reg (
    .clk(idx_between_2_6_reg_clk),
    .done(idx_between_2_6_reg_done),
    .in(idx_between_2_6_reg_in),
    .out(idx_between_2_6_reg_out),
    .reset(idx_between_2_6_reg_reset),
    .write_en(idx_between_2_6_reg_write_en)
);
std_lt # (
    .WIDTH(5)
) index_lt_6 (
    .left(index_lt_6_left),
    .out(index_lt_6_out),
    .right(index_lt_6_right)
);
std_ge # (
    .WIDTH(5)
) index_ge_2 (
    .left(index_ge_2_left),
    .out(index_ge_2_out),
    .right(index_ge_2_right)
);
std_and # (
    .WIDTH(1)
) idx_between_2_6_comb (
    .left(idx_between_2_6_comb_left),
    .out(idx_between_2_6_comb_out),
    .right(idx_between_2_6_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_11_15_reg (
    .clk(idx_between_11_15_reg_clk),
    .done(idx_between_11_15_reg_done),
    .in(idx_between_11_15_reg_in),
    .out(idx_between_11_15_reg_out),
    .reset(idx_between_11_15_reg_reset),
    .write_en(idx_between_11_15_reg_write_en)
);
std_and # (
    .WIDTH(1)
) idx_between_11_15_comb (
    .left(idx_between_11_15_comb_left),
    .out(idx_between_11_15_comb_out),
    .right(idx_between_11_15_comb_right)
);
std_reg # (
    .WIDTH(1)
) idx_between_7_11_reg (
    .clk(idx_between_7_11_reg_clk),
    .done(idx_between_7_11_reg_done),
    .in(idx_between_7_11_reg_in),
    .out(idx_between_7_11_reg_out),
    .reset(idx_between_7_11_reg_reset),
    .write_en(idx_between_7_11_reg_write_en)
);
std_ge # (
    .WIDTH(5)
) index_ge_7 (
    .left(index_ge_7_left),
    .out(index_ge_7_out),
    .right(index_ge_7_right)
);
std_and # (
    .WIDTH(1)
) idx_between_7_11_comb (
    .left(idx_between_7_11_comb_left),
    .out(idx_between_7_11_comb_out),
    .right(idx_between_7_11_comb_right)
);
std_reg # (
    .WIDTH(1)
) cond (
    .clk(cond_clk),
    .done(cond_done),
    .in(cond_in),
    .out(cond_out),
    .reset(cond_reset),
    .write_en(cond_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire (
    .in(cond_wire_in),
    .out(cond_wire_out)
);
std_reg # (
    .WIDTH(1)
) cond0 (
    .clk(cond0_clk),
    .done(cond0_done),
    .in(cond0_in),
    .out(cond0_out),
    .reset(cond0_reset),
    .write_en(cond0_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire0 (
    .in(cond_wire0_in),
    .out(cond_wire0_out)
);
std_reg # (
    .WIDTH(1)
) cond1 (
    .clk(cond1_clk),
    .done(cond1_done),
    .in(cond1_in),
    .out(cond1_out),
    .reset(cond1_reset),
    .write_en(cond1_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire1 (
    .in(cond_wire1_in),
    .out(cond_wire1_out)
);
std_reg # (
    .WIDTH(1)
) cond2 (
    .clk(cond2_clk),
    .done(cond2_done),
    .in(cond2_in),
    .out(cond2_out),
    .reset(cond2_reset),
    .write_en(cond2_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire2 (
    .in(cond_wire2_in),
    .out(cond_wire2_out)
);
std_reg # (
    .WIDTH(1)
) cond3 (
    .clk(cond3_clk),
    .done(cond3_done),
    .in(cond3_in),
    .out(cond3_out),
    .reset(cond3_reset),
    .write_en(cond3_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire3 (
    .in(cond_wire3_in),
    .out(cond_wire3_out)
);
std_reg # (
    .WIDTH(1)
) cond4 (
    .clk(cond4_clk),
    .done(cond4_done),
    .in(cond4_in),
    .out(cond4_out),
    .reset(cond4_reset),
    .write_en(cond4_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire4 (
    .in(cond_wire4_in),
    .out(cond_wire4_out)
);
std_reg # (
    .WIDTH(1)
) cond5 (
    .clk(cond5_clk),
    .done(cond5_done),
    .in(cond5_in),
    .out(cond5_out),
    .reset(cond5_reset),
    .write_en(cond5_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire5 (
    .in(cond_wire5_in),
    .out(cond_wire5_out)
);
std_reg # (
    .WIDTH(1)
) cond6 (
    .clk(cond6_clk),
    .done(cond6_done),
    .in(cond6_in),
    .out(cond6_out),
    .reset(cond6_reset),
    .write_en(cond6_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire6 (
    .in(cond_wire6_in),
    .out(cond_wire6_out)
);
std_reg # (
    .WIDTH(1)
) cond7 (
    .clk(cond7_clk),
    .done(cond7_done),
    .in(cond7_in),
    .out(cond7_out),
    .reset(cond7_reset),
    .write_en(cond7_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire7 (
    .in(cond_wire7_in),
    .out(cond_wire7_out)
);
std_reg # (
    .WIDTH(1)
) cond8 (
    .clk(cond8_clk),
    .done(cond8_done),
    .in(cond8_in),
    .out(cond8_out),
    .reset(cond8_reset),
    .write_en(cond8_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire8 (
    .in(cond_wire8_in),
    .out(cond_wire8_out)
);
std_reg # (
    .WIDTH(1)
) cond9 (
    .clk(cond9_clk),
    .done(cond9_done),
    .in(cond9_in),
    .out(cond9_out),
    .reset(cond9_reset),
    .write_en(cond9_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire9 (
    .in(cond_wire9_in),
    .out(cond_wire9_out)
);
std_reg # (
    .WIDTH(1)
) cond10 (
    .clk(cond10_clk),
    .done(cond10_done),
    .in(cond10_in),
    .out(cond10_out),
    .reset(cond10_reset),
    .write_en(cond10_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire10 (
    .in(cond_wire10_in),
    .out(cond_wire10_out)
);
std_reg # (
    .WIDTH(1)
) cond11 (
    .clk(cond11_clk),
    .done(cond11_done),
    .in(cond11_in),
    .out(cond11_out),
    .reset(cond11_reset),
    .write_en(cond11_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire11 (
    .in(cond_wire11_in),
    .out(cond_wire11_out)
);
std_reg # (
    .WIDTH(1)
) cond12 (
    .clk(cond12_clk),
    .done(cond12_done),
    .in(cond12_in),
    .out(cond12_out),
    .reset(cond12_reset),
    .write_en(cond12_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire12 (
    .in(cond_wire12_in),
    .out(cond_wire12_out)
);
std_reg # (
    .WIDTH(1)
) cond13 (
    .clk(cond13_clk),
    .done(cond13_done),
    .in(cond13_in),
    .out(cond13_out),
    .reset(cond13_reset),
    .write_en(cond13_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire13 (
    .in(cond_wire13_in),
    .out(cond_wire13_out)
);
std_reg # (
    .WIDTH(1)
) cond14 (
    .clk(cond14_clk),
    .done(cond14_done),
    .in(cond14_in),
    .out(cond14_out),
    .reset(cond14_reset),
    .write_en(cond14_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire14 (
    .in(cond_wire14_in),
    .out(cond_wire14_out)
);
std_reg # (
    .WIDTH(1)
) cond15 (
    .clk(cond15_clk),
    .done(cond15_done),
    .in(cond15_in),
    .out(cond15_out),
    .reset(cond15_reset),
    .write_en(cond15_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire15 (
    .in(cond_wire15_in),
    .out(cond_wire15_out)
);
std_reg # (
    .WIDTH(1)
) cond16 (
    .clk(cond16_clk),
    .done(cond16_done),
    .in(cond16_in),
    .out(cond16_out),
    .reset(cond16_reset),
    .write_en(cond16_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire16 (
    .in(cond_wire16_in),
    .out(cond_wire16_out)
);
std_reg # (
    .WIDTH(1)
) cond17 (
    .clk(cond17_clk),
    .done(cond17_done),
    .in(cond17_in),
    .out(cond17_out),
    .reset(cond17_reset),
    .write_en(cond17_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire17 (
    .in(cond_wire17_in),
    .out(cond_wire17_out)
);
std_reg # (
    .WIDTH(1)
) cond18 (
    .clk(cond18_clk),
    .done(cond18_done),
    .in(cond18_in),
    .out(cond18_out),
    .reset(cond18_reset),
    .write_en(cond18_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire18 (
    .in(cond_wire18_in),
    .out(cond_wire18_out)
);
std_reg # (
    .WIDTH(1)
) cond19 (
    .clk(cond19_clk),
    .done(cond19_done),
    .in(cond19_in),
    .out(cond19_out),
    .reset(cond19_reset),
    .write_en(cond19_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire19 (
    .in(cond_wire19_in),
    .out(cond_wire19_out)
);
std_reg # (
    .WIDTH(1)
) cond20 (
    .clk(cond20_clk),
    .done(cond20_done),
    .in(cond20_in),
    .out(cond20_out),
    .reset(cond20_reset),
    .write_en(cond20_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire20 (
    .in(cond_wire20_in),
    .out(cond_wire20_out)
);
std_reg # (
    .WIDTH(1)
) cond21 (
    .clk(cond21_clk),
    .done(cond21_done),
    .in(cond21_in),
    .out(cond21_out),
    .reset(cond21_reset),
    .write_en(cond21_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire21 (
    .in(cond_wire21_in),
    .out(cond_wire21_out)
);
std_reg # (
    .WIDTH(1)
) cond22 (
    .clk(cond22_clk),
    .done(cond22_done),
    .in(cond22_in),
    .out(cond22_out),
    .reset(cond22_reset),
    .write_en(cond22_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire22 (
    .in(cond_wire22_in),
    .out(cond_wire22_out)
);
std_reg # (
    .WIDTH(1)
) cond23 (
    .clk(cond23_clk),
    .done(cond23_done),
    .in(cond23_in),
    .out(cond23_out),
    .reset(cond23_reset),
    .write_en(cond23_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire23 (
    .in(cond_wire23_in),
    .out(cond_wire23_out)
);
std_reg # (
    .WIDTH(1)
) cond24 (
    .clk(cond24_clk),
    .done(cond24_done),
    .in(cond24_in),
    .out(cond24_out),
    .reset(cond24_reset),
    .write_en(cond24_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire24 (
    .in(cond_wire24_in),
    .out(cond_wire24_out)
);
std_reg # (
    .WIDTH(1)
) cond25 (
    .clk(cond25_clk),
    .done(cond25_done),
    .in(cond25_in),
    .out(cond25_out),
    .reset(cond25_reset),
    .write_en(cond25_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire25 (
    .in(cond_wire25_in),
    .out(cond_wire25_out)
);
std_reg # (
    .WIDTH(1)
) cond26 (
    .clk(cond26_clk),
    .done(cond26_done),
    .in(cond26_in),
    .out(cond26_out),
    .reset(cond26_reset),
    .write_en(cond26_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire26 (
    .in(cond_wire26_in),
    .out(cond_wire26_out)
);
std_reg # (
    .WIDTH(1)
) cond27 (
    .clk(cond27_clk),
    .done(cond27_done),
    .in(cond27_in),
    .out(cond27_out),
    .reset(cond27_reset),
    .write_en(cond27_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire27 (
    .in(cond_wire27_in),
    .out(cond_wire27_out)
);
std_reg # (
    .WIDTH(1)
) cond28 (
    .clk(cond28_clk),
    .done(cond28_done),
    .in(cond28_in),
    .out(cond28_out),
    .reset(cond28_reset),
    .write_en(cond28_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire28 (
    .in(cond_wire28_in),
    .out(cond_wire28_out)
);
std_reg # (
    .WIDTH(1)
) cond29 (
    .clk(cond29_clk),
    .done(cond29_done),
    .in(cond29_in),
    .out(cond29_out),
    .reset(cond29_reset),
    .write_en(cond29_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire29 (
    .in(cond_wire29_in),
    .out(cond_wire29_out)
);
std_reg # (
    .WIDTH(1)
) cond30 (
    .clk(cond30_clk),
    .done(cond30_done),
    .in(cond30_in),
    .out(cond30_out),
    .reset(cond30_reset),
    .write_en(cond30_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire30 (
    .in(cond_wire30_in),
    .out(cond_wire30_out)
);
std_reg # (
    .WIDTH(1)
) cond31 (
    .clk(cond31_clk),
    .done(cond31_done),
    .in(cond31_in),
    .out(cond31_out),
    .reset(cond31_reset),
    .write_en(cond31_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire31 (
    .in(cond_wire31_in),
    .out(cond_wire31_out)
);
std_reg # (
    .WIDTH(1)
) cond32 (
    .clk(cond32_clk),
    .done(cond32_done),
    .in(cond32_in),
    .out(cond32_out),
    .reset(cond32_reset),
    .write_en(cond32_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire32 (
    .in(cond_wire32_in),
    .out(cond_wire32_out)
);
std_reg # (
    .WIDTH(1)
) cond33 (
    .clk(cond33_clk),
    .done(cond33_done),
    .in(cond33_in),
    .out(cond33_out),
    .reset(cond33_reset),
    .write_en(cond33_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire33 (
    .in(cond_wire33_in),
    .out(cond_wire33_out)
);
std_reg # (
    .WIDTH(1)
) cond34 (
    .clk(cond34_clk),
    .done(cond34_done),
    .in(cond34_in),
    .out(cond34_out),
    .reset(cond34_reset),
    .write_en(cond34_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire34 (
    .in(cond_wire34_in),
    .out(cond_wire34_out)
);
std_reg # (
    .WIDTH(1)
) cond35 (
    .clk(cond35_clk),
    .done(cond35_done),
    .in(cond35_in),
    .out(cond35_out),
    .reset(cond35_reset),
    .write_en(cond35_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire35 (
    .in(cond_wire35_in),
    .out(cond_wire35_out)
);
std_reg # (
    .WIDTH(1)
) cond36 (
    .clk(cond36_clk),
    .done(cond36_done),
    .in(cond36_in),
    .out(cond36_out),
    .reset(cond36_reset),
    .write_en(cond36_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire36 (
    .in(cond_wire36_in),
    .out(cond_wire36_out)
);
std_reg # (
    .WIDTH(1)
) cond37 (
    .clk(cond37_clk),
    .done(cond37_done),
    .in(cond37_in),
    .out(cond37_out),
    .reset(cond37_reset),
    .write_en(cond37_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire37 (
    .in(cond_wire37_in),
    .out(cond_wire37_out)
);
std_reg # (
    .WIDTH(1)
) cond38 (
    .clk(cond38_clk),
    .done(cond38_done),
    .in(cond38_in),
    .out(cond38_out),
    .reset(cond38_reset),
    .write_en(cond38_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire38 (
    .in(cond_wire38_in),
    .out(cond_wire38_out)
);
std_reg # (
    .WIDTH(1)
) cond39 (
    .clk(cond39_clk),
    .done(cond39_done),
    .in(cond39_in),
    .out(cond39_out),
    .reset(cond39_reset),
    .write_en(cond39_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire39 (
    .in(cond_wire39_in),
    .out(cond_wire39_out)
);
std_reg # (
    .WIDTH(1)
) cond40 (
    .clk(cond40_clk),
    .done(cond40_done),
    .in(cond40_in),
    .out(cond40_out),
    .reset(cond40_reset),
    .write_en(cond40_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire40 (
    .in(cond_wire40_in),
    .out(cond_wire40_out)
);
std_reg # (
    .WIDTH(1)
) cond41 (
    .clk(cond41_clk),
    .done(cond41_done),
    .in(cond41_in),
    .out(cond41_out),
    .reset(cond41_reset),
    .write_en(cond41_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire41 (
    .in(cond_wire41_in),
    .out(cond_wire41_out)
);
std_reg # (
    .WIDTH(1)
) cond42 (
    .clk(cond42_clk),
    .done(cond42_done),
    .in(cond42_in),
    .out(cond42_out),
    .reset(cond42_reset),
    .write_en(cond42_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire42 (
    .in(cond_wire42_in),
    .out(cond_wire42_out)
);
std_reg # (
    .WIDTH(1)
) cond43 (
    .clk(cond43_clk),
    .done(cond43_done),
    .in(cond43_in),
    .out(cond43_out),
    .reset(cond43_reset),
    .write_en(cond43_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire43 (
    .in(cond_wire43_in),
    .out(cond_wire43_out)
);
std_reg # (
    .WIDTH(1)
) cond44 (
    .clk(cond44_clk),
    .done(cond44_done),
    .in(cond44_in),
    .out(cond44_out),
    .reset(cond44_reset),
    .write_en(cond44_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire44 (
    .in(cond_wire44_in),
    .out(cond_wire44_out)
);
std_reg # (
    .WIDTH(1)
) cond45 (
    .clk(cond45_clk),
    .done(cond45_done),
    .in(cond45_in),
    .out(cond45_out),
    .reset(cond45_reset),
    .write_en(cond45_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire45 (
    .in(cond_wire45_in),
    .out(cond_wire45_out)
);
std_reg # (
    .WIDTH(1)
) cond46 (
    .clk(cond46_clk),
    .done(cond46_done),
    .in(cond46_in),
    .out(cond46_out),
    .reset(cond46_reset),
    .write_en(cond46_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire46 (
    .in(cond_wire46_in),
    .out(cond_wire46_out)
);
std_reg # (
    .WIDTH(1)
) cond47 (
    .clk(cond47_clk),
    .done(cond47_done),
    .in(cond47_in),
    .out(cond47_out),
    .reset(cond47_reset),
    .write_en(cond47_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire47 (
    .in(cond_wire47_in),
    .out(cond_wire47_out)
);
std_reg # (
    .WIDTH(1)
) cond48 (
    .clk(cond48_clk),
    .done(cond48_done),
    .in(cond48_in),
    .out(cond48_out),
    .reset(cond48_reset),
    .write_en(cond48_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire48 (
    .in(cond_wire48_in),
    .out(cond_wire48_out)
);
std_reg # (
    .WIDTH(1)
) cond49 (
    .clk(cond49_clk),
    .done(cond49_done),
    .in(cond49_in),
    .out(cond49_out),
    .reset(cond49_reset),
    .write_en(cond49_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire49 (
    .in(cond_wire49_in),
    .out(cond_wire49_out)
);
std_reg # (
    .WIDTH(1)
) cond50 (
    .clk(cond50_clk),
    .done(cond50_done),
    .in(cond50_in),
    .out(cond50_out),
    .reset(cond50_reset),
    .write_en(cond50_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire50 (
    .in(cond_wire50_in),
    .out(cond_wire50_out)
);
std_reg # (
    .WIDTH(1)
) cond51 (
    .clk(cond51_clk),
    .done(cond51_done),
    .in(cond51_in),
    .out(cond51_out),
    .reset(cond51_reset),
    .write_en(cond51_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire51 (
    .in(cond_wire51_in),
    .out(cond_wire51_out)
);
std_reg # (
    .WIDTH(1)
) cond52 (
    .clk(cond52_clk),
    .done(cond52_done),
    .in(cond52_in),
    .out(cond52_out),
    .reset(cond52_reset),
    .write_en(cond52_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire52 (
    .in(cond_wire52_in),
    .out(cond_wire52_out)
);
std_reg # (
    .WIDTH(1)
) cond53 (
    .clk(cond53_clk),
    .done(cond53_done),
    .in(cond53_in),
    .out(cond53_out),
    .reset(cond53_reset),
    .write_en(cond53_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire53 (
    .in(cond_wire53_in),
    .out(cond_wire53_out)
);
std_reg # (
    .WIDTH(1)
) cond54 (
    .clk(cond54_clk),
    .done(cond54_done),
    .in(cond54_in),
    .out(cond54_out),
    .reset(cond54_reset),
    .write_en(cond54_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire54 (
    .in(cond_wire54_in),
    .out(cond_wire54_out)
);
std_reg # (
    .WIDTH(1)
) cond55 (
    .clk(cond55_clk),
    .done(cond55_done),
    .in(cond55_in),
    .out(cond55_out),
    .reset(cond55_reset),
    .write_en(cond55_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire55 (
    .in(cond_wire55_in),
    .out(cond_wire55_out)
);
std_reg # (
    .WIDTH(1)
) cond56 (
    .clk(cond56_clk),
    .done(cond56_done),
    .in(cond56_in),
    .out(cond56_out),
    .reset(cond56_reset),
    .write_en(cond56_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire56 (
    .in(cond_wire56_in),
    .out(cond_wire56_out)
);
std_reg # (
    .WIDTH(1)
) cond57 (
    .clk(cond57_clk),
    .done(cond57_done),
    .in(cond57_in),
    .out(cond57_out),
    .reset(cond57_reset),
    .write_en(cond57_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire57 (
    .in(cond_wire57_in),
    .out(cond_wire57_out)
);
std_reg # (
    .WIDTH(1)
) cond58 (
    .clk(cond58_clk),
    .done(cond58_done),
    .in(cond58_in),
    .out(cond58_out),
    .reset(cond58_reset),
    .write_en(cond58_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire58 (
    .in(cond_wire58_in),
    .out(cond_wire58_out)
);
std_reg # (
    .WIDTH(1)
) cond59 (
    .clk(cond59_clk),
    .done(cond59_done),
    .in(cond59_in),
    .out(cond59_out),
    .reset(cond59_reset),
    .write_en(cond59_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire59 (
    .in(cond_wire59_in),
    .out(cond_wire59_out)
);
std_reg # (
    .WIDTH(1)
) cond60 (
    .clk(cond60_clk),
    .done(cond60_done),
    .in(cond60_in),
    .out(cond60_out),
    .reset(cond60_reset),
    .write_en(cond60_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire60 (
    .in(cond_wire60_in),
    .out(cond_wire60_out)
);
std_reg # (
    .WIDTH(1)
) cond61 (
    .clk(cond61_clk),
    .done(cond61_done),
    .in(cond61_in),
    .out(cond61_out),
    .reset(cond61_reset),
    .write_en(cond61_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire61 (
    .in(cond_wire61_in),
    .out(cond_wire61_out)
);
std_reg # (
    .WIDTH(1)
) cond62 (
    .clk(cond62_clk),
    .done(cond62_done),
    .in(cond62_in),
    .out(cond62_out),
    .reset(cond62_reset),
    .write_en(cond62_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire62 (
    .in(cond_wire62_in),
    .out(cond_wire62_out)
);
std_reg # (
    .WIDTH(1)
) cond63 (
    .clk(cond63_clk),
    .done(cond63_done),
    .in(cond63_in),
    .out(cond63_out),
    .reset(cond63_reset),
    .write_en(cond63_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire63 (
    .in(cond_wire63_in),
    .out(cond_wire63_out)
);
std_reg # (
    .WIDTH(1)
) cond64 (
    .clk(cond64_clk),
    .done(cond64_done),
    .in(cond64_in),
    .out(cond64_out),
    .reset(cond64_reset),
    .write_en(cond64_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire64 (
    .in(cond_wire64_in),
    .out(cond_wire64_out)
);
std_reg # (
    .WIDTH(1)
) cond65 (
    .clk(cond65_clk),
    .done(cond65_done),
    .in(cond65_in),
    .out(cond65_out),
    .reset(cond65_reset),
    .write_en(cond65_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire65 (
    .in(cond_wire65_in),
    .out(cond_wire65_out)
);
std_reg # (
    .WIDTH(1)
) cond66 (
    .clk(cond66_clk),
    .done(cond66_done),
    .in(cond66_in),
    .out(cond66_out),
    .reset(cond66_reset),
    .write_en(cond66_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire66 (
    .in(cond_wire66_in),
    .out(cond_wire66_out)
);
std_reg # (
    .WIDTH(1)
) cond67 (
    .clk(cond67_clk),
    .done(cond67_done),
    .in(cond67_in),
    .out(cond67_out),
    .reset(cond67_reset),
    .write_en(cond67_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire67 (
    .in(cond_wire67_in),
    .out(cond_wire67_out)
);
std_reg # (
    .WIDTH(1)
) cond68 (
    .clk(cond68_clk),
    .done(cond68_done),
    .in(cond68_in),
    .out(cond68_out),
    .reset(cond68_reset),
    .write_en(cond68_write_en)
);
std_wire # (
    .WIDTH(1)
) cond_wire68 (
    .in(cond_wire68_in),
    .out(cond_wire68_out)
);
std_reg # (
    .WIDTH(1)
) fsm (
    .clk(fsm_clk),
    .done(fsm_done),
    .in(fsm_in),
    .out(fsm_out),
    .reset(fsm_reset),
    .write_en(fsm_write_en)
);
std_reg # (
    .WIDTH(5)
) fsm0 (
    .clk(fsm0_clk),
    .done(fsm0_done),
    .in(fsm0_in),
    .out(fsm0_out),
    .reset(fsm0_reset),
    .write_en(fsm0_write_en)
);
undef # (
    .WIDTH(1)
) ud (
    .out(ud_out)
);
std_add # (
    .WIDTH(5)
) adder (
    .left(adder_left),
    .out(adder_out),
    .right(adder_right)
);
undef # (
    .WIDTH(1)
) ud0 (
    .out(ud0_out)
);
std_add # (
    .WIDTH(1)
) adder0 (
    .left(adder0_left),
    .out(adder0_out),
    .right(adder0_right)
);
std_reg # (
    .WIDTH(1)
) signal_reg (
    .clk(signal_reg_clk),
    .done(signal_reg_done),
    .in(signal_reg_in),
    .out(signal_reg_out),
    .reset(signal_reg_reset),
    .write_en(signal_reg_write_en)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_seq_go (
    .in(early_reset_static_seq_go_in),
    .out(early_reset_static_seq_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_seq_done (
    .in(early_reset_static_seq_done_in),
    .out(early_reset_static_seq_done_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par0_go (
    .in(early_reset_static_par0_go_in),
    .out(early_reset_static_par0_go_out)
);
std_wire # (
    .WIDTH(1)
) early_reset_static_par0_done (
    .in(early_reset_static_par0_done_in),
    .out(early_reset_static_par0_done_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_seq_go (
    .in(wrapper_early_reset_static_seq_go_in),
    .out(wrapper_early_reset_static_seq_go_out)
);
std_wire # (
    .WIDTH(1)
) wrapper_early_reset_static_seq_done (
    .in(wrapper_early_reset_static_seq_done_in),
    .out(wrapper_early_reset_static_seq_done_out)
);
wire _guard0 = 1;
wire _guard1 = cond_wire14_out;
wire _guard2 = early_reset_static_par0_go_out;
wire _guard3 = _guard1 & _guard2;
wire _guard4 = cond_wire14_out;
wire _guard5 = early_reset_static_par0_go_out;
wire _guard6 = _guard4 & _guard5;
wire _guard7 = cond_wire19_out;
wire _guard8 = early_reset_static_par0_go_out;
wire _guard9 = _guard7 & _guard8;
wire _guard10 = cond_wire19_out;
wire _guard11 = early_reset_static_par0_go_out;
wire _guard12 = _guard10 & _guard11;
wire _guard13 = fsm0_out == 5'd0;
wire _guard14 = early_reset_static_seq_go_out;
wire _guard15 = _guard13 & _guard14;
wire _guard16 = early_reset_static_par0_go_out;
wire _guard17 = _guard15 | _guard16;
wire _guard18 = early_reset_static_par0_go_out;
wire _guard19 = fsm0_out == 5'd0;
wire _guard20 = early_reset_static_seq_go_out;
wire _guard21 = _guard19 & _guard20;
wire _guard22 = fsm0_out == 5'd0;
wire _guard23 = early_reset_static_seq_go_out;
wire _guard24 = _guard22 & _guard23;
wire _guard25 = early_reset_static_par0_go_out;
wire _guard26 = _guard24 | _guard25;
wire _guard27 = fsm0_out == 5'd0;
wire _guard28 = early_reset_static_seq_go_out;
wire _guard29 = _guard27 & _guard28;
wire _guard30 = early_reset_static_par0_go_out;
wire _guard31 = early_reset_static_par0_go_out;
wire _guard32 = early_reset_static_par0_go_out;
wire _guard33 = early_reset_static_par0_go_out;
wire _guard34 = early_reset_static_par0_go_out;
wire _guard35 = ~_guard0;
wire _guard36 = early_reset_static_par0_go_out;
wire _guard37 = _guard35 & _guard36;
wire _guard38 = early_reset_static_par0_go_out;
wire _guard39 = ~_guard0;
wire _guard40 = early_reset_static_par0_go_out;
wire _guard41 = _guard39 & _guard40;
wire _guard42 = early_reset_static_par0_go_out;
wire _guard43 = early_reset_static_par0_go_out;
wire _guard44 = ~_guard0;
wire _guard45 = early_reset_static_par0_go_out;
wire _guard46 = _guard44 & _guard45;
wire _guard47 = early_reset_static_par0_go_out;
wire _guard48 = ~_guard0;
wire _guard49 = early_reset_static_par0_go_out;
wire _guard50 = _guard48 & _guard49;
wire _guard51 = ~_guard0;
wire _guard52 = early_reset_static_par0_go_out;
wire _guard53 = _guard51 & _guard52;
wire _guard54 = early_reset_static_par0_go_out;
wire _guard55 = early_reset_static_par0_go_out;
wire _guard56 = early_reset_static_par0_go_out;
wire _guard57 = early_reset_static_par0_go_out;
wire _guard58 = ~_guard0;
wire _guard59 = early_reset_static_par0_go_out;
wire _guard60 = _guard58 & _guard59;
wire _guard61 = early_reset_static_par0_go_out;
wire _guard62 = early_reset_static_par0_go_out;
wire _guard63 = cond_wire11_out;
wire _guard64 = early_reset_static_par0_go_out;
wire _guard65 = _guard63 & _guard64;
wire _guard66 = cond_wire11_out;
wire _guard67 = early_reset_static_par0_go_out;
wire _guard68 = _guard66 & _guard67;
wire _guard69 = cond_wire1_out;
wire _guard70 = early_reset_static_par0_go_out;
wire _guard71 = _guard69 & _guard70;
wire _guard72 = cond_wire1_out;
wire _guard73 = early_reset_static_par0_go_out;
wire _guard74 = _guard72 & _guard73;
wire _guard75 = cond_wire30_out;
wire _guard76 = early_reset_static_par0_go_out;
wire _guard77 = _guard75 & _guard76;
wire _guard78 = cond_wire28_out;
wire _guard79 = early_reset_static_par0_go_out;
wire _guard80 = _guard78 & _guard79;
wire _guard81 = fsm_out == 1'd0;
wire _guard82 = cond_wire28_out;
wire _guard83 = _guard81 & _guard82;
wire _guard84 = fsm_out == 1'd0;
wire _guard85 = _guard83 & _guard84;
wire _guard86 = fsm_out == 1'd0;
wire _guard87 = cond_wire30_out;
wire _guard88 = _guard86 & _guard87;
wire _guard89 = fsm_out == 1'd0;
wire _guard90 = _guard88 & _guard89;
wire _guard91 = _guard85 | _guard90;
wire _guard92 = early_reset_static_par0_go_out;
wire _guard93 = _guard91 & _guard92;
wire _guard94 = fsm_out == 1'd0;
wire _guard95 = cond_wire28_out;
wire _guard96 = _guard94 & _guard95;
wire _guard97 = fsm_out == 1'd0;
wire _guard98 = _guard96 & _guard97;
wire _guard99 = fsm_out == 1'd0;
wire _guard100 = cond_wire30_out;
wire _guard101 = _guard99 & _guard100;
wire _guard102 = fsm_out == 1'd0;
wire _guard103 = _guard101 & _guard102;
wire _guard104 = _guard98 | _guard103;
wire _guard105 = early_reset_static_par0_go_out;
wire _guard106 = _guard104 & _guard105;
wire _guard107 = fsm_out == 1'd0;
wire _guard108 = cond_wire28_out;
wire _guard109 = _guard107 & _guard108;
wire _guard110 = fsm_out == 1'd0;
wire _guard111 = _guard109 & _guard110;
wire _guard112 = fsm_out == 1'd0;
wire _guard113 = cond_wire30_out;
wire _guard114 = _guard112 & _guard113;
wire _guard115 = fsm_out == 1'd0;
wire _guard116 = _guard114 & _guard115;
wire _guard117 = _guard111 | _guard116;
wire _guard118 = early_reset_static_par0_go_out;
wire _guard119 = _guard117 & _guard118;
wire _guard120 = cond_wire34_out;
wire _guard121 = early_reset_static_par0_go_out;
wire _guard122 = _guard120 & _guard121;
wire _guard123 = cond_wire32_out;
wire _guard124 = early_reset_static_par0_go_out;
wire _guard125 = _guard123 & _guard124;
wire _guard126 = fsm_out == 1'd0;
wire _guard127 = cond_wire32_out;
wire _guard128 = _guard126 & _guard127;
wire _guard129 = fsm_out == 1'd0;
wire _guard130 = _guard128 & _guard129;
wire _guard131 = fsm_out == 1'd0;
wire _guard132 = cond_wire34_out;
wire _guard133 = _guard131 & _guard132;
wire _guard134 = fsm_out == 1'd0;
wire _guard135 = _guard133 & _guard134;
wire _guard136 = _guard130 | _guard135;
wire _guard137 = early_reset_static_par0_go_out;
wire _guard138 = _guard136 & _guard137;
wire _guard139 = fsm_out == 1'd0;
wire _guard140 = cond_wire32_out;
wire _guard141 = _guard139 & _guard140;
wire _guard142 = fsm_out == 1'd0;
wire _guard143 = _guard141 & _guard142;
wire _guard144 = fsm_out == 1'd0;
wire _guard145 = cond_wire34_out;
wire _guard146 = _guard144 & _guard145;
wire _guard147 = fsm_out == 1'd0;
wire _guard148 = _guard146 & _guard147;
wire _guard149 = _guard143 | _guard148;
wire _guard150 = early_reset_static_par0_go_out;
wire _guard151 = _guard149 & _guard150;
wire _guard152 = fsm_out == 1'd0;
wire _guard153 = cond_wire32_out;
wire _guard154 = _guard152 & _guard153;
wire _guard155 = fsm_out == 1'd0;
wire _guard156 = _guard154 & _guard155;
wire _guard157 = fsm_out == 1'd0;
wire _guard158 = cond_wire34_out;
wire _guard159 = _guard157 & _guard158;
wire _guard160 = fsm_out == 1'd0;
wire _guard161 = _guard159 & _guard160;
wire _guard162 = _guard156 | _guard161;
wire _guard163 = early_reset_static_par0_go_out;
wire _guard164 = _guard162 & _guard163;
wire _guard165 = cond_wire29_out;
wire _guard166 = early_reset_static_par0_go_out;
wire _guard167 = _guard165 & _guard166;
wire _guard168 = cond_wire29_out;
wire _guard169 = early_reset_static_par0_go_out;
wire _guard170 = _guard168 & _guard169;
wire _guard171 = fsm0_out == 5'd0;
wire _guard172 = early_reset_static_seq_go_out;
wire _guard173 = _guard171 & _guard172;
wire _guard174 = cond_wire53_out;
wire _guard175 = early_reset_static_par0_go_out;
wire _guard176 = _guard174 & _guard175;
wire _guard177 = _guard173 | _guard176;
wire _guard178 = cond_wire53_out;
wire _guard179 = early_reset_static_par0_go_out;
wire _guard180 = _guard178 & _guard179;
wire _guard181 = fsm0_out == 5'd0;
wire _guard182 = early_reset_static_seq_go_out;
wire _guard183 = _guard181 & _guard182;
wire _guard184 = early_reset_static_par0_go_out;
wire _guard185 = early_reset_static_par0_go_out;
wire _guard186 = early_reset_static_par0_go_out;
wire _guard187 = early_reset_static_par0_go_out;
wire _guard188 = early_reset_static_par0_go_out;
wire _guard189 = early_reset_static_par0_go_out;
wire _guard190 = fsm0_out == 5'd0;
wire _guard191 = early_reset_static_seq_go_out;
wire _guard192 = _guard190 & _guard191;
wire _guard193 = early_reset_static_par0_go_out;
wire _guard194 = _guard192 | _guard193;
wire _guard195 = early_reset_static_par0_go_out;
wire _guard196 = fsm0_out == 5'd0;
wire _guard197 = early_reset_static_seq_go_out;
wire _guard198 = _guard196 & _guard197;
wire _guard199 = fsm0_out == 5'd0;
wire _guard200 = early_reset_static_seq_go_out;
wire _guard201 = _guard199 & _guard200;
wire _guard202 = early_reset_static_par0_go_out;
wire _guard203 = _guard201 | _guard202;
wire _guard204 = early_reset_static_par0_go_out;
wire _guard205 = fsm0_out == 5'd0;
wire _guard206 = early_reset_static_seq_go_out;
wire _guard207 = _guard205 & _guard206;
wire _guard208 = wrapper_early_reset_static_seq_done_out;
wire _guard209 = cond_wire9_out;
wire _guard210 = early_reset_static_par0_go_out;
wire _guard211 = _guard209 & _guard210;
wire _guard212 = cond_wire_out;
wire _guard213 = early_reset_static_par0_go_out;
wire _guard214 = _guard212 & _guard213;
wire _guard215 = cond_wire31_out;
wire _guard216 = early_reset_static_par0_go_out;
wire _guard217 = _guard215 & _guard216;
wire _guard218 = cond_wire23_out;
wire _guard219 = early_reset_static_par0_go_out;
wire _guard220 = _guard218 & _guard219;
wire _guard221 = cond_wire27_out;
wire _guard222 = early_reset_static_par0_go_out;
wire _guard223 = _guard221 & _guard222;
wire _guard224 = cond_wire35_out;
wire _guard225 = early_reset_static_par0_go_out;
wire _guard226 = _guard224 & _guard225;
wire _guard227 = cond_wire8_out;
wire _guard228 = early_reset_static_par0_go_out;
wire _guard229 = _guard227 & _guard228;
wire _guard230 = cond_wire18_out;
wire _guard231 = early_reset_static_par0_go_out;
wire _guard232 = _guard230 & _guard231;
wire _guard233 = cond_wire13_out;
wire _guard234 = early_reset_static_par0_go_out;
wire _guard235 = _guard233 & _guard234;
wire _guard236 = cond_wire3_out;
wire _guard237 = early_reset_static_par0_go_out;
wire _guard238 = _guard236 & _guard237;
wire _guard239 = cond_wire65_out;
wire _guard240 = early_reset_static_par0_go_out;
wire _guard241 = _guard239 & _guard240;
wire _guard242 = cond_wire57_out;
wire _guard243 = early_reset_static_par0_go_out;
wire _guard244 = _guard242 & _guard243;
wire _guard245 = cond_wire61_out;
wire _guard246 = early_reset_static_par0_go_out;
wire _guard247 = _guard245 & _guard246;
wire _guard248 = cond_wire68_out;
wire _guard249 = early_reset_static_par0_go_out;
wire _guard250 = _guard248 & _guard249;
wire _guard251 = cond_wire19_out;
wire _guard252 = early_reset_static_par0_go_out;
wire _guard253 = _guard251 & _guard252;
wire _guard254 = cond_wire53_out;
wire _guard255 = early_reset_static_par0_go_out;
wire _guard256 = _guard254 & _guard255;
wire _guard257 = cond_wire44_out;
wire _guard258 = early_reset_static_par0_go_out;
wire _guard259 = _guard257 & _guard258;
wire _guard260 = cond_wire52_out;
wire _guard261 = early_reset_static_par0_go_out;
wire _guard262 = _guard260 & _guard261;
wire _guard263 = cond_wire40_out;
wire _guard264 = early_reset_static_par0_go_out;
wire _guard265 = _guard263 & _guard264;
wire _guard266 = cond_wire48_out;
wire _guard267 = early_reset_static_par0_go_out;
wire _guard268 = _guard266 & _guard267;
wire _guard269 = cond_wire31_out;
wire _guard270 = early_reset_static_par0_go_out;
wire _guard271 = _guard269 & _guard270;
wire _guard272 = cond_wire35_out;
wire _guard273 = early_reset_static_par0_go_out;
wire _guard274 = _guard272 & _guard273;
wire _guard275 = cond_wire23_out;
wire _guard276 = early_reset_static_par0_go_out;
wire _guard277 = _guard275 & _guard276;
wire _guard278 = cond_wire27_out;
wire _guard279 = early_reset_static_par0_go_out;
wire _guard280 = _guard278 & _guard279;
wire _guard281 = fsm_out == 1'd0;
wire _guard282 = cond_wire23_out;
wire _guard283 = _guard281 & _guard282;
wire _guard284 = fsm_out == 1'd0;
wire _guard285 = _guard283 & _guard284;
wire _guard286 = fsm_out == 1'd0;
wire _guard287 = cond_wire27_out;
wire _guard288 = _guard286 & _guard287;
wire _guard289 = fsm_out == 1'd0;
wire _guard290 = _guard288 & _guard289;
wire _guard291 = _guard285 | _guard290;
wire _guard292 = fsm_out == 1'd0;
wire _guard293 = cond_wire31_out;
wire _guard294 = _guard292 & _guard293;
wire _guard295 = fsm_out == 1'd0;
wire _guard296 = _guard294 & _guard295;
wire _guard297 = _guard291 | _guard296;
wire _guard298 = fsm_out == 1'd0;
wire _guard299 = cond_wire35_out;
wire _guard300 = _guard298 & _guard299;
wire _guard301 = fsm_out == 1'd0;
wire _guard302 = _guard300 & _guard301;
wire _guard303 = _guard297 | _guard302;
wire _guard304 = early_reset_static_par0_go_out;
wire _guard305 = _guard303 & _guard304;
wire _guard306 = cond_wire_out;
wire _guard307 = early_reset_static_par0_go_out;
wire _guard308 = _guard306 & _guard307;
wire _guard309 = cond_wire4_out;
wire _guard310 = early_reset_static_par0_go_out;
wire _guard311 = _guard309 & _guard310;
wire _guard312 = fsm_out == 1'd0;
wire _guard313 = cond_wire3_out;
wire _guard314 = _guard312 & _guard313;
wire _guard315 = fsm_out == 1'd0;
wire _guard316 = _guard314 & _guard315;
wire _guard317 = fsm_out == 1'd0;
wire _guard318 = cond_wire8_out;
wire _guard319 = _guard317 & _guard318;
wire _guard320 = fsm_out == 1'd0;
wire _guard321 = _guard319 & _guard320;
wire _guard322 = _guard316 | _guard321;
wire _guard323 = fsm_out == 1'd0;
wire _guard324 = cond_wire13_out;
wire _guard325 = _guard323 & _guard324;
wire _guard326 = fsm_out == 1'd0;
wire _guard327 = _guard325 & _guard326;
wire _guard328 = _guard322 | _guard327;
wire _guard329 = fsm_out == 1'd0;
wire _guard330 = cond_wire18_out;
wire _guard331 = _guard329 & _guard330;
wire _guard332 = fsm_out == 1'd0;
wire _guard333 = _guard331 & _guard332;
wire _guard334 = _guard328 | _guard333;
wire _guard335 = early_reset_static_par0_go_out;
wire _guard336 = _guard334 & _guard335;
wire _guard337 = fsm_out == 1'd0;
wire _guard338 = cond_wire40_out;
wire _guard339 = _guard337 & _guard338;
wire _guard340 = fsm_out == 1'd0;
wire _guard341 = _guard339 & _guard340;
wire _guard342 = fsm_out == 1'd0;
wire _guard343 = cond_wire44_out;
wire _guard344 = _guard342 & _guard343;
wire _guard345 = fsm_out == 1'd0;
wire _guard346 = _guard344 & _guard345;
wire _guard347 = _guard341 | _guard346;
wire _guard348 = fsm_out == 1'd0;
wire _guard349 = cond_wire48_out;
wire _guard350 = _guard348 & _guard349;
wire _guard351 = fsm_out == 1'd0;
wire _guard352 = _guard350 & _guard351;
wire _guard353 = _guard347 | _guard352;
wire _guard354 = fsm_out == 1'd0;
wire _guard355 = cond_wire52_out;
wire _guard356 = _guard354 & _guard355;
wire _guard357 = fsm_out == 1'd0;
wire _guard358 = _guard356 & _guard357;
wire _guard359 = _guard353 | _guard358;
wire _guard360 = early_reset_static_par0_go_out;
wire _guard361 = _guard359 & _guard360;
wire _guard362 = fsm_out == 1'd0;
wire _guard363 = cond_wire57_out;
wire _guard364 = _guard362 & _guard363;
wire _guard365 = fsm_out == 1'd0;
wire _guard366 = _guard364 & _guard365;
wire _guard367 = fsm_out == 1'd0;
wire _guard368 = cond_wire61_out;
wire _guard369 = _guard367 & _guard368;
wire _guard370 = fsm_out == 1'd0;
wire _guard371 = _guard369 & _guard370;
wire _guard372 = _guard366 | _guard371;
wire _guard373 = fsm_out == 1'd0;
wire _guard374 = cond_wire65_out;
wire _guard375 = _guard373 & _guard374;
wire _guard376 = fsm_out == 1'd0;
wire _guard377 = _guard375 & _guard376;
wire _guard378 = _guard372 | _guard377;
wire _guard379 = fsm_out == 1'd0;
wire _guard380 = cond_wire68_out;
wire _guard381 = _guard379 & _guard380;
wire _guard382 = fsm_out == 1'd0;
wire _guard383 = _guard381 & _guard382;
wire _guard384 = _guard378 | _guard383;
wire _guard385 = early_reset_static_par0_go_out;
wire _guard386 = _guard384 & _guard385;
wire _guard387 = cond_wire36_out;
wire _guard388 = early_reset_static_par0_go_out;
wire _guard389 = _guard387 & _guard388;
wire _guard390 = cond_wire13_out;
wire _guard391 = early_reset_static_par0_go_out;
wire _guard392 = _guard390 & _guard391;
wire _guard393 = cond_wire3_out;
wire _guard394 = early_reset_static_par0_go_out;
wire _guard395 = _guard393 & _guard394;
wire _guard396 = cond_wire8_out;
wire _guard397 = early_reset_static_par0_go_out;
wire _guard398 = _guard396 & _guard397;
wire _guard399 = cond_wire18_out;
wire _guard400 = early_reset_static_par0_go_out;
wire _guard401 = _guard399 & _guard400;
wire _guard402 = cond_wire65_out;
wire _guard403 = early_reset_static_par0_go_out;
wire _guard404 = _guard402 & _guard403;
wire _guard405 = cond_wire57_out;
wire _guard406 = early_reset_static_par0_go_out;
wire _guard407 = _guard405 & _guard406;
wire _guard408 = cond_wire61_out;
wire _guard409 = early_reset_static_par0_go_out;
wire _guard410 = _guard408 & _guard409;
wire _guard411 = cond_wire68_out;
wire _guard412 = early_reset_static_par0_go_out;
wire _guard413 = _guard411 & _guard412;
wire _guard414 = cond_wire14_out;
wire _guard415 = early_reset_static_par0_go_out;
wire _guard416 = _guard414 & _guard415;
wire _guard417 = cond_wire48_out;
wire _guard418 = early_reset_static_par0_go_out;
wire _guard419 = _guard417 & _guard418;
wire _guard420 = cond_wire40_out;
wire _guard421 = early_reset_static_par0_go_out;
wire _guard422 = _guard420 & _guard421;
wire _guard423 = cond_wire44_out;
wire _guard424 = early_reset_static_par0_go_out;
wire _guard425 = _guard423 & _guard424;
wire _guard426 = cond_wire52_out;
wire _guard427 = early_reset_static_par0_go_out;
wire _guard428 = _guard426 & _guard427;
wire _guard429 = early_reset_static_par0_go_out;
wire _guard430 = ~_guard0;
wire _guard431 = early_reset_static_par0_go_out;
wire _guard432 = _guard430 & _guard431;
wire _guard433 = early_reset_static_par0_go_out;
wire _guard434 = ~_guard0;
wire _guard435 = early_reset_static_par0_go_out;
wire _guard436 = _guard434 & _guard435;
wire _guard437 = early_reset_static_par0_go_out;
wire _guard438 = early_reset_static_par0_go_out;
wire _guard439 = ~_guard0;
wire _guard440 = early_reset_static_par0_go_out;
wire _guard441 = _guard439 & _guard440;
wire _guard442 = early_reset_static_par0_go_out;
wire _guard443 = early_reset_static_par0_go_out;
wire _guard444 = ~_guard0;
wire _guard445 = early_reset_static_par0_go_out;
wire _guard446 = _guard444 & _guard445;
wire _guard447 = early_reset_static_par0_go_out;
wire _guard448 = early_reset_static_par0_go_out;
wire _guard449 = early_reset_static_par0_go_out;
wire _guard450 = ~_guard0;
wire _guard451 = early_reset_static_par0_go_out;
wire _guard452 = _guard450 & _guard451;
wire _guard453 = ~_guard0;
wire _guard454 = early_reset_static_par0_go_out;
wire _guard455 = _guard453 & _guard454;
wire _guard456 = early_reset_static_par0_go_out;
wire _guard457 = early_reset_static_par0_go_out;
wire _guard458 = early_reset_static_par0_go_out;
wire _guard459 = early_reset_static_par0_go_out;
wire _guard460 = early_reset_static_par0_go_out;
wire _guard461 = early_reset_static_par0_go_out;
wire _guard462 = fsm_out == 1'd0;
wire _guard463 = early_reset_static_par0_go_out;
wire _guard464 = _guard462 & _guard463;
wire _guard465 = fsm_out != 1'd0;
wire _guard466 = early_reset_static_par0_go_out;
wire _guard467 = _guard465 & _guard466;
wire _guard468 = early_reset_static_seq_go_out;
wire _guard469 = early_reset_static_seq_go_out;
wire _guard470 = fsm0_out >= 5'd1;
wire _guard471 = fsm0_out < 5'd17;
wire _guard472 = _guard470 & _guard471;
wire _guard473 = early_reset_static_seq_go_out;
wire _guard474 = _guard472 & _guard473;
wire _guard475 = fsm0_out == 5'd0;
wire _guard476 = early_reset_static_seq_go_out;
wire _guard477 = _guard475 & _guard476;
wire _guard478 = cond_wire_out;
wire _guard479 = early_reset_static_par0_go_out;
wire _guard480 = _guard478 & _guard479;
wire _guard481 = _guard477 | _guard480;
wire _guard482 = cond_wire_out;
wire _guard483 = early_reset_static_par0_go_out;
wire _guard484 = _guard482 & _guard483;
wire _guard485 = fsm0_out == 5'd0;
wire _guard486 = early_reset_static_seq_go_out;
wire _guard487 = _guard485 & _guard486;
wire _guard488 = fsm0_out == 5'd0;
wire _guard489 = early_reset_static_seq_go_out;
wire _guard490 = _guard488 & _guard489;
wire _guard491 = early_reset_static_par0_go_out;
wire _guard492 = _guard490 | _guard491;
wire _guard493 = early_reset_static_par0_go_out;
wire _guard494 = fsm0_out == 5'd0;
wire _guard495 = early_reset_static_seq_go_out;
wire _guard496 = _guard494 & _guard495;
wire _guard497 = early_reset_static_par0_go_out;
wire _guard498 = early_reset_static_par0_go_out;
wire _guard499 = early_reset_static_par0_go_out;
wire _guard500 = early_reset_static_par0_go_out;
wire _guard501 = fsm0_out == 5'd0;
wire _guard502 = early_reset_static_seq_go_out;
wire _guard503 = _guard501 & _guard502;
wire _guard504 = early_reset_static_par0_go_out;
wire _guard505 = _guard503 | _guard504;
wire _guard506 = fsm0_out == 5'd0;
wire _guard507 = early_reset_static_seq_go_out;
wire _guard508 = _guard506 & _guard507;
wire _guard509 = early_reset_static_par0_go_out;
wire _guard510 = early_reset_static_par0_go_out;
wire _guard511 = early_reset_static_par0_go_out;
wire _guard512 = early_reset_static_par0_go_out;
wire _guard513 = early_reset_static_par0_go_out;
wire _guard514 = ~_guard0;
wire _guard515 = early_reset_static_par0_go_out;
wire _guard516 = _guard514 & _guard515;
wire _guard517 = early_reset_static_par0_go_out;
wire _guard518 = early_reset_static_par0_go_out;
wire _guard519 = early_reset_static_par0_go_out;
wire _guard520 = ~_guard0;
wire _guard521 = early_reset_static_par0_go_out;
wire _guard522 = _guard520 & _guard521;
wire _guard523 = early_reset_static_par0_go_out;
wire _guard524 = ~_guard0;
wire _guard525 = early_reset_static_par0_go_out;
wire _guard526 = _guard524 & _guard525;
wire _guard527 = early_reset_static_par0_go_out;
wire _guard528 = early_reset_static_par0_go_out;
wire _guard529 = early_reset_static_par0_go_out;
wire _guard530 = early_reset_static_par0_go_out;
wire _guard531 = ~_guard0;
wire _guard532 = early_reset_static_par0_go_out;
wire _guard533 = _guard531 & _guard532;
wire _guard534 = ~_guard0;
wire _guard535 = early_reset_static_par0_go_out;
wire _guard536 = _guard534 & _guard535;
wire _guard537 = early_reset_static_par0_go_out;
wire _guard538 = cond_wire7_out;
wire _guard539 = early_reset_static_par0_go_out;
wire _guard540 = _guard538 & _guard539;
wire _guard541 = cond_wire5_out;
wire _guard542 = early_reset_static_par0_go_out;
wire _guard543 = _guard541 & _guard542;
wire _guard544 = fsm_out == 1'd0;
wire _guard545 = cond_wire5_out;
wire _guard546 = _guard544 & _guard545;
wire _guard547 = fsm_out == 1'd0;
wire _guard548 = _guard546 & _guard547;
wire _guard549 = fsm_out == 1'd0;
wire _guard550 = cond_wire7_out;
wire _guard551 = _guard549 & _guard550;
wire _guard552 = fsm_out == 1'd0;
wire _guard553 = _guard551 & _guard552;
wire _guard554 = _guard548 | _guard553;
wire _guard555 = early_reset_static_par0_go_out;
wire _guard556 = _guard554 & _guard555;
wire _guard557 = fsm_out == 1'd0;
wire _guard558 = cond_wire5_out;
wire _guard559 = _guard557 & _guard558;
wire _guard560 = fsm_out == 1'd0;
wire _guard561 = _guard559 & _guard560;
wire _guard562 = fsm_out == 1'd0;
wire _guard563 = cond_wire7_out;
wire _guard564 = _guard562 & _guard563;
wire _guard565 = fsm_out == 1'd0;
wire _guard566 = _guard564 & _guard565;
wire _guard567 = _guard561 | _guard566;
wire _guard568 = early_reset_static_par0_go_out;
wire _guard569 = _guard567 & _guard568;
wire _guard570 = fsm_out == 1'd0;
wire _guard571 = cond_wire5_out;
wire _guard572 = _guard570 & _guard571;
wire _guard573 = fsm_out == 1'd0;
wire _guard574 = _guard572 & _guard573;
wire _guard575 = fsm_out == 1'd0;
wire _guard576 = cond_wire7_out;
wire _guard577 = _guard575 & _guard576;
wire _guard578 = fsm_out == 1'd0;
wire _guard579 = _guard577 & _guard578;
wire _guard580 = _guard574 | _guard579;
wire _guard581 = early_reset_static_par0_go_out;
wire _guard582 = _guard580 & _guard581;
wire _guard583 = cond_wire25_out;
wire _guard584 = early_reset_static_par0_go_out;
wire _guard585 = _guard583 & _guard584;
wire _guard586 = cond_wire25_out;
wire _guard587 = early_reset_static_par0_go_out;
wire _guard588 = _guard586 & _guard587;
wire _guard589 = cond_wire42_out;
wire _guard590 = early_reset_static_par0_go_out;
wire _guard591 = _guard589 & _guard590;
wire _guard592 = cond_wire42_out;
wire _guard593 = early_reset_static_par0_go_out;
wire _guard594 = _guard592 & _guard593;
wire _guard595 = cond_wire53_out;
wire _guard596 = early_reset_static_par0_go_out;
wire _guard597 = _guard595 & _guard596;
wire _guard598 = cond_wire53_out;
wire _guard599 = early_reset_static_par0_go_out;
wire _guard600 = _guard598 & _guard599;
wire _guard601 = early_reset_static_par0_go_out;
wire _guard602 = early_reset_static_par0_go_out;
wire _guard603 = early_reset_static_par0_go_out;
wire _guard604 = early_reset_static_par0_go_out;
wire _guard605 = fsm0_out == 5'd0;
wire _guard606 = early_reset_static_seq_go_out;
wire _guard607 = _guard605 & _guard606;
wire _guard608 = early_reset_static_par0_go_out;
wire _guard609 = _guard607 | _guard608;
wire _guard610 = fsm0_out == 5'd0;
wire _guard611 = early_reset_static_seq_go_out;
wire _guard612 = _guard610 & _guard611;
wire _guard613 = early_reset_static_par0_go_out;
wire _guard614 = early_reset_static_par0_go_out;
wire _guard615 = early_reset_static_par0_go_out;
wire _guard616 = early_reset_static_par0_go_out;
wire _guard617 = early_reset_static_par0_go_out;
wire _guard618 = early_reset_static_par0_go_out;
wire _guard619 = early_reset_static_par0_go_out;
wire _guard620 = early_reset_static_par0_go_out;
wire _guard621 = early_reset_static_par0_go_out;
wire _guard622 = early_reset_static_par0_go_out;
wire _guard623 = early_reset_static_par0_go_out;
wire _guard624 = early_reset_static_par0_go_out;
wire _guard625 = ~_guard0;
wire _guard626 = early_reset_static_par0_go_out;
wire _guard627 = _guard625 & _guard626;
wire _guard628 = early_reset_static_par0_go_out;
wire _guard629 = early_reset_static_par0_go_out;
wire _guard630 = early_reset_static_par0_go_out;
wire _guard631 = ~_guard0;
wire _guard632 = early_reset_static_par0_go_out;
wire _guard633 = _guard631 & _guard632;
wire _guard634 = early_reset_static_par0_go_out;
wire _guard635 = ~_guard0;
wire _guard636 = early_reset_static_par0_go_out;
wire _guard637 = _guard635 & _guard636;
wire _guard638 = early_reset_static_par0_go_out;
wire _guard639 = ~_guard0;
wire _guard640 = early_reset_static_par0_go_out;
wire _guard641 = _guard639 & _guard640;
wire _guard642 = early_reset_static_par0_go_out;
wire _guard643 = early_reset_static_par0_go_out;
wire _guard644 = cond_wire22_out;
wire _guard645 = early_reset_static_par0_go_out;
wire _guard646 = _guard644 & _guard645;
wire _guard647 = cond_wire20_out;
wire _guard648 = early_reset_static_par0_go_out;
wire _guard649 = _guard647 & _guard648;
wire _guard650 = fsm_out == 1'd0;
wire _guard651 = cond_wire20_out;
wire _guard652 = _guard650 & _guard651;
wire _guard653 = fsm_out == 1'd0;
wire _guard654 = _guard652 & _guard653;
wire _guard655 = fsm_out == 1'd0;
wire _guard656 = cond_wire22_out;
wire _guard657 = _guard655 & _guard656;
wire _guard658 = fsm_out == 1'd0;
wire _guard659 = _guard657 & _guard658;
wire _guard660 = _guard654 | _guard659;
wire _guard661 = early_reset_static_par0_go_out;
wire _guard662 = _guard660 & _guard661;
wire _guard663 = fsm_out == 1'd0;
wire _guard664 = cond_wire20_out;
wire _guard665 = _guard663 & _guard664;
wire _guard666 = fsm_out == 1'd0;
wire _guard667 = _guard665 & _guard666;
wire _guard668 = fsm_out == 1'd0;
wire _guard669 = cond_wire22_out;
wire _guard670 = _guard668 & _guard669;
wire _guard671 = fsm_out == 1'd0;
wire _guard672 = _guard670 & _guard671;
wire _guard673 = _guard667 | _guard672;
wire _guard674 = early_reset_static_par0_go_out;
wire _guard675 = _guard673 & _guard674;
wire _guard676 = fsm_out == 1'd0;
wire _guard677 = cond_wire20_out;
wire _guard678 = _guard676 & _guard677;
wire _guard679 = fsm_out == 1'd0;
wire _guard680 = _guard678 & _guard679;
wire _guard681 = fsm_out == 1'd0;
wire _guard682 = cond_wire22_out;
wire _guard683 = _guard681 & _guard682;
wire _guard684 = fsm_out == 1'd0;
wire _guard685 = _guard683 & _guard684;
wire _guard686 = _guard680 | _guard685;
wire _guard687 = early_reset_static_par0_go_out;
wire _guard688 = _guard686 & _guard687;
wire _guard689 = cond_wire19_out;
wire _guard690 = early_reset_static_par0_go_out;
wire _guard691 = _guard689 & _guard690;
wire _guard692 = cond_wire19_out;
wire _guard693 = early_reset_static_par0_go_out;
wire _guard694 = _guard692 & _guard693;
wire _guard695 = cond_wire21_out;
wire _guard696 = early_reset_static_par0_go_out;
wire _guard697 = _guard695 & _guard696;
wire _guard698 = cond_wire21_out;
wire _guard699 = early_reset_static_par0_go_out;
wire _guard700 = _guard698 & _guard699;
wire _guard701 = cond_wire11_out;
wire _guard702 = early_reset_static_par0_go_out;
wire _guard703 = _guard701 & _guard702;
wire _guard704 = cond_wire11_out;
wire _guard705 = early_reset_static_par0_go_out;
wire _guard706 = _guard704 & _guard705;
wire _guard707 = cond_wire36_out;
wire _guard708 = early_reset_static_par0_go_out;
wire _guard709 = _guard707 & _guard708;
wire _guard710 = cond_wire36_out;
wire _guard711 = early_reset_static_par0_go_out;
wire _guard712 = _guard710 & _guard711;
wire _guard713 = cond_wire55_out;
wire _guard714 = early_reset_static_par0_go_out;
wire _guard715 = _guard713 & _guard714;
wire _guard716 = cond_wire55_out;
wire _guard717 = early_reset_static_par0_go_out;
wire _guard718 = _guard716 & _guard717;
wire _guard719 = cond_wire64_out;
wire _guard720 = early_reset_static_par0_go_out;
wire _guard721 = _guard719 & _guard720;
wire _guard722 = cond_wire62_out;
wire _guard723 = early_reset_static_par0_go_out;
wire _guard724 = _guard722 & _guard723;
wire _guard725 = fsm_out == 1'd0;
wire _guard726 = cond_wire62_out;
wire _guard727 = _guard725 & _guard726;
wire _guard728 = fsm_out == 1'd0;
wire _guard729 = _guard727 & _guard728;
wire _guard730 = fsm_out == 1'd0;
wire _guard731 = cond_wire64_out;
wire _guard732 = _guard730 & _guard731;
wire _guard733 = fsm_out == 1'd0;
wire _guard734 = _guard732 & _guard733;
wire _guard735 = _guard729 | _guard734;
wire _guard736 = early_reset_static_par0_go_out;
wire _guard737 = _guard735 & _guard736;
wire _guard738 = fsm_out == 1'd0;
wire _guard739 = cond_wire62_out;
wire _guard740 = _guard738 & _guard739;
wire _guard741 = fsm_out == 1'd0;
wire _guard742 = _guard740 & _guard741;
wire _guard743 = fsm_out == 1'd0;
wire _guard744 = cond_wire64_out;
wire _guard745 = _guard743 & _guard744;
wire _guard746 = fsm_out == 1'd0;
wire _guard747 = _guard745 & _guard746;
wire _guard748 = _guard742 | _guard747;
wire _guard749 = early_reset_static_par0_go_out;
wire _guard750 = _guard748 & _guard749;
wire _guard751 = fsm_out == 1'd0;
wire _guard752 = cond_wire62_out;
wire _guard753 = _guard751 & _guard752;
wire _guard754 = fsm_out == 1'd0;
wire _guard755 = _guard753 & _guard754;
wire _guard756 = fsm_out == 1'd0;
wire _guard757 = cond_wire64_out;
wire _guard758 = _guard756 & _guard757;
wire _guard759 = fsm_out == 1'd0;
wire _guard760 = _guard758 & _guard759;
wire _guard761 = _guard755 | _guard760;
wire _guard762 = early_reset_static_par0_go_out;
wire _guard763 = _guard761 & _guard762;
wire _guard764 = fsm0_out == 5'd0;
wire _guard765 = early_reset_static_seq_go_out;
wire _guard766 = _guard764 & _guard765;
wire _guard767 = cond_wire4_out;
wire _guard768 = early_reset_static_par0_go_out;
wire _guard769 = _guard767 & _guard768;
wire _guard770 = _guard766 | _guard769;
wire _guard771 = cond_wire4_out;
wire _guard772 = early_reset_static_par0_go_out;
wire _guard773 = _guard771 & _guard772;
wire _guard774 = fsm0_out == 5'd0;
wire _guard775 = early_reset_static_seq_go_out;
wire _guard776 = _guard774 & _guard775;
wire _guard777 = early_reset_static_par0_go_out;
wire _guard778 = early_reset_static_par0_go_out;
wire _guard779 = early_reset_static_par0_go_out;
wire _guard780 = ~_guard0;
wire _guard781 = early_reset_static_par0_go_out;
wire _guard782 = _guard780 & _guard781;
wire _guard783 = early_reset_static_par0_go_out;
wire _guard784 = ~_guard0;
wire _guard785 = early_reset_static_par0_go_out;
wire _guard786 = _guard784 & _guard785;
wire _guard787 = early_reset_static_par0_go_out;
wire _guard788 = ~_guard0;
wire _guard789 = early_reset_static_par0_go_out;
wire _guard790 = _guard788 & _guard789;
wire _guard791 = early_reset_static_par0_go_out;
wire _guard792 = ~_guard0;
wire _guard793 = early_reset_static_par0_go_out;
wire _guard794 = _guard792 & _guard793;
wire _guard795 = cond_wire_out;
wire _guard796 = early_reset_static_par0_go_out;
wire _guard797 = _guard795 & _guard796;
wire _guard798 = cond_wire_out;
wire _guard799 = early_reset_static_par0_go_out;
wire _guard800 = _guard798 & _guard799;
wire _guard801 = cond_wire17_out;
wire _guard802 = early_reset_static_par0_go_out;
wire _guard803 = _guard801 & _guard802;
wire _guard804 = cond_wire15_out;
wire _guard805 = early_reset_static_par0_go_out;
wire _guard806 = _guard804 & _guard805;
wire _guard807 = fsm_out == 1'd0;
wire _guard808 = cond_wire15_out;
wire _guard809 = _guard807 & _guard808;
wire _guard810 = fsm_out == 1'd0;
wire _guard811 = _guard809 & _guard810;
wire _guard812 = fsm_out == 1'd0;
wire _guard813 = cond_wire17_out;
wire _guard814 = _guard812 & _guard813;
wire _guard815 = fsm_out == 1'd0;
wire _guard816 = _guard814 & _guard815;
wire _guard817 = _guard811 | _guard816;
wire _guard818 = early_reset_static_par0_go_out;
wire _guard819 = _guard817 & _guard818;
wire _guard820 = fsm_out == 1'd0;
wire _guard821 = cond_wire15_out;
wire _guard822 = _guard820 & _guard821;
wire _guard823 = fsm_out == 1'd0;
wire _guard824 = _guard822 & _guard823;
wire _guard825 = fsm_out == 1'd0;
wire _guard826 = cond_wire17_out;
wire _guard827 = _guard825 & _guard826;
wire _guard828 = fsm_out == 1'd0;
wire _guard829 = _guard827 & _guard828;
wire _guard830 = _guard824 | _guard829;
wire _guard831 = early_reset_static_par0_go_out;
wire _guard832 = _guard830 & _guard831;
wire _guard833 = fsm_out == 1'd0;
wire _guard834 = cond_wire15_out;
wire _guard835 = _guard833 & _guard834;
wire _guard836 = fsm_out == 1'd0;
wire _guard837 = _guard835 & _guard836;
wire _guard838 = fsm_out == 1'd0;
wire _guard839 = cond_wire17_out;
wire _guard840 = _guard838 & _guard839;
wire _guard841 = fsm_out == 1'd0;
wire _guard842 = _guard840 & _guard841;
wire _guard843 = _guard837 | _guard842;
wire _guard844 = early_reset_static_par0_go_out;
wire _guard845 = _guard843 & _guard844;
wire _guard846 = cond_wire16_out;
wire _guard847 = early_reset_static_par0_go_out;
wire _guard848 = _guard846 & _guard847;
wire _guard849 = cond_wire16_out;
wire _guard850 = early_reset_static_par0_go_out;
wire _guard851 = _guard849 & _guard850;
wire _guard852 = cond_wire46_out;
wire _guard853 = early_reset_static_par0_go_out;
wire _guard854 = _guard852 & _guard853;
wire _guard855 = cond_wire46_out;
wire _guard856 = early_reset_static_par0_go_out;
wire _guard857 = _guard855 & _guard856;
wire _guard858 = cond_wire56_out;
wire _guard859 = early_reset_static_par0_go_out;
wire _guard860 = _guard858 & _guard859;
wire _guard861 = cond_wire54_out;
wire _guard862 = early_reset_static_par0_go_out;
wire _guard863 = _guard861 & _guard862;
wire _guard864 = fsm_out == 1'd0;
wire _guard865 = cond_wire54_out;
wire _guard866 = _guard864 & _guard865;
wire _guard867 = fsm_out == 1'd0;
wire _guard868 = _guard866 & _guard867;
wire _guard869 = fsm_out == 1'd0;
wire _guard870 = cond_wire56_out;
wire _guard871 = _guard869 & _guard870;
wire _guard872 = fsm_out == 1'd0;
wire _guard873 = _guard871 & _guard872;
wire _guard874 = _guard868 | _guard873;
wire _guard875 = early_reset_static_par0_go_out;
wire _guard876 = _guard874 & _guard875;
wire _guard877 = fsm_out == 1'd0;
wire _guard878 = cond_wire54_out;
wire _guard879 = _guard877 & _guard878;
wire _guard880 = fsm_out == 1'd0;
wire _guard881 = _guard879 & _guard880;
wire _guard882 = fsm_out == 1'd0;
wire _guard883 = cond_wire56_out;
wire _guard884 = _guard882 & _guard883;
wire _guard885 = fsm_out == 1'd0;
wire _guard886 = _guard884 & _guard885;
wire _guard887 = _guard881 | _guard886;
wire _guard888 = early_reset_static_par0_go_out;
wire _guard889 = _guard887 & _guard888;
wire _guard890 = fsm_out == 1'd0;
wire _guard891 = cond_wire54_out;
wire _guard892 = _guard890 & _guard891;
wire _guard893 = fsm_out == 1'd0;
wire _guard894 = _guard892 & _guard893;
wire _guard895 = fsm_out == 1'd0;
wire _guard896 = cond_wire56_out;
wire _guard897 = _guard895 & _guard896;
wire _guard898 = fsm_out == 1'd0;
wire _guard899 = _guard897 & _guard898;
wire _guard900 = _guard894 | _guard899;
wire _guard901 = early_reset_static_par0_go_out;
wire _guard902 = _guard900 & _guard901;
wire _guard903 = cond_wire46_out;
wire _guard904 = early_reset_static_par0_go_out;
wire _guard905 = _guard903 & _guard904;
wire _guard906 = cond_wire46_out;
wire _guard907 = early_reset_static_par0_go_out;
wire _guard908 = _guard906 & _guard907;
wire _guard909 = early_reset_static_par0_go_out;
wire _guard910 = early_reset_static_par0_go_out;
wire _guard911 = early_reset_static_par0_go_out;
wire _guard912 = early_reset_static_par0_go_out;
wire _guard913 = early_reset_static_par0_go_out;
wire _guard914 = early_reset_static_par0_go_out;
wire _guard915 = ~_guard0;
wire _guard916 = early_reset_static_par0_go_out;
wire _guard917 = _guard915 & _guard916;
wire _guard918 = early_reset_static_par0_go_out;
wire _guard919 = early_reset_static_par0_go_out;
wire _guard920 = early_reset_static_par0_go_out;
wire _guard921 = early_reset_static_par0_go_out;
wire _guard922 = ~_guard0;
wire _guard923 = early_reset_static_par0_go_out;
wire _guard924 = _guard922 & _guard923;
wire _guard925 = early_reset_static_par0_go_out;
wire _guard926 = early_reset_static_par0_go_out;
wire _guard927 = early_reset_static_par0_go_out;
wire _guard928 = early_reset_static_par0_go_out;
wire _guard929 = early_reset_static_par0_go_out;
wire _guard930 = early_reset_static_par0_go_out;
wire _guard931 = early_reset_static_par0_go_out;
wire _guard932 = ~_guard0;
wire _guard933 = early_reset_static_par0_go_out;
wire _guard934 = _guard932 & _guard933;
wire _guard935 = early_reset_static_par0_go_out;
wire _guard936 = ~_guard0;
wire _guard937 = early_reset_static_par0_go_out;
wire _guard938 = _guard936 & _guard937;
wire _guard939 = cond_wire12_out;
wire _guard940 = early_reset_static_par0_go_out;
wire _guard941 = _guard939 & _guard940;
wire _guard942 = cond_wire10_out;
wire _guard943 = early_reset_static_par0_go_out;
wire _guard944 = _guard942 & _guard943;
wire _guard945 = fsm_out == 1'd0;
wire _guard946 = cond_wire10_out;
wire _guard947 = _guard945 & _guard946;
wire _guard948 = fsm_out == 1'd0;
wire _guard949 = _guard947 & _guard948;
wire _guard950 = fsm_out == 1'd0;
wire _guard951 = cond_wire12_out;
wire _guard952 = _guard950 & _guard951;
wire _guard953 = fsm_out == 1'd0;
wire _guard954 = _guard952 & _guard953;
wire _guard955 = _guard949 | _guard954;
wire _guard956 = early_reset_static_par0_go_out;
wire _guard957 = _guard955 & _guard956;
wire _guard958 = fsm_out == 1'd0;
wire _guard959 = cond_wire10_out;
wire _guard960 = _guard958 & _guard959;
wire _guard961 = fsm_out == 1'd0;
wire _guard962 = _guard960 & _guard961;
wire _guard963 = fsm_out == 1'd0;
wire _guard964 = cond_wire12_out;
wire _guard965 = _guard963 & _guard964;
wire _guard966 = fsm_out == 1'd0;
wire _guard967 = _guard965 & _guard966;
wire _guard968 = _guard962 | _guard967;
wire _guard969 = early_reset_static_par0_go_out;
wire _guard970 = _guard968 & _guard969;
wire _guard971 = fsm_out == 1'd0;
wire _guard972 = cond_wire10_out;
wire _guard973 = _guard971 & _guard972;
wire _guard974 = fsm_out == 1'd0;
wire _guard975 = _guard973 & _guard974;
wire _guard976 = fsm_out == 1'd0;
wire _guard977 = cond_wire12_out;
wire _guard978 = _guard976 & _guard977;
wire _guard979 = fsm_out == 1'd0;
wire _guard980 = _guard978 & _guard979;
wire _guard981 = _guard975 | _guard980;
wire _guard982 = early_reset_static_par0_go_out;
wire _guard983 = _guard981 & _guard982;
wire _guard984 = fsm0_out == 5'd0;
wire _guard985 = early_reset_static_seq_go_out;
wire _guard986 = _guard984 & _guard985;
wire _guard987 = cond_wire_out;
wire _guard988 = early_reset_static_par0_go_out;
wire _guard989 = _guard987 & _guard988;
wire _guard990 = _guard986 | _guard989;
wire _guard991 = cond_wire_out;
wire _guard992 = early_reset_static_par0_go_out;
wire _guard993 = _guard991 & _guard992;
wire _guard994 = fsm0_out == 5'd0;
wire _guard995 = early_reset_static_seq_go_out;
wire _guard996 = _guard994 & _guard995;
wire _guard997 = fsm0_out == 5'd0;
wire _guard998 = early_reset_static_seq_go_out;
wire _guard999 = _guard997 & _guard998;
wire _guard1000 = cond_wire19_out;
wire _guard1001 = early_reset_static_par0_go_out;
wire _guard1002 = _guard1000 & _guard1001;
wire _guard1003 = _guard999 | _guard1002;
wire _guard1004 = cond_wire19_out;
wire _guard1005 = early_reset_static_par0_go_out;
wire _guard1006 = _guard1004 & _guard1005;
wire _guard1007 = fsm0_out == 5'd0;
wire _guard1008 = early_reset_static_seq_go_out;
wire _guard1009 = _guard1007 & _guard1008;
wire _guard1010 = early_reset_static_par0_go_out;
wire _guard1011 = early_reset_static_par0_go_out;
wire _guard1012 = fsm0_out == 5'd0;
wire _guard1013 = early_reset_static_seq_go_out;
wire _guard1014 = _guard1012 & _guard1013;
wire _guard1015 = early_reset_static_par0_go_out;
wire _guard1016 = _guard1014 | _guard1015;
wire _guard1017 = fsm0_out == 5'd0;
wire _guard1018 = early_reset_static_seq_go_out;
wire _guard1019 = _guard1017 & _guard1018;
wire _guard1020 = early_reset_static_par0_go_out;
wire _guard1021 = early_reset_static_par0_go_out;
wire _guard1022 = early_reset_static_par0_go_out;
wire _guard1023 = early_reset_static_par0_go_out;
wire _guard1024 = early_reset_static_par0_go_out;
wire _guard1025 = early_reset_static_par0_go_out;
wire _guard1026 = early_reset_static_par0_go_out;
wire _guard1027 = early_reset_static_par0_go_out;
wire _guard1028 = early_reset_static_par0_go_out;
wire _guard1029 = early_reset_static_par0_go_out;
wire _guard1030 = early_reset_static_par0_go_out;
wire _guard1031 = early_reset_static_par0_go_out;
wire _guard1032 = early_reset_static_par0_go_out;
wire _guard1033 = early_reset_static_par0_go_out;
wire _guard1034 = early_reset_static_par0_go_out;
wire _guard1035 = early_reset_static_par0_go_out;
wire _guard1036 = early_reset_static_par0_go_out;
wire _guard1037 = early_reset_static_par0_go_out;
wire _guard1038 = early_reset_static_par0_go_out;
wire _guard1039 = early_reset_static_par0_go_out;
wire _guard1040 = early_reset_static_par0_go_out;
wire _guard1041 = cond_wire43_out;
wire _guard1042 = early_reset_static_par0_go_out;
wire _guard1043 = _guard1041 & _guard1042;
wire _guard1044 = cond_wire41_out;
wire _guard1045 = early_reset_static_par0_go_out;
wire _guard1046 = _guard1044 & _guard1045;
wire _guard1047 = fsm_out == 1'd0;
wire _guard1048 = cond_wire41_out;
wire _guard1049 = _guard1047 & _guard1048;
wire _guard1050 = fsm_out == 1'd0;
wire _guard1051 = _guard1049 & _guard1050;
wire _guard1052 = fsm_out == 1'd0;
wire _guard1053 = cond_wire43_out;
wire _guard1054 = _guard1052 & _guard1053;
wire _guard1055 = fsm_out == 1'd0;
wire _guard1056 = _guard1054 & _guard1055;
wire _guard1057 = _guard1051 | _guard1056;
wire _guard1058 = early_reset_static_par0_go_out;
wire _guard1059 = _guard1057 & _guard1058;
wire _guard1060 = fsm_out == 1'd0;
wire _guard1061 = cond_wire41_out;
wire _guard1062 = _guard1060 & _guard1061;
wire _guard1063 = fsm_out == 1'd0;
wire _guard1064 = _guard1062 & _guard1063;
wire _guard1065 = fsm_out == 1'd0;
wire _guard1066 = cond_wire43_out;
wire _guard1067 = _guard1065 & _guard1066;
wire _guard1068 = fsm_out == 1'd0;
wire _guard1069 = _guard1067 & _guard1068;
wire _guard1070 = _guard1064 | _guard1069;
wire _guard1071 = early_reset_static_par0_go_out;
wire _guard1072 = _guard1070 & _guard1071;
wire _guard1073 = fsm_out == 1'd0;
wire _guard1074 = cond_wire41_out;
wire _guard1075 = _guard1073 & _guard1074;
wire _guard1076 = fsm_out == 1'd0;
wire _guard1077 = _guard1075 & _guard1076;
wire _guard1078 = fsm_out == 1'd0;
wire _guard1079 = cond_wire43_out;
wire _guard1080 = _guard1078 & _guard1079;
wire _guard1081 = fsm_out == 1'd0;
wire _guard1082 = _guard1080 & _guard1081;
wire _guard1083 = _guard1077 | _guard1082;
wire _guard1084 = early_reset_static_par0_go_out;
wire _guard1085 = _guard1083 & _guard1084;
wire _guard1086 = cond_wire51_out;
wire _guard1087 = early_reset_static_par0_go_out;
wire _guard1088 = _guard1086 & _guard1087;
wire _guard1089 = cond_wire49_out;
wire _guard1090 = early_reset_static_par0_go_out;
wire _guard1091 = _guard1089 & _guard1090;
wire _guard1092 = fsm_out == 1'd0;
wire _guard1093 = cond_wire49_out;
wire _guard1094 = _guard1092 & _guard1093;
wire _guard1095 = fsm_out == 1'd0;
wire _guard1096 = _guard1094 & _guard1095;
wire _guard1097 = fsm_out == 1'd0;
wire _guard1098 = cond_wire51_out;
wire _guard1099 = _guard1097 & _guard1098;
wire _guard1100 = fsm_out == 1'd0;
wire _guard1101 = _guard1099 & _guard1100;
wire _guard1102 = _guard1096 | _guard1101;
wire _guard1103 = early_reset_static_par0_go_out;
wire _guard1104 = _guard1102 & _guard1103;
wire _guard1105 = fsm_out == 1'd0;
wire _guard1106 = cond_wire49_out;
wire _guard1107 = _guard1105 & _guard1106;
wire _guard1108 = fsm_out == 1'd0;
wire _guard1109 = _guard1107 & _guard1108;
wire _guard1110 = fsm_out == 1'd0;
wire _guard1111 = cond_wire51_out;
wire _guard1112 = _guard1110 & _guard1111;
wire _guard1113 = fsm_out == 1'd0;
wire _guard1114 = _guard1112 & _guard1113;
wire _guard1115 = _guard1109 | _guard1114;
wire _guard1116 = early_reset_static_par0_go_out;
wire _guard1117 = _guard1115 & _guard1116;
wire _guard1118 = fsm_out == 1'd0;
wire _guard1119 = cond_wire49_out;
wire _guard1120 = _guard1118 & _guard1119;
wire _guard1121 = fsm_out == 1'd0;
wire _guard1122 = _guard1120 & _guard1121;
wire _guard1123 = fsm_out == 1'd0;
wire _guard1124 = cond_wire51_out;
wire _guard1125 = _guard1123 & _guard1124;
wire _guard1126 = fsm_out == 1'd0;
wire _guard1127 = _guard1125 & _guard1126;
wire _guard1128 = _guard1122 | _guard1127;
wire _guard1129 = early_reset_static_par0_go_out;
wire _guard1130 = _guard1128 & _guard1129;
wire _guard1131 = cond_wire60_out;
wire _guard1132 = early_reset_static_par0_go_out;
wire _guard1133 = _guard1131 & _guard1132;
wire _guard1134 = cond_wire58_out;
wire _guard1135 = early_reset_static_par0_go_out;
wire _guard1136 = _guard1134 & _guard1135;
wire _guard1137 = fsm_out == 1'd0;
wire _guard1138 = cond_wire58_out;
wire _guard1139 = _guard1137 & _guard1138;
wire _guard1140 = fsm_out == 1'd0;
wire _guard1141 = _guard1139 & _guard1140;
wire _guard1142 = fsm_out == 1'd0;
wire _guard1143 = cond_wire60_out;
wire _guard1144 = _guard1142 & _guard1143;
wire _guard1145 = fsm_out == 1'd0;
wire _guard1146 = _guard1144 & _guard1145;
wire _guard1147 = _guard1141 | _guard1146;
wire _guard1148 = early_reset_static_par0_go_out;
wire _guard1149 = _guard1147 & _guard1148;
wire _guard1150 = fsm_out == 1'd0;
wire _guard1151 = cond_wire58_out;
wire _guard1152 = _guard1150 & _guard1151;
wire _guard1153 = fsm_out == 1'd0;
wire _guard1154 = _guard1152 & _guard1153;
wire _guard1155 = fsm_out == 1'd0;
wire _guard1156 = cond_wire60_out;
wire _guard1157 = _guard1155 & _guard1156;
wire _guard1158 = fsm_out == 1'd0;
wire _guard1159 = _guard1157 & _guard1158;
wire _guard1160 = _guard1154 | _guard1159;
wire _guard1161 = early_reset_static_par0_go_out;
wire _guard1162 = _guard1160 & _guard1161;
wire _guard1163 = fsm_out == 1'd0;
wire _guard1164 = cond_wire58_out;
wire _guard1165 = _guard1163 & _guard1164;
wire _guard1166 = fsm_out == 1'd0;
wire _guard1167 = _guard1165 & _guard1166;
wire _guard1168 = fsm_out == 1'd0;
wire _guard1169 = cond_wire60_out;
wire _guard1170 = _guard1168 & _guard1169;
wire _guard1171 = fsm_out == 1'd0;
wire _guard1172 = _guard1170 & _guard1171;
wire _guard1173 = _guard1167 | _guard1172;
wire _guard1174 = early_reset_static_par0_go_out;
wire _guard1175 = _guard1173 & _guard1174;
wire _guard1176 = early_reset_static_par0_go_out;
wire _guard1177 = early_reset_static_par0_go_out;
wire _guard1178 = early_reset_static_par0_go_out;
wire _guard1179 = ~_guard0;
wire _guard1180 = early_reset_static_par0_go_out;
wire _guard1181 = _guard1179 & _guard1180;
wire _guard1182 = early_reset_static_par0_go_out;
wire _guard1183 = early_reset_static_par0_go_out;
wire _guard1184 = early_reset_static_par0_go_out;
wire _guard1185 = early_reset_static_par0_go_out;
wire _guard1186 = early_reset_static_par0_go_out;
wire _guard1187 = ~_guard0;
wire _guard1188 = early_reset_static_par0_go_out;
wire _guard1189 = _guard1187 & _guard1188;
wire _guard1190 = early_reset_static_par0_go_out;
wire _guard1191 = early_reset_static_par0_go_out;
wire _guard1192 = early_reset_static_par0_go_out;
wire _guard1193 = early_reset_static_par0_go_out;
wire _guard1194 = early_reset_static_par0_go_out;
wire _guard1195 = early_reset_static_par0_go_out;
wire _guard1196 = early_reset_static_seq_go_out;
wire _guard1197 = fsm0_out != 5'd16;
wire _guard1198 = early_reset_static_seq_go_out;
wire _guard1199 = _guard1197 & _guard1198;
wire _guard1200 = fsm0_out == 5'd16;
wire _guard1201 = early_reset_static_seq_go_out;
wire _guard1202 = _guard1200 & _guard1201;
wire _guard1203 = cond_wire21_out;
wire _guard1204 = early_reset_static_par0_go_out;
wire _guard1205 = _guard1203 & _guard1204;
wire _guard1206 = cond_wire21_out;
wire _guard1207 = early_reset_static_par0_go_out;
wire _guard1208 = _guard1206 & _guard1207;
wire _guard1209 = cond_wire38_out;
wire _guard1210 = early_reset_static_par0_go_out;
wire _guard1211 = _guard1209 & _guard1210;
wire _guard1212 = cond_wire38_out;
wire _guard1213 = early_reset_static_par0_go_out;
wire _guard1214 = _guard1212 & _guard1213;
wire _guard1215 = cond_wire42_out;
wire _guard1216 = early_reset_static_par0_go_out;
wire _guard1217 = _guard1215 & _guard1216;
wire _guard1218 = cond_wire42_out;
wire _guard1219 = early_reset_static_par0_go_out;
wire _guard1220 = _guard1218 & _guard1219;
wire _guard1221 = fsm0_out == 5'd0;
wire _guard1222 = early_reset_static_seq_go_out;
wire _guard1223 = _guard1221 & _guard1222;
wire _guard1224 = early_reset_static_par0_go_out;
wire _guard1225 = _guard1223 | _guard1224;
wire _guard1226 = fsm0_out == 5'd0;
wire _guard1227 = early_reset_static_seq_go_out;
wire _guard1228 = _guard1226 & _guard1227;
wire _guard1229 = early_reset_static_par0_go_out;
wire _guard1230 = fsm0_out == 5'd0;
wire _guard1231 = early_reset_static_seq_go_out;
wire _guard1232 = _guard1230 & _guard1231;
wire _guard1233 = early_reset_static_par0_go_out;
wire _guard1234 = _guard1232 | _guard1233;
wire _guard1235 = fsm0_out == 5'd0;
wire _guard1236 = early_reset_static_seq_go_out;
wire _guard1237 = _guard1235 & _guard1236;
wire _guard1238 = early_reset_static_par0_go_out;
wire _guard1239 = fsm0_out == 5'd0;
wire _guard1240 = early_reset_static_seq_go_out;
wire _guard1241 = _guard1239 & _guard1240;
wire _guard1242 = early_reset_static_par0_go_out;
wire _guard1243 = _guard1241 | _guard1242;
wire _guard1244 = early_reset_static_par0_go_out;
wire _guard1245 = fsm0_out == 5'd0;
wire _guard1246 = early_reset_static_seq_go_out;
wire _guard1247 = _guard1245 & _guard1246;
wire _guard1248 = early_reset_static_par0_go_out;
wire _guard1249 = early_reset_static_par0_go_out;
wire _guard1250 = early_reset_static_par0_go_out;
wire _guard1251 = early_reset_static_par0_go_out;
wire _guard1252 = early_reset_static_par0_go_out;
wire _guard1253 = ~_guard0;
wire _guard1254 = early_reset_static_par0_go_out;
wire _guard1255 = _guard1253 & _guard1254;
wire _guard1256 = early_reset_static_par0_go_out;
wire _guard1257 = early_reset_static_par0_go_out;
wire _guard1258 = early_reset_static_par0_go_out;
wire _guard1259 = early_reset_static_par0_go_out;
wire _guard1260 = ~_guard0;
wire _guard1261 = early_reset_static_par0_go_out;
wire _guard1262 = _guard1260 & _guard1261;
wire _guard1263 = early_reset_static_par0_go_out;
wire _guard1264 = early_reset_static_par0_go_out;
wire _guard1265 = early_reset_static_par0_go_out;
wire _guard1266 = early_reset_static_par0_go_out;
wire _guard1267 = early_reset_static_par0_go_out;
wire _guard1268 = early_reset_static_par0_go_out;
wire _guard1269 = ~_guard0;
wire _guard1270 = early_reset_static_par0_go_out;
wire _guard1271 = _guard1269 & _guard1270;
wire _guard1272 = early_reset_static_par0_go_out;
wire _guard1273 = early_reset_static_par0_go_out;
wire _guard1274 = ~_guard0;
wire _guard1275 = early_reset_static_par0_go_out;
wire _guard1276 = _guard1274 & _guard1275;
wire _guard1277 = early_reset_static_par0_go_out;
wire _guard1278 = ~_guard0;
wire _guard1279 = early_reset_static_par0_go_out;
wire _guard1280 = _guard1278 & _guard1279;
wire _guard1281 = early_reset_static_par0_go_out;
wire _guard1282 = fsm0_out == 5'd0;
wire _guard1283 = signal_reg_out;
wire _guard1284 = _guard1282 & _guard1283;
wire _guard1285 = cond_wire4_out;
wire _guard1286 = early_reset_static_par0_go_out;
wire _guard1287 = _guard1285 & _guard1286;
wire _guard1288 = cond_wire4_out;
wire _guard1289 = early_reset_static_par0_go_out;
wire _guard1290 = _guard1288 & _guard1289;
wire _guard1291 = cond_wire6_out;
wire _guard1292 = early_reset_static_par0_go_out;
wire _guard1293 = _guard1291 & _guard1292;
wire _guard1294 = cond_wire6_out;
wire _guard1295 = early_reset_static_par0_go_out;
wire _guard1296 = _guard1294 & _guard1295;
wire _guard1297 = cond_wire33_out;
wire _guard1298 = early_reset_static_par0_go_out;
wire _guard1299 = _guard1297 & _guard1298;
wire _guard1300 = cond_wire33_out;
wire _guard1301 = early_reset_static_par0_go_out;
wire _guard1302 = _guard1300 & _guard1301;
wire _guard1303 = cond_wire53_out;
wire _guard1304 = early_reset_static_par0_go_out;
wire _guard1305 = _guard1303 & _guard1304;
wire _guard1306 = cond_wire53_out;
wire _guard1307 = early_reset_static_par0_go_out;
wire _guard1308 = _guard1306 & _guard1307;
wire _guard1309 = early_reset_static_par0_go_out;
wire _guard1310 = early_reset_static_par0_go_out;
wire _guard1311 = early_reset_static_par0_go_out;
wire _guard1312 = early_reset_static_par0_go_out;
wire _guard1313 = early_reset_static_par0_go_out;
wire _guard1314 = early_reset_static_par0_go_out;
wire _guard1315 = early_reset_static_par0_go_out;
wire _guard1316 = early_reset_static_par0_go_out;
wire _guard1317 = early_reset_static_par0_go_out;
wire _guard1318 = early_reset_static_par0_go_out;
wire _guard1319 = fsm0_out == 5'd0;
wire _guard1320 = early_reset_static_seq_go_out;
wire _guard1321 = _guard1319 & _guard1320;
wire _guard1322 = early_reset_static_par0_go_out;
wire _guard1323 = _guard1321 | _guard1322;
wire _guard1324 = early_reset_static_par0_go_out;
wire _guard1325 = fsm0_out == 5'd0;
wire _guard1326 = early_reset_static_seq_go_out;
wire _guard1327 = _guard1325 & _guard1326;
wire _guard1328 = fsm0_out == 5'd0;
wire _guard1329 = early_reset_static_seq_go_out;
wire _guard1330 = _guard1328 & _guard1329;
wire _guard1331 = early_reset_static_par0_go_out;
wire _guard1332 = _guard1330 | _guard1331;
wire _guard1333 = early_reset_static_par0_go_out;
wire _guard1334 = fsm0_out == 5'd0;
wire _guard1335 = early_reset_static_seq_go_out;
wire _guard1336 = _guard1334 & _guard1335;
wire _guard1337 = fsm0_out == 5'd0;
wire _guard1338 = early_reset_static_seq_go_out;
wire _guard1339 = _guard1337 & _guard1338;
wire _guard1340 = early_reset_static_par0_go_out;
wire _guard1341 = _guard1339 | _guard1340;
wire _guard1342 = fsm0_out == 5'd0;
wire _guard1343 = early_reset_static_seq_go_out;
wire _guard1344 = _guard1342 & _guard1343;
wire _guard1345 = early_reset_static_par0_go_out;
wire _guard1346 = early_reset_static_par0_go_out;
wire _guard1347 = early_reset_static_par0_go_out;
wire _guard1348 = early_reset_static_par0_go_out;
wire _guard1349 = early_reset_static_par0_go_out;
wire _guard1350 = early_reset_static_par0_go_out;
wire _guard1351 = early_reset_static_par0_go_out;
wire _guard1352 = early_reset_static_par0_go_out;
wire _guard1353 = early_reset_static_par0_go_out;
wire _guard1354 = ~_guard0;
wire _guard1355 = early_reset_static_par0_go_out;
wire _guard1356 = _guard1354 & _guard1355;
wire _guard1357 = early_reset_static_par0_go_out;
wire _guard1358 = early_reset_static_par0_go_out;
wire _guard1359 = early_reset_static_par0_go_out;
wire _guard1360 = ~_guard0;
wire _guard1361 = early_reset_static_par0_go_out;
wire _guard1362 = _guard1360 & _guard1361;
wire _guard1363 = early_reset_static_par0_go_out;
wire _guard1364 = early_reset_static_par0_go_out;
wire _guard1365 = early_reset_static_par0_go_out;
wire _guard1366 = early_reset_static_par0_go_out;
wire _guard1367 = ~_guard0;
wire _guard1368 = early_reset_static_par0_go_out;
wire _guard1369 = _guard1367 & _guard1368;
wire _guard1370 = early_reset_static_par0_go_out;
wire _guard1371 = early_reset_static_par0_go_out;
wire _guard1372 = early_reset_static_par0_go_out;
wire _guard1373 = ~_guard0;
wire _guard1374 = early_reset_static_par0_go_out;
wire _guard1375 = _guard1373 & _guard1374;
wire _guard1376 = early_reset_static_par0_go_out;
wire _guard1377 = early_reset_static_par0_go_out;
wire _guard1378 = wrapper_early_reset_static_seq_go_out;
wire _guard1379 = cond_wire9_out;
wire _guard1380 = early_reset_static_par0_go_out;
wire _guard1381 = _guard1379 & _guard1380;
wire _guard1382 = cond_wire9_out;
wire _guard1383 = early_reset_static_par0_go_out;
wire _guard1384 = _guard1382 & _guard1383;
wire _guard1385 = cond_wire6_out;
wire _guard1386 = early_reset_static_par0_go_out;
wire _guard1387 = _guard1385 & _guard1386;
wire _guard1388 = cond_wire6_out;
wire _guard1389 = early_reset_static_par0_go_out;
wire _guard1390 = _guard1388 & _guard1389;
wire _guard1391 = cond_wire59_out;
wire _guard1392 = early_reset_static_par0_go_out;
wire _guard1393 = _guard1391 & _guard1392;
wire _guard1394 = cond_wire59_out;
wire _guard1395 = early_reset_static_par0_go_out;
wire _guard1396 = _guard1394 & _guard1395;
wire _guard1397 = cond_wire_out;
wire _guard1398 = early_reset_static_par0_go_out;
wire _guard1399 = _guard1397 & _guard1398;
wire _guard1400 = cond_wire_out;
wire _guard1401 = early_reset_static_par0_go_out;
wire _guard1402 = _guard1400 & _guard1401;
wire _guard1403 = cond_wire_out;
wire _guard1404 = early_reset_static_par0_go_out;
wire _guard1405 = _guard1403 & _guard1404;
wire _guard1406 = cond_wire_out;
wire _guard1407 = early_reset_static_par0_go_out;
wire _guard1408 = _guard1406 & _guard1407;
wire _guard1409 = early_reset_static_par0_go_out;
wire _guard1410 = early_reset_static_par0_go_out;
wire _guard1411 = early_reset_static_par0_go_out;
wire _guard1412 = early_reset_static_par0_go_out;
wire _guard1413 = fsm0_out == 5'd0;
wire _guard1414 = early_reset_static_seq_go_out;
wire _guard1415 = _guard1413 & _guard1414;
wire _guard1416 = early_reset_static_par0_go_out;
wire _guard1417 = _guard1415 | _guard1416;
wire _guard1418 = early_reset_static_par0_go_out;
wire _guard1419 = fsm0_out == 5'd0;
wire _guard1420 = early_reset_static_seq_go_out;
wire _guard1421 = _guard1419 & _guard1420;
wire _guard1422 = early_reset_static_par0_go_out;
wire _guard1423 = early_reset_static_par0_go_out;
wire _guard1424 = early_reset_static_par0_go_out;
wire _guard1425 = early_reset_static_par0_go_out;
wire _guard1426 = early_reset_static_par0_go_out;
wire _guard1427 = ~_guard0;
wire _guard1428 = early_reset_static_par0_go_out;
wire _guard1429 = _guard1427 & _guard1428;
wire _guard1430 = ~_guard0;
wire _guard1431 = early_reset_static_par0_go_out;
wire _guard1432 = _guard1430 & _guard1431;
wire _guard1433 = early_reset_static_par0_go_out;
wire _guard1434 = early_reset_static_par0_go_out;
wire _guard1435 = early_reset_static_par0_go_out;
wire _guard1436 = early_reset_static_par0_go_out;
wire _guard1437 = ~_guard0;
wire _guard1438 = early_reset_static_par0_go_out;
wire _guard1439 = _guard1437 & _guard1438;
wire _guard1440 = early_reset_static_par0_go_out;
wire _guard1441 = early_reset_static_par0_go_out;
wire _guard1442 = early_reset_static_par0_go_out;
wire _guard1443 = early_reset_static_par0_go_out;
wire _guard1444 = early_reset_static_par0_go_out;
wire _guard1445 = early_reset_static_par0_go_out;
wire _guard1446 = early_reset_static_par0_go_out;
wire _guard1447 = early_reset_static_par0_go_out;
wire _guard1448 = early_reset_static_par0_go_out;
wire _guard1449 = ~_guard0;
wire _guard1450 = early_reset_static_par0_go_out;
wire _guard1451 = _guard1449 & _guard1450;
wire _guard1452 = ~_guard0;
wire _guard1453 = early_reset_static_par0_go_out;
wire _guard1454 = _guard1452 & _guard1453;
wire _guard1455 = early_reset_static_par0_go_out;
wire _guard1456 = early_reset_static_par0_go_out;
wire _guard1457 = early_reset_static_par0_go_out;
wire _guard1458 = ~_guard0;
wire _guard1459 = early_reset_static_par0_go_out;
wire _guard1460 = _guard1458 & _guard1459;
wire _guard1461 = early_reset_static_par0_go_out;
wire _guard1462 = ~_guard0;
wire _guard1463 = early_reset_static_par0_go_out;
wire _guard1464 = _guard1462 & _guard1463;
wire _guard1465 = early_reset_static_par0_go_out;
wire _guard1466 = early_reset_static_par0_go_out;
wire _guard1467 = early_reset_static_par0_go_out;
wire _guard1468 = fsm0_out == 5'd0;
wire _guard1469 = signal_reg_out;
wire _guard1470 = _guard1468 & _guard1469;
wire _guard1471 = fsm0_out == 5'd0;
wire _guard1472 = signal_reg_out;
wire _guard1473 = ~_guard1472;
wire _guard1474 = _guard1471 & _guard1473;
wire _guard1475 = wrapper_early_reset_static_seq_go_out;
wire _guard1476 = _guard1474 & _guard1475;
wire _guard1477 = _guard1470 | _guard1476;
wire _guard1478 = fsm0_out == 5'd0;
wire _guard1479 = signal_reg_out;
wire _guard1480 = ~_guard1479;
wire _guard1481 = _guard1478 & _guard1480;
wire _guard1482 = wrapper_early_reset_static_seq_go_out;
wire _guard1483 = _guard1481 & _guard1482;
wire _guard1484 = fsm0_out == 5'd0;
wire _guard1485 = signal_reg_out;
wire _guard1486 = _guard1484 & _guard1485;
wire _guard1487 = cond_wire39_out;
wire _guard1488 = early_reset_static_par0_go_out;
wire _guard1489 = _guard1487 & _guard1488;
wire _guard1490 = cond_wire37_out;
wire _guard1491 = early_reset_static_par0_go_out;
wire _guard1492 = _guard1490 & _guard1491;
wire _guard1493 = fsm_out == 1'd0;
wire _guard1494 = cond_wire37_out;
wire _guard1495 = _guard1493 & _guard1494;
wire _guard1496 = fsm_out == 1'd0;
wire _guard1497 = _guard1495 & _guard1496;
wire _guard1498 = fsm_out == 1'd0;
wire _guard1499 = cond_wire39_out;
wire _guard1500 = _guard1498 & _guard1499;
wire _guard1501 = fsm_out == 1'd0;
wire _guard1502 = _guard1500 & _guard1501;
wire _guard1503 = _guard1497 | _guard1502;
wire _guard1504 = early_reset_static_par0_go_out;
wire _guard1505 = _guard1503 & _guard1504;
wire _guard1506 = fsm_out == 1'd0;
wire _guard1507 = cond_wire37_out;
wire _guard1508 = _guard1506 & _guard1507;
wire _guard1509 = fsm_out == 1'd0;
wire _guard1510 = _guard1508 & _guard1509;
wire _guard1511 = fsm_out == 1'd0;
wire _guard1512 = cond_wire39_out;
wire _guard1513 = _guard1511 & _guard1512;
wire _guard1514 = fsm_out == 1'd0;
wire _guard1515 = _guard1513 & _guard1514;
wire _guard1516 = _guard1510 | _guard1515;
wire _guard1517 = early_reset_static_par0_go_out;
wire _guard1518 = _guard1516 & _guard1517;
wire _guard1519 = fsm_out == 1'd0;
wire _guard1520 = cond_wire37_out;
wire _guard1521 = _guard1519 & _guard1520;
wire _guard1522 = fsm_out == 1'd0;
wire _guard1523 = _guard1521 & _guard1522;
wire _guard1524 = fsm_out == 1'd0;
wire _guard1525 = cond_wire39_out;
wire _guard1526 = _guard1524 & _guard1525;
wire _guard1527 = fsm_out == 1'd0;
wire _guard1528 = _guard1526 & _guard1527;
wire _guard1529 = _guard1523 | _guard1528;
wire _guard1530 = early_reset_static_par0_go_out;
wire _guard1531 = _guard1529 & _guard1530;
wire _guard1532 = cond_wire38_out;
wire _guard1533 = early_reset_static_par0_go_out;
wire _guard1534 = _guard1532 & _guard1533;
wire _guard1535 = cond_wire38_out;
wire _guard1536 = early_reset_static_par0_go_out;
wire _guard1537 = _guard1535 & _guard1536;
wire _guard1538 = cond_wire29_out;
wire _guard1539 = early_reset_static_par0_go_out;
wire _guard1540 = _guard1538 & _guard1539;
wire _guard1541 = cond_wire29_out;
wire _guard1542 = early_reset_static_par0_go_out;
wire _guard1543 = _guard1541 & _guard1542;
wire _guard1544 = cond_wire4_out;
wire _guard1545 = early_reset_static_par0_go_out;
wire _guard1546 = _guard1544 & _guard1545;
wire _guard1547 = cond_wire4_out;
wire _guard1548 = early_reset_static_par0_go_out;
wire _guard1549 = _guard1547 & _guard1548;
wire _guard1550 = fsm0_out == 5'd0;
wire _guard1551 = early_reset_static_seq_go_out;
wire _guard1552 = _guard1550 & _guard1551;
wire _guard1553 = cond_wire14_out;
wire _guard1554 = early_reset_static_par0_go_out;
wire _guard1555 = _guard1553 & _guard1554;
wire _guard1556 = _guard1552 | _guard1555;
wire _guard1557 = cond_wire14_out;
wire _guard1558 = early_reset_static_par0_go_out;
wire _guard1559 = _guard1557 & _guard1558;
wire _guard1560 = fsm0_out == 5'd0;
wire _guard1561 = early_reset_static_seq_go_out;
wire _guard1562 = _guard1560 & _guard1561;
wire _guard1563 = early_reset_static_par0_go_out;
wire _guard1564 = early_reset_static_par0_go_out;
wire _guard1565 = early_reset_static_par0_go_out;
wire _guard1566 = early_reset_static_par0_go_out;
wire _guard1567 = early_reset_static_par0_go_out;
wire _guard1568 = ~_guard0;
wire _guard1569 = early_reset_static_par0_go_out;
wire _guard1570 = _guard1568 & _guard1569;
wire _guard1571 = ~_guard0;
wire _guard1572 = early_reset_static_par0_go_out;
wire _guard1573 = _guard1571 & _guard1572;
wire _guard1574 = early_reset_static_par0_go_out;
wire _guard1575 = early_reset_static_par0_go_out;
wire _guard1576 = early_reset_static_par0_go_out;
wire _guard1577 = early_reset_static_par0_go_out;
wire _guard1578 = early_reset_static_par0_go_out;
wire _guard1579 = early_reset_static_par0_go_out;
wire _guard1580 = ~_guard0;
wire _guard1581 = early_reset_static_par0_go_out;
wire _guard1582 = _guard1580 & _guard1581;
wire _guard1583 = early_reset_static_par0_go_out;
wire _guard1584 = ~_guard0;
wire _guard1585 = early_reset_static_par0_go_out;
wire _guard1586 = _guard1584 & _guard1585;
wire _guard1587 = cond_wire2_out;
wire _guard1588 = early_reset_static_par0_go_out;
wire _guard1589 = _guard1587 & _guard1588;
wire _guard1590 = cond_wire0_out;
wire _guard1591 = early_reset_static_par0_go_out;
wire _guard1592 = _guard1590 & _guard1591;
wire _guard1593 = fsm_out == 1'd0;
wire _guard1594 = cond_wire0_out;
wire _guard1595 = _guard1593 & _guard1594;
wire _guard1596 = fsm_out == 1'd0;
wire _guard1597 = _guard1595 & _guard1596;
wire _guard1598 = fsm_out == 1'd0;
wire _guard1599 = cond_wire2_out;
wire _guard1600 = _guard1598 & _guard1599;
wire _guard1601 = fsm_out == 1'd0;
wire _guard1602 = _guard1600 & _guard1601;
wire _guard1603 = _guard1597 | _guard1602;
wire _guard1604 = early_reset_static_par0_go_out;
wire _guard1605 = _guard1603 & _guard1604;
wire _guard1606 = fsm_out == 1'd0;
wire _guard1607 = cond_wire0_out;
wire _guard1608 = _guard1606 & _guard1607;
wire _guard1609 = fsm_out == 1'd0;
wire _guard1610 = _guard1608 & _guard1609;
wire _guard1611 = fsm_out == 1'd0;
wire _guard1612 = cond_wire2_out;
wire _guard1613 = _guard1611 & _guard1612;
wire _guard1614 = fsm_out == 1'd0;
wire _guard1615 = _guard1613 & _guard1614;
wire _guard1616 = _guard1610 | _guard1615;
wire _guard1617 = early_reset_static_par0_go_out;
wire _guard1618 = _guard1616 & _guard1617;
wire _guard1619 = fsm_out == 1'd0;
wire _guard1620 = cond_wire0_out;
wire _guard1621 = _guard1619 & _guard1620;
wire _guard1622 = fsm_out == 1'd0;
wire _guard1623 = _guard1621 & _guard1622;
wire _guard1624 = fsm_out == 1'd0;
wire _guard1625 = cond_wire2_out;
wire _guard1626 = _guard1624 & _guard1625;
wire _guard1627 = fsm_out == 1'd0;
wire _guard1628 = _guard1626 & _guard1627;
wire _guard1629 = _guard1623 | _guard1628;
wire _guard1630 = early_reset_static_par0_go_out;
wire _guard1631 = _guard1629 & _guard1630;
wire _guard1632 = cond_wire67_out;
wire _guard1633 = early_reset_static_par0_go_out;
wire _guard1634 = _guard1632 & _guard1633;
wire _guard1635 = cond_wire66_out;
wire _guard1636 = early_reset_static_par0_go_out;
wire _guard1637 = _guard1635 & _guard1636;
wire _guard1638 = fsm_out == 1'd0;
wire _guard1639 = cond_wire66_out;
wire _guard1640 = _guard1638 & _guard1639;
wire _guard1641 = fsm_out == 1'd0;
wire _guard1642 = _guard1640 & _guard1641;
wire _guard1643 = fsm_out == 1'd0;
wire _guard1644 = cond_wire67_out;
wire _guard1645 = _guard1643 & _guard1644;
wire _guard1646 = fsm_out == 1'd0;
wire _guard1647 = _guard1645 & _guard1646;
wire _guard1648 = _guard1642 | _guard1647;
wire _guard1649 = early_reset_static_par0_go_out;
wire _guard1650 = _guard1648 & _guard1649;
wire _guard1651 = fsm_out == 1'd0;
wire _guard1652 = cond_wire66_out;
wire _guard1653 = _guard1651 & _guard1652;
wire _guard1654 = fsm_out == 1'd0;
wire _guard1655 = _guard1653 & _guard1654;
wire _guard1656 = fsm_out == 1'd0;
wire _guard1657 = cond_wire67_out;
wire _guard1658 = _guard1656 & _guard1657;
wire _guard1659 = fsm_out == 1'd0;
wire _guard1660 = _guard1658 & _guard1659;
wire _guard1661 = _guard1655 | _guard1660;
wire _guard1662 = early_reset_static_par0_go_out;
wire _guard1663 = _guard1661 & _guard1662;
wire _guard1664 = fsm_out == 1'd0;
wire _guard1665 = cond_wire66_out;
wire _guard1666 = _guard1664 & _guard1665;
wire _guard1667 = fsm_out == 1'd0;
wire _guard1668 = _guard1666 & _guard1667;
wire _guard1669 = fsm_out == 1'd0;
wire _guard1670 = cond_wire67_out;
wire _guard1671 = _guard1669 & _guard1670;
wire _guard1672 = fsm_out == 1'd0;
wire _guard1673 = _guard1671 & _guard1672;
wire _guard1674 = _guard1668 | _guard1673;
wire _guard1675 = early_reset_static_par0_go_out;
wire _guard1676 = _guard1674 & _guard1675;
wire _guard1677 = cond_wire50_out;
wire _guard1678 = early_reset_static_par0_go_out;
wire _guard1679 = _guard1677 & _guard1678;
wire _guard1680 = cond_wire50_out;
wire _guard1681 = early_reset_static_par0_go_out;
wire _guard1682 = _guard1680 & _guard1681;
wire _guard1683 = cond_wire9_out;
wire _guard1684 = early_reset_static_par0_go_out;
wire _guard1685 = _guard1683 & _guard1684;
wire _guard1686 = cond_wire9_out;
wire _guard1687 = early_reset_static_par0_go_out;
wire _guard1688 = _guard1686 & _guard1687;
wire _guard1689 = early_reset_static_par0_go_out;
wire _guard1690 = early_reset_static_par0_go_out;
wire _guard1691 = early_reset_static_par0_go_out;
wire _guard1692 = early_reset_static_par0_go_out;
wire _guard1693 = early_reset_static_par0_go_out;
wire _guard1694 = early_reset_static_par0_go_out;
wire _guard1695 = early_reset_static_par0_go_out;
wire _guard1696 = early_reset_static_par0_go_out;
wire _guard1697 = early_reset_static_par0_go_out;
wire _guard1698 = early_reset_static_par0_go_out;
wire _guard1699 = early_reset_static_par0_go_out;
wire _guard1700 = early_reset_static_par0_go_out;
wire _guard1701 = early_reset_static_par0_go_out;
wire _guard1702 = ~_guard0;
wire _guard1703 = early_reset_static_par0_go_out;
wire _guard1704 = _guard1702 & _guard1703;
wire _guard1705 = early_reset_static_par0_go_out;
wire _guard1706 = ~_guard0;
wire _guard1707 = early_reset_static_par0_go_out;
wire _guard1708 = _guard1706 & _guard1707;
wire _guard1709 = early_reset_static_par0_go_out;
wire _guard1710 = ~_guard0;
wire _guard1711 = early_reset_static_par0_go_out;
wire _guard1712 = _guard1710 & _guard1711;
wire _guard1713 = early_reset_static_par0_go_out;
wire _guard1714 = ~_guard0;
wire _guard1715 = early_reset_static_par0_go_out;
wire _guard1716 = _guard1714 & _guard1715;
wire _guard1717 = ~_guard0;
wire _guard1718 = early_reset_static_par0_go_out;
wire _guard1719 = _guard1717 & _guard1718;
wire _guard1720 = early_reset_static_par0_go_out;
wire _guard1721 = ~_guard0;
wire _guard1722 = early_reset_static_par0_go_out;
wire _guard1723 = _guard1721 & _guard1722;
wire _guard1724 = early_reset_static_par0_go_out;
wire _guard1725 = early_reset_static_par0_go_out;
wire _guard1726 = ~_guard0;
wire _guard1727 = early_reset_static_par0_go_out;
wire _guard1728 = _guard1726 & _guard1727;
wire _guard1729 = early_reset_static_par0_go_out;
wire _guard1730 = early_reset_static_par0_go_out;
wire _guard1731 = early_reset_static_par0_go_out;
wire _guard1732 = ~_guard0;
wire _guard1733 = early_reset_static_par0_go_out;
wire _guard1734 = _guard1732 & _guard1733;
wire _guard1735 = early_reset_static_par0_go_out;
wire _guard1736 = early_reset_static_par0_go_out;
wire _guard1737 = early_reset_static_par0_go_out;
wire _guard1738 = early_reset_static_par0_go_out;
wire _guard1739 = early_reset_static_par0_go_out;
wire _guard1740 = early_reset_static_par0_go_out;
wire _guard1741 = cond_wire14_out;
wire _guard1742 = early_reset_static_par0_go_out;
wire _guard1743 = _guard1741 & _guard1742;
wire _guard1744 = cond_wire14_out;
wire _guard1745 = early_reset_static_par0_go_out;
wire _guard1746 = _guard1744 & _guard1745;
wire _guard1747 = cond_wire25_out;
wire _guard1748 = early_reset_static_par0_go_out;
wire _guard1749 = _guard1747 & _guard1748;
wire _guard1750 = cond_wire25_out;
wire _guard1751 = early_reset_static_par0_go_out;
wire _guard1752 = _guard1750 & _guard1751;
wire _guard1753 = cond_wire63_out;
wire _guard1754 = early_reset_static_par0_go_out;
wire _guard1755 = _guard1753 & _guard1754;
wire _guard1756 = cond_wire63_out;
wire _guard1757 = early_reset_static_par0_go_out;
wire _guard1758 = _guard1756 & _guard1757;
wire _guard1759 = fsm0_out == 5'd0;
wire _guard1760 = early_reset_static_seq_go_out;
wire _guard1761 = _guard1759 & _guard1760;
wire _guard1762 = cond_wire9_out;
wire _guard1763 = early_reset_static_par0_go_out;
wire _guard1764 = _guard1762 & _guard1763;
wire _guard1765 = _guard1761 | _guard1764;
wire _guard1766 = cond_wire9_out;
wire _guard1767 = early_reset_static_par0_go_out;
wire _guard1768 = _guard1766 & _guard1767;
wire _guard1769 = fsm0_out == 5'd0;
wire _guard1770 = early_reset_static_seq_go_out;
wire _guard1771 = _guard1769 & _guard1770;
wire _guard1772 = fsm0_out == 5'd0;
wire _guard1773 = early_reset_static_seq_go_out;
wire _guard1774 = _guard1772 & _guard1773;
wire _guard1775 = cond_wire36_out;
wire _guard1776 = early_reset_static_par0_go_out;
wire _guard1777 = _guard1775 & _guard1776;
wire _guard1778 = _guard1774 | _guard1777;
wire _guard1779 = fsm0_out == 5'd0;
wire _guard1780 = early_reset_static_seq_go_out;
wire _guard1781 = _guard1779 & _guard1780;
wire _guard1782 = cond_wire36_out;
wire _guard1783 = early_reset_static_par0_go_out;
wire _guard1784 = _guard1782 & _guard1783;
wire _guard1785 = early_reset_static_par0_go_out;
wire _guard1786 = early_reset_static_par0_go_out;
wire _guard1787 = early_reset_static_par0_go_out;
wire _guard1788 = early_reset_static_par0_go_out;
wire _guard1789 = early_reset_static_par0_go_out;
wire _guard1790 = early_reset_static_par0_go_out;
wire _guard1791 = early_reset_static_par0_go_out;
wire _guard1792 = early_reset_static_par0_go_out;
wire _guard1793 = early_reset_static_par0_go_out;
wire _guard1794 = early_reset_static_par0_go_out;
wire _guard1795 = ~_guard0;
wire _guard1796 = early_reset_static_par0_go_out;
wire _guard1797 = _guard1795 & _guard1796;
wire _guard1798 = early_reset_static_par0_go_out;
wire _guard1799 = early_reset_static_par0_go_out;
wire _guard1800 = early_reset_static_par0_go_out;
wire _guard1801 = early_reset_static_par0_go_out;
wire _guard1802 = early_reset_static_par0_go_out;
wire _guard1803 = ~_guard0;
wire _guard1804 = early_reset_static_par0_go_out;
wire _guard1805 = _guard1803 & _guard1804;
wire _guard1806 = early_reset_static_par0_go_out;
wire _guard1807 = early_reset_static_par0_go_out;
wire _guard1808 = early_reset_static_par0_go_out;
wire _guard1809 = early_reset_static_par0_go_out;
wire _guard1810 = early_reset_static_par0_go_out;
wire _guard1811 = ~_guard0;
wire _guard1812 = early_reset_static_par0_go_out;
wire _guard1813 = _guard1811 & _guard1812;
wire _guard1814 = early_reset_static_par0_go_out;
wire _guard1815 = early_reset_static_par0_go_out;
wire _guard1816 = ~_guard0;
wire _guard1817 = early_reset_static_par0_go_out;
wire _guard1818 = _guard1816 & _guard1817;
wire _guard1819 = cond_wire_out;
wire _guard1820 = early_reset_static_par0_go_out;
wire _guard1821 = _guard1819 & _guard1820;
wire _guard1822 = cond_wire_out;
wire _guard1823 = early_reset_static_par0_go_out;
wire _guard1824 = _guard1822 & _guard1823;
wire _guard1825 = cond_wire26_out;
wire _guard1826 = early_reset_static_par0_go_out;
wire _guard1827 = _guard1825 & _guard1826;
wire _guard1828 = cond_wire24_out;
wire _guard1829 = early_reset_static_par0_go_out;
wire _guard1830 = _guard1828 & _guard1829;
wire _guard1831 = fsm_out == 1'd0;
wire _guard1832 = cond_wire24_out;
wire _guard1833 = _guard1831 & _guard1832;
wire _guard1834 = fsm_out == 1'd0;
wire _guard1835 = _guard1833 & _guard1834;
wire _guard1836 = fsm_out == 1'd0;
wire _guard1837 = cond_wire26_out;
wire _guard1838 = _guard1836 & _guard1837;
wire _guard1839 = fsm_out == 1'd0;
wire _guard1840 = _guard1838 & _guard1839;
wire _guard1841 = _guard1835 | _guard1840;
wire _guard1842 = early_reset_static_par0_go_out;
wire _guard1843 = _guard1841 & _guard1842;
wire _guard1844 = fsm_out == 1'd0;
wire _guard1845 = cond_wire24_out;
wire _guard1846 = _guard1844 & _guard1845;
wire _guard1847 = fsm_out == 1'd0;
wire _guard1848 = _guard1846 & _guard1847;
wire _guard1849 = fsm_out == 1'd0;
wire _guard1850 = cond_wire26_out;
wire _guard1851 = _guard1849 & _guard1850;
wire _guard1852 = fsm_out == 1'd0;
wire _guard1853 = _guard1851 & _guard1852;
wire _guard1854 = _guard1848 | _guard1853;
wire _guard1855 = early_reset_static_par0_go_out;
wire _guard1856 = _guard1854 & _guard1855;
wire _guard1857 = fsm_out == 1'd0;
wire _guard1858 = cond_wire24_out;
wire _guard1859 = _guard1857 & _guard1858;
wire _guard1860 = fsm_out == 1'd0;
wire _guard1861 = _guard1859 & _guard1860;
wire _guard1862 = fsm_out == 1'd0;
wire _guard1863 = cond_wire26_out;
wire _guard1864 = _guard1862 & _guard1863;
wire _guard1865 = fsm_out == 1'd0;
wire _guard1866 = _guard1864 & _guard1865;
wire _guard1867 = _guard1861 | _guard1866;
wire _guard1868 = early_reset_static_par0_go_out;
wire _guard1869 = _guard1867 & _guard1868;
wire _guard1870 = early_reset_static_par0_go_out;
wire _guard1871 = early_reset_static_par0_go_out;
wire _guard1872 = early_reset_static_par0_go_out;
wire _guard1873 = early_reset_static_par0_go_out;
wire _guard1874 = fsm0_out == 5'd0;
wire _guard1875 = early_reset_static_seq_go_out;
wire _guard1876 = _guard1874 & _guard1875;
wire _guard1877 = early_reset_static_par0_go_out;
wire _guard1878 = _guard1876 | _guard1877;
wire _guard1879 = early_reset_static_par0_go_out;
wire _guard1880 = fsm0_out == 5'd0;
wire _guard1881 = early_reset_static_seq_go_out;
wire _guard1882 = _guard1880 & _guard1881;
wire _guard1883 = early_reset_static_par0_go_out;
wire _guard1884 = early_reset_static_par0_go_out;
wire _guard1885 = fsm0_out == 5'd0;
wire _guard1886 = early_reset_static_seq_go_out;
wire _guard1887 = _guard1885 & _guard1886;
wire _guard1888 = early_reset_static_par0_go_out;
wire _guard1889 = _guard1887 | _guard1888;
wire _guard1890 = early_reset_static_par0_go_out;
wire _guard1891 = fsm0_out == 5'd0;
wire _guard1892 = early_reset_static_seq_go_out;
wire _guard1893 = _guard1891 & _guard1892;
wire _guard1894 = fsm0_out == 5'd0;
wire _guard1895 = early_reset_static_seq_go_out;
wire _guard1896 = _guard1894 & _guard1895;
wire _guard1897 = early_reset_static_par0_go_out;
wire _guard1898 = _guard1896 | _guard1897;
wire _guard1899 = fsm0_out == 5'd0;
wire _guard1900 = early_reset_static_seq_go_out;
wire _guard1901 = _guard1899 & _guard1900;
wire _guard1902 = early_reset_static_par0_go_out;
wire _guard1903 = fsm0_out == 5'd0;
wire _guard1904 = early_reset_static_seq_go_out;
wire _guard1905 = _guard1903 & _guard1904;
wire _guard1906 = early_reset_static_par0_go_out;
wire _guard1907 = _guard1905 | _guard1906;
wire _guard1908 = fsm0_out == 5'd0;
wire _guard1909 = early_reset_static_seq_go_out;
wire _guard1910 = _guard1908 & _guard1909;
wire _guard1911 = early_reset_static_par0_go_out;
wire _guard1912 = early_reset_static_par0_go_out;
wire _guard1913 = ~_guard0;
wire _guard1914 = early_reset_static_par0_go_out;
wire _guard1915 = _guard1913 & _guard1914;
wire _guard1916 = early_reset_static_par0_go_out;
wire _guard1917 = early_reset_static_par0_go_out;
wire _guard1918 = early_reset_static_par0_go_out;
wire _guard1919 = early_reset_static_par0_go_out;
wire _guard1920 = early_reset_static_par0_go_out;
wire _guard1921 = early_reset_static_par0_go_out;
wire _guard1922 = early_reset_static_par0_go_out;
wire _guard1923 = ~_guard0;
wire _guard1924 = early_reset_static_par0_go_out;
wire _guard1925 = _guard1923 & _guard1924;
wire _guard1926 = early_reset_static_par0_go_out;
wire _guard1927 = ~_guard0;
wire _guard1928 = early_reset_static_par0_go_out;
wire _guard1929 = _guard1927 & _guard1928;
wire _guard1930 = early_reset_static_par0_go_out;
wire _guard1931 = early_reset_static_par0_go_out;
wire _guard1932 = ~_guard0;
wire _guard1933 = early_reset_static_par0_go_out;
wire _guard1934 = _guard1932 & _guard1933;
wire _guard1935 = early_reset_static_par0_go_out;
wire _guard1936 = cond_wire1_out;
wire _guard1937 = early_reset_static_par0_go_out;
wire _guard1938 = _guard1936 & _guard1937;
wire _guard1939 = cond_wire1_out;
wire _guard1940 = early_reset_static_par0_go_out;
wire _guard1941 = _guard1939 & _guard1940;
wire _guard1942 = cond_wire47_out;
wire _guard1943 = early_reset_static_par0_go_out;
wire _guard1944 = _guard1942 & _guard1943;
wire _guard1945 = cond_wire45_out;
wire _guard1946 = early_reset_static_par0_go_out;
wire _guard1947 = _guard1945 & _guard1946;
wire _guard1948 = fsm_out == 1'd0;
wire _guard1949 = cond_wire45_out;
wire _guard1950 = _guard1948 & _guard1949;
wire _guard1951 = fsm_out == 1'd0;
wire _guard1952 = _guard1950 & _guard1951;
wire _guard1953 = fsm_out == 1'd0;
wire _guard1954 = cond_wire47_out;
wire _guard1955 = _guard1953 & _guard1954;
wire _guard1956 = fsm_out == 1'd0;
wire _guard1957 = _guard1955 & _guard1956;
wire _guard1958 = _guard1952 | _guard1957;
wire _guard1959 = early_reset_static_par0_go_out;
wire _guard1960 = _guard1958 & _guard1959;
wire _guard1961 = fsm_out == 1'd0;
wire _guard1962 = cond_wire45_out;
wire _guard1963 = _guard1961 & _guard1962;
wire _guard1964 = fsm_out == 1'd0;
wire _guard1965 = _guard1963 & _guard1964;
wire _guard1966 = fsm_out == 1'd0;
wire _guard1967 = cond_wire47_out;
wire _guard1968 = _guard1966 & _guard1967;
wire _guard1969 = fsm_out == 1'd0;
wire _guard1970 = _guard1968 & _guard1969;
wire _guard1971 = _guard1965 | _guard1970;
wire _guard1972 = early_reset_static_par0_go_out;
wire _guard1973 = _guard1971 & _guard1972;
wire _guard1974 = fsm_out == 1'd0;
wire _guard1975 = cond_wire45_out;
wire _guard1976 = _guard1974 & _guard1975;
wire _guard1977 = fsm_out == 1'd0;
wire _guard1978 = _guard1976 & _guard1977;
wire _guard1979 = fsm_out == 1'd0;
wire _guard1980 = cond_wire47_out;
wire _guard1981 = _guard1979 & _guard1980;
wire _guard1982 = fsm_out == 1'd0;
wire _guard1983 = _guard1981 & _guard1982;
wire _guard1984 = _guard1978 | _guard1983;
wire _guard1985 = early_reset_static_par0_go_out;
wire _guard1986 = _guard1984 & _guard1985;
wire _guard1987 = cond_wire36_out;
wire _guard1988 = early_reset_static_par0_go_out;
wire _guard1989 = _guard1987 & _guard1988;
wire _guard1990 = cond_wire36_out;
wire _guard1991 = early_reset_static_par0_go_out;
wire _guard1992 = _guard1990 & _guard1991;
wire _guard1993 = early_reset_static_par0_go_out;
wire _guard1994 = early_reset_static_par0_go_out;
wire _guard1995 = early_reset_static_par0_go_out;
wire _guard1996 = early_reset_static_par0_go_out;
wire _guard1997 = fsm0_out == 5'd0;
wire _guard1998 = early_reset_static_seq_go_out;
wire _guard1999 = _guard1997 & _guard1998;
wire _guard2000 = early_reset_static_par0_go_out;
wire _guard2001 = _guard1999 | _guard2000;
wire _guard2002 = fsm0_out == 5'd0;
wire _guard2003 = early_reset_static_seq_go_out;
wire _guard2004 = _guard2002 & _guard2003;
wire _guard2005 = early_reset_static_par0_go_out;
wire _guard2006 = early_reset_static_par0_go_out;
wire _guard2007 = early_reset_static_par0_go_out;
wire _guard2008 = early_reset_static_par0_go_out;
wire _guard2009 = ~_guard0;
wire _guard2010 = early_reset_static_par0_go_out;
wire _guard2011 = _guard2009 & _guard2010;
wire _guard2012 = ~_guard0;
wire _guard2013 = early_reset_static_par0_go_out;
wire _guard2014 = _guard2012 & _guard2013;
wire _guard2015 = early_reset_static_par0_go_out;
wire _guard2016 = early_reset_static_par0_go_out;
wire _guard2017 = early_reset_static_par0_go_out;
wire _guard2018 = early_reset_static_par0_go_out;
wire _guard2019 = early_reset_static_par0_go_out;
wire _guard2020 = ~_guard0;
wire _guard2021 = early_reset_static_par0_go_out;
wire _guard2022 = _guard2020 & _guard2021;
wire _guard2023 = early_reset_static_par0_go_out;
wire _guard2024 = early_reset_static_par0_go_out;
wire _guard2025 = early_reset_static_par0_go_out;
assign t3_add_left = 3'd1;
assign t3_add_right = t3_idx_out;
assign l1_add_left = 3'd1;
assign l1_add_right = l1_idx_out;
assign idx_between_3_7_reg_write_en = _guard17;
assign idx_between_3_7_reg_clk = clk;
assign idx_between_3_7_reg_reset = reset;
assign idx_between_3_7_reg_in =
  _guard18 ? idx_between_3_7_comb_out :
  _guard21 ? 1'd0 :
  'x;
assign idx_between_0_4_reg_write_en = _guard26;
assign idx_between_0_4_reg_clk = clk;
assign idx_between_0_4_reg_reset = reset;
assign idx_between_0_4_reg_in =
  _guard29 ? 1'd1 :
  _guard30 ? index_lt_4_out :
  'x;
assign index_lt_5_left = idx_add_out;
assign index_lt_5_right = 5'd5;
assign index_ge_15_left = idx_add_out;
assign index_ge_15_right = 5'd15;
assign cond_wire3_in =
  _guard37 ? cond3_out :
  _guard38 ? idx_between_9_10_reg_out :
  1'd0;
assign cond_wire30_in =
  _guard41 ? cond30_out :
  _guard42 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire38_in =
  _guard43 ? idx_between_3_7_reg_out :
  _guard46 ? cond38_out :
  1'd0;
assign cond_wire39_in =
  _guard47 ? idx_between_7_11_reg_out :
  _guard50 ? cond39_out :
  1'd0;
assign cond_wire47_in =
  _guard53 ? cond47_out :
  _guard54 ? idx_between_9_13_reg_out :
  1'd0;
assign cond53_write_en = _guard55;
assign cond53_clk = clk;
assign cond53_reset = reset;
assign cond53_in =
  _guard56 ? idx_between_3_7_reg_out :
  1'd0;
assign cond_wire54_in =
  _guard57 ? idx_between_4_8_reg_out :
  _guard60 ? cond54_out :
  1'd0;
assign cond65_write_en = _guard61;
assign cond65_clk = clk;
assign cond65_reset = reset;
assign cond65_in =
  _guard62 ? idx_between_14_15_reg_out :
  1'd0;
assign left_0_3_write_en = _guard65;
assign left_0_3_clk = clk;
assign left_0_3_reset = reset;
assign left_0_3_in = left_0_2_out;
assign top_1_0_write_en = _guard71;
assign top_1_0_clk = clk;
assign top_1_0_reset = reset;
assign top_1_0_in = top_0_0_out;
assign pe_1_2_mul_ready =
  _guard77 ? 1'd1 :
  _guard80 ? 1'd0 :
  1'd0;
assign pe_1_2_clk = clk;
assign pe_1_2_top =
  _guard93 ? top_1_2_out :
  32'd0;
assign pe_1_2_left =
  _guard106 ? left_1_2_out :
  32'd0;
assign pe_1_2_reset = reset;
assign pe_1_2_go = _guard119;
assign pe_1_3_mul_ready =
  _guard122 ? 1'd1 :
  _guard125 ? 1'd0 :
  1'd0;
assign pe_1_3_clk = clk;
assign pe_1_3_top =
  _guard138 ? top_1_3_out :
  32'd0;
assign pe_1_3_left =
  _guard151 ? left_1_3_out :
  32'd0;
assign pe_1_3_reset = reset;
assign pe_1_3_go = _guard164;
assign left_1_3_write_en = _guard167;
assign left_1_3_clk = clk;
assign left_1_3_reset = reset;
assign left_1_3_in = left_1_2_out;
assign l3_idx_write_en = _guard177;
assign l3_idx_clk = clk;
assign l3_idx_reset = reset;
assign l3_idx_in =
  _guard180 ? l3_add_out :
  _guard183 ? 3'd0 :
  'x;
assign index_lt_13_left = idx_add_out;
assign index_lt_13_right = 5'd13;
assign index_ge_8_left = idx_add_out;
assign index_ge_8_right = 5'd8;
assign index_ge_14_left = idx_add_out;
assign index_ge_14_right = 5'd14;
assign idx_between_15_16_reg_write_en = _guard194;
assign idx_between_15_16_reg_clk = clk;
assign idx_between_15_16_reg_reset = reset;
assign idx_between_15_16_reg_in =
  _guard195 ? idx_between_15_16_comb_out :
  _guard198 ? 1'd0 :
  'x;
assign idx_between_6_10_reg_write_en = _guard203;
assign idx_between_6_10_reg_clk = clk;
assign idx_between_6_10_reg_reset = reset;
assign idx_between_6_10_reg_in =
  _guard204 ? idx_between_6_10_comb_out :
  _guard207 ? 1'd0 :
  'x;
assign done = _guard208;
assign t2_addr0 =
  _guard211 ? t2_idx_out :
  3'd0;
assign t3_reset = reset;
assign t0_reset = reset;
assign out_mem_2_reset = reset;
assign t2_clk = clk;
assign l0_addr0 =
  _guard214 ? l0_idx_out :
  3'd0;
assign l3_clk = clk;
assign out_mem_1_addr0 =
  _guard217 ? 3'd2 :
  _guard220 ? 3'd0 :
  _guard223 ? 3'd1 :
  _guard226 ? 3'd3 :
  3'd0;
assign out_mem_1_clk = clk;
assign out_mem_3_reset = reset;
assign out_mem_0_write_data =
  _guard229 ? pe_0_1_out :
  _guard232 ? pe_0_3_out :
  _guard235 ? pe_0_2_out :
  _guard238 ? pe_0_0_out :
  32'd0;
assign t0_clk = clk;
assign out_mem_1_reset = reset;
assign out_mem_3_write_data =
  _guard241 ? pe_3_2_out :
  _guard244 ? pe_3_0_out :
  _guard247 ? pe_3_1_out :
  _guard250 ? pe_3_3_out :
  32'd0;
assign l0_reset = reset;
assign l1_addr0 =
  _guard253 ? l1_idx_out :
  3'd0;
assign out_mem_0_clk = clk;
assign t1_reset = reset;
assign out_mem_3_clk = clk;
assign l3_addr0 =
  _guard256 ? l3_idx_out :
  3'd0;
assign out_mem_2_write_data =
  _guard259 ? pe_2_1_out :
  _guard262 ? pe_2_3_out :
  _guard265 ? pe_2_0_out :
  _guard268 ? pe_2_2_out :
  32'd0;
assign out_mem_0_reset = reset;
assign out_mem_1_write_data =
  _guard271 ? pe_1_2_out :
  _guard274 ? pe_1_3_out :
  _guard277 ? pe_1_0_out :
  _guard280 ? pe_1_1_out :
  32'd0;
assign out_mem_1_write_en = _guard305;
assign t0_addr0 =
  _guard308 ? t0_idx_out :
  3'd0;
assign t1_addr0 =
  _guard311 ? t1_idx_out :
  3'd0;
assign t1_clk = clk;
assign l1_reset = reset;
assign l2_clk = clk;
assign l2_reset = reset;
assign out_mem_0_write_en = _guard336;
assign out_mem_2_write_en = _guard361;
assign out_mem_2_clk = clk;
assign t3_clk = clk;
assign out_mem_3_write_en = _guard386;
assign l0_clk = clk;
assign l1_clk = clk;
assign l2_addr0 =
  _guard389 ? l2_idx_out :
  3'd0;
assign l3_reset = reset;
assign out_mem_0_addr0 =
  _guard392 ? 3'd2 :
  _guard395 ? 3'd0 :
  _guard398 ? 3'd1 :
  _guard401 ? 3'd3 :
  3'd0;
assign out_mem_3_addr0 =
  _guard404 ? 3'd2 :
  _guard407 ? 3'd0 :
  _guard410 ? 3'd1 :
  _guard413 ? 3'd3 :
  3'd0;
assign t2_reset = reset;
assign t3_addr0 =
  _guard416 ? t3_idx_out :
  3'd0;
assign out_mem_2_addr0 =
  _guard419 ? 3'd2 :
  _guard422 ? 3'd0 :
  _guard425 ? 3'd1 :
  _guard428 ? 3'd3 :
  3'd0;
assign cond_wire0_in =
  _guard429 ? idx_between_1_5_reg_out :
  _guard432 ? cond0_out :
  1'd0;
assign cond_wire4_in =
  _guard433 ? idx_between_1_5_reg_out :
  _guard436 ? cond4_out :
  1'd0;
assign cond6_write_en = _guard437;
assign cond6_clk = clk;
assign cond6_reset = reset;
assign cond6_in =
  _guard438 ? idx_between_2_6_reg_out :
  1'd0;
assign cond_wire13_in =
  _guard441 ? cond13_out :
  _guard442 ? idx_between_11_12_reg_out :
  1'd0;
assign cond_wire16_in =
  _guard443 ? idx_between_4_8_reg_out :
  _guard446 ? cond16_out :
  1'd0;
assign cond30_write_en = _guard447;
assign cond30_clk = clk;
assign cond30_reset = reset;
assign cond30_in =
  _guard448 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire32_in =
  _guard449 ? idx_between_5_9_reg_out :
  _guard452 ? cond32_out :
  1'd0;
assign cond_wire40_in =
  _guard455 ? cond40_out :
  _guard456 ? idx_between_11_12_reg_out :
  1'd0;
assign cond44_write_en = _guard457;
assign cond44_clk = clk;
assign cond44_reset = reset;
assign cond44_in =
  _guard458 ? idx_between_12_13_reg_out :
  1'd0;
assign cond45_write_en = _guard459;
assign cond45_clk = clk;
assign cond45_reset = reset;
assign cond45_in =
  _guard460 ? idx_between_5_9_reg_out :
  1'd0;
assign fsm_write_en = _guard461;
assign fsm_clk = clk;
assign fsm_reset = reset;
assign fsm_in =
  _guard464 ? 1'd0 :
  _guard467 ? adder0_out :
  1'd0;
assign adder_left =
  _guard468 ? fsm0_out :
  5'd0;
assign adder_right =
  _guard469 ? 5'd1 :
  5'd0;
assign early_reset_static_par0_go_in = _guard474;
assign l0_idx_write_en = _guard481;
assign l0_idx_clk = clk;
assign l0_idx_reset = reset;
assign l0_idx_in =
  _guard484 ? l0_add_out :
  _guard487 ? 3'd0 :
  'x;
assign idx_between_13_14_reg_write_en = _guard492;
assign idx_between_13_14_reg_clk = clk;
assign idx_between_13_14_reg_reset = reset;
assign idx_between_13_14_reg_in =
  _guard493 ? idx_between_13_14_comb_out :
  _guard496 ? 1'd0 :
  'x;
assign index_lt_11_left = idx_add_out;
assign index_lt_11_right = 5'd11;
assign idx_between_15_16_comb_left = index_ge_15_out;
assign idx_between_15_16_comb_right = index_lt_16_out;
assign idx_between_7_11_reg_write_en = _guard505;
assign idx_between_7_11_reg_clk = clk;
assign idx_between_7_11_reg_reset = reset;
assign idx_between_7_11_reg_in =
  _guard508 ? 1'd0 :
  _guard509 ? idx_between_7_11_comb_out :
  'x;
assign cond11_write_en = _guard510;
assign cond11_clk = clk;
assign cond11_reset = reset;
assign cond11_in =
  _guard511 ? idx_between_3_7_reg_out :
  1'd0;
assign cond15_write_en = _guard512;
assign cond15_clk = clk;
assign cond15_reset = reset;
assign cond15_in =
  _guard513 ? idx_between_4_8_reg_out :
  1'd0;
assign cond_wire27_in =
  _guard516 ? cond27_out :
  _guard517 ? idx_between_11_12_reg_out :
  1'd0;
assign cond43_write_en = _guard518;
assign cond43_clk = clk;
assign cond43_reset = reset;
assign cond43_in =
  _guard519 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire43_in =
  _guard522 ? cond43_out :
  _guard523 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire44_in =
  _guard526 ? cond44_out :
  _guard527 ? idx_between_12_13_reg_out :
  1'd0;
assign cond62_write_en = _guard528;
assign cond62_clk = clk;
assign cond62_reset = reset;
assign cond62_in =
  _guard529 ? idx_between_6_10_reg_out :
  1'd0;
assign cond_wire63_in =
  _guard530 ? idx_between_6_10_reg_out :
  _guard533 ? cond63_out :
  1'd0;
assign cond_wire67_in =
  _guard536 ? cond67_out :
  _guard537 ? idx_between_11_15_reg_out :
  1'd0;
assign pe_0_1_mul_ready =
  _guard540 ? 1'd1 :
  _guard543 ? 1'd0 :
  1'd0;
assign pe_0_1_clk = clk;
assign pe_0_1_top =
  _guard556 ? top_0_1_out :
  32'd0;
assign pe_0_1_left =
  _guard569 ? left_0_1_out :
  32'd0;
assign pe_0_1_reset = reset;
assign pe_0_1_go = _guard582;
assign left_1_2_write_en = _guard585;
assign left_1_2_clk = clk;
assign left_1_2_reset = reset;
assign left_1_2_in = left_1_1_out;
assign left_2_2_write_en = _guard591;
assign left_2_2_clk = clk;
assign left_2_2_reset = reset;
assign left_2_2_in = left_2_1_out;
assign l3_add_left = 3'd1;
assign l3_add_right = l3_idx_out;
assign index_ge_3_left = idx_add_out;
assign index_ge_3_right = 5'd3;
assign index_ge_12_left = idx_add_out;
assign index_ge_12_right = 5'd12;
assign idx_between_4_8_reg_write_en = _guard609;
assign idx_between_4_8_reg_clk = clk;
assign idx_between_4_8_reg_reset = reset;
assign idx_between_4_8_reg_in =
  _guard612 ? 1'd0 :
  _guard613 ? idx_between_4_8_comb_out :
  'x;
assign idx_between_5_9_comb_left = index_ge_5_out;
assign idx_between_5_9_comb_right = index_lt_9_out;
assign idx_between_9_13_comb_left = index_ge_9_out;
assign idx_between_9_13_comb_right = index_lt_13_out;
assign idx_between_10_14_comb_left = index_ge_10_out;
assign idx_between_10_14_comb_right = index_lt_14_out;
assign idx_between_6_10_comb_left = index_ge_6_out;
assign idx_between_6_10_comb_right = index_lt_10_out;
assign cond_write_en = _guard622;
assign cond_clk = clk;
assign cond_reset = reset;
assign cond_in =
  _guard623 ? idx_between_0_4_reg_out :
  1'd0;
assign cond_wire26_in =
  _guard624 ? idx_between_7_11_reg_out :
  _guard627 ? cond26_out :
  1'd0;
assign cond35_write_en = _guard628;
assign cond35_clk = clk;
assign cond35_reset = reset;
assign cond35_in =
  _guard629 ? idx_between_13_14_reg_out :
  1'd0;
assign cond_wire35_in =
  _guard630 ? idx_between_13_14_reg_out :
  _guard633 ? cond35_out :
  1'd0;
assign cond_wire50_in =
  _guard634 ? idx_between_6_10_reg_out :
  _guard637 ? cond50_out :
  1'd0;
assign cond_wire56_in =
  _guard638 ? idx_between_8_12_reg_out :
  _guard641 ? cond56_out :
  1'd0;
assign cond60_write_en = _guard642;
assign cond60_clk = clk;
assign cond60_reset = reset;
assign cond60_in =
  _guard643 ? idx_between_9_13_reg_out :
  1'd0;
assign pe_1_0_mul_ready =
  _guard646 ? 1'd1 :
  _guard649 ? 1'd0 :
  1'd0;
assign pe_1_0_clk = clk;
assign pe_1_0_top =
  _guard662 ? top_1_0_out :
  32'd0;
assign pe_1_0_left =
  _guard675 ? left_1_0_out :
  32'd0;
assign pe_1_0_reset = reset;
assign pe_1_0_go = _guard688;
assign left_1_0_write_en = _guard691;
assign left_1_0_clk = clk;
assign left_1_0_reset = reset;
assign left_1_0_in = l1_read_data;
assign left_1_1_write_en = _guard697;
assign left_1_1_clk = clk;
assign left_1_1_reset = reset;
assign left_1_1_in = left_1_0_out;
assign top_1_2_write_en = _guard703;
assign top_1_2_clk = clk;
assign top_1_2_reset = reset;
assign top_1_2_in = top_0_2_out;
assign left_2_0_write_en = _guard709;
assign left_2_0_clk = clk;
assign left_2_0_reset = reset;
assign left_2_0_in = l2_read_data;
assign left_3_1_write_en = _guard715;
assign left_3_1_clk = clk;
assign left_3_1_reset = reset;
assign left_3_1_in = left_3_0_out;
assign pe_3_2_mul_ready =
  _guard721 ? 1'd1 :
  _guard724 ? 1'd0 :
  1'd0;
assign pe_3_2_clk = clk;
assign pe_3_2_top =
  _guard737 ? top_3_2_out :
  32'd0;
assign pe_3_2_left =
  _guard750 ? left_3_2_out :
  32'd0;
assign pe_3_2_reset = reset;
assign pe_3_2_go = _guard763;
assign t1_idx_write_en = _guard770;
assign t1_idx_clk = clk;
assign t1_idx_reset = reset;
assign t1_idx_in =
  _guard773 ? t1_add_out :
  _guard776 ? 3'd0 :
  'x;
assign cond18_write_en = _guard777;
assign cond18_clk = clk;
assign cond18_reset = reset;
assign cond18_in =
  _guard778 ? idx_between_12_13_reg_out :
  1'd0;
assign cond_wire24_in =
  _guard779 ? idx_between_3_7_reg_out :
  _guard782 ? cond24_out :
  1'd0;
assign cond_wire31_in =
  _guard783 ? idx_between_12_13_reg_out :
  _guard786 ? cond31_out :
  1'd0;
assign cond_wire46_in =
  _guard787 ? idx_between_5_9_reg_out :
  _guard790 ? cond46_out :
  1'd0;
assign cond_wire48_in =
  _guard791 ? idx_between_13_14_reg_out :
  _guard794 ? cond48_out :
  1'd0;
assign left_0_0_write_en = _guard797;
assign left_0_0_clk = clk;
assign left_0_0_reset = reset;
assign left_0_0_in = l0_read_data;
assign pe_0_3_mul_ready =
  _guard803 ? 1'd1 :
  _guard806 ? 1'd0 :
  1'd0;
assign pe_0_3_clk = clk;
assign pe_0_3_top =
  _guard819 ? top_0_3_out :
  32'd0;
assign pe_0_3_left =
  _guard832 ? left_0_3_out :
  32'd0;
assign pe_0_3_reset = reset;
assign pe_0_3_go = _guard845;
assign top_1_3_write_en = _guard848;
assign top_1_3_clk = clk;
assign top_1_3_reset = reset;
assign top_1_3_in = top_0_3_out;
assign left_2_3_write_en = _guard854;
assign left_2_3_clk = clk;
assign left_2_3_reset = reset;
assign left_2_3_in = left_2_2_out;
assign pe_3_0_mul_ready =
  _guard860 ? 1'd1 :
  _guard863 ? 1'd0 :
  1'd0;
assign pe_3_0_clk = clk;
assign pe_3_0_top =
  _guard876 ? top_3_0_out :
  32'd0;
assign pe_3_0_left =
  _guard889 ? left_3_0_out :
  32'd0;
assign pe_3_0_reset = reset;
assign pe_3_0_go = _guard902;
assign top_3_2_write_en = _guard905;
assign top_3_2_clk = clk;
assign top_3_2_reset = reset;
assign top_3_2_in = top_2_2_out;
assign idx_between_14_15_comb_left = index_ge_14_out;
assign idx_between_14_15_comb_right = index_lt_15_out;
assign idx_between_9_10_comb_left = index_ge_9_out;
assign idx_between_9_10_comb_right = index_lt_10_out;
assign idx_between_10_11_comb_left = index_ge_10_out;
assign idx_between_10_11_comb_right = index_lt_11_out;
assign cond_wire18_in =
  _guard917 ? cond18_out :
  _guard918 ? idx_between_12_13_reg_out :
  1'd0;
assign cond19_write_en = _guard919;
assign cond19_clk = clk;
assign cond19_reset = reset;
assign cond19_in =
  _guard920 ? idx_between_1_5_reg_out :
  1'd0;
assign cond_wire29_in =
  _guard921 ? idx_between_4_8_reg_out :
  _guard924 ? cond29_out :
  1'd0;
assign cond34_write_en = _guard925;
assign cond34_clk = clk;
assign cond34_reset = reset;
assign cond34_in =
  _guard926 ? idx_between_9_13_reg_out :
  1'd0;
assign cond40_write_en = _guard927;
assign cond40_clk = clk;
assign cond40_reset = reset;
assign cond40_in =
  _guard928 ? idx_between_11_12_reg_out :
  1'd0;
assign cond57_write_en = _guard929;
assign cond57_clk = clk;
assign cond57_reset = reset;
assign cond57_in =
  _guard930 ? idx_between_12_13_reg_out :
  1'd0;
assign cond_wire59_in =
  _guard931 ? idx_between_5_9_reg_out :
  _guard934 ? cond59_out :
  1'd0;
assign cond_wire61_in =
  _guard935 ? idx_between_13_14_reg_out :
  _guard938 ? cond61_out :
  1'd0;
assign pe_0_2_mul_ready =
  _guard941 ? 1'd1 :
  _guard944 ? 1'd0 :
  1'd0;
assign pe_0_2_clk = clk;
assign pe_0_2_top =
  _guard957 ? top_0_2_out :
  32'd0;
assign pe_0_2_left =
  _guard970 ? left_0_2_out :
  32'd0;
assign pe_0_2_reset = reset;
assign pe_0_2_go = _guard983;
assign t0_idx_write_en = _guard990;
assign t0_idx_clk = clk;
assign t0_idx_reset = reset;
assign t0_idx_in =
  _guard993 ? t0_add_out :
  _guard996 ? 3'd0 :
  'x;
assign l1_idx_write_en = _guard1003;
assign l1_idx_clk = clk;
assign l1_idx_reset = reset;
assign l1_idx_in =
  _guard1006 ? l1_add_out :
  _guard1009 ? 3'd0 :
  'x;
assign idx_add_left = idx_out;
assign idx_add_right = 5'd1;
assign idx_between_8_12_reg_write_en = _guard1016;
assign idx_between_8_12_reg_clk = clk;
assign idx_between_8_12_reg_reset = reset;
assign idx_between_8_12_reg_in =
  _guard1019 ? 1'd0 :
  _guard1020 ? idx_between_8_12_comb_out :
  'x;
assign index_lt_16_left = idx_add_out;
assign index_lt_16_right = 5'd16;
assign index_ge_7_left = idx_add_out;
assign index_ge_7_right = 5'd7;
assign cond3_write_en = _guard1025;
assign cond3_clk = clk;
assign cond3_reset = reset;
assign cond3_in =
  _guard1026 ? idx_between_9_10_reg_out :
  1'd0;
assign cond13_write_en = _guard1027;
assign cond13_clk = clk;
assign cond13_reset = reset;
assign cond13_in =
  _guard1028 ? idx_between_11_12_reg_out :
  1'd0;
assign cond29_write_en = _guard1029;
assign cond29_clk = clk;
assign cond29_reset = reset;
assign cond29_in =
  _guard1030 ? idx_between_4_8_reg_out :
  1'd0;
assign cond41_write_en = _guard1031;
assign cond41_clk = clk;
assign cond41_reset = reset;
assign cond41_in =
  _guard1032 ? idx_between_4_8_reg_out :
  1'd0;
assign cond54_write_en = _guard1033;
assign cond54_clk = clk;
assign cond54_reset = reset;
assign cond54_in =
  _guard1034 ? idx_between_4_8_reg_out :
  1'd0;
assign cond64_write_en = _guard1035;
assign cond64_clk = clk;
assign cond64_reset = reset;
assign cond64_in =
  _guard1036 ? idx_between_10_14_reg_out :
  1'd0;
assign cond67_write_en = _guard1037;
assign cond67_clk = clk;
assign cond67_reset = reset;
assign cond67_in =
  _guard1038 ? idx_between_11_15_reg_out :
  1'd0;
assign cond68_write_en = _guard1039;
assign cond68_clk = clk;
assign cond68_reset = reset;
assign cond68_in =
  _guard1040 ? idx_between_15_16_reg_out :
  1'd0;
assign early_reset_static_par0_done_in = ud0_out;
assign pe_2_1_mul_ready =
  _guard1043 ? 1'd1 :
  _guard1046 ? 1'd0 :
  1'd0;
assign pe_2_1_clk = clk;
assign pe_2_1_top =
  _guard1059 ? top_2_1_out :
  32'd0;
assign pe_2_1_left =
  _guard1072 ? left_2_1_out :
  32'd0;
assign pe_2_1_reset = reset;
assign pe_2_1_go = _guard1085;
assign pe_2_3_mul_ready =
  _guard1088 ? 1'd1 :
  _guard1091 ? 1'd0 :
  1'd0;
assign pe_2_3_clk = clk;
assign pe_2_3_top =
  _guard1104 ? top_2_3_out :
  32'd0;
assign pe_2_3_left =
  _guard1117 ? left_2_3_out :
  32'd0;
assign pe_2_3_reset = reset;
assign pe_2_3_go = _guard1130;
assign pe_3_1_mul_ready =
  _guard1133 ? 1'd1 :
  _guard1136 ? 1'd0 :
  1'd0;
assign pe_3_1_clk = clk;
assign pe_3_1_top =
  _guard1149 ? top_3_1_out :
  32'd0;
assign pe_3_1_left =
  _guard1162 ? left_3_1_out :
  32'd0;
assign pe_3_1_reset = reset;
assign pe_3_1_go = _guard1175;
assign cond17_write_en = _guard1176;
assign cond17_clk = clk;
assign cond17_reset = reset;
assign cond17_in =
  _guard1177 ? idx_between_8_12_reg_out :
  1'd0;
assign cond_wire22_in =
  _guard1178 ? idx_between_6_10_reg_out :
  _guard1181 ? cond22_out :
  1'd0;
assign cond23_write_en = _guard1182;
assign cond23_clk = clk;
assign cond23_reset = reset;
assign cond23_in =
  _guard1183 ? idx_between_10_11_reg_out :
  1'd0;
assign cond25_write_en = _guard1184;
assign cond25_clk = clk;
assign cond25_reset = reset;
assign cond25_in =
  _guard1185 ? idx_between_3_7_reg_out :
  1'd0;
assign cond_wire33_in =
  _guard1186 ? idx_between_5_9_reg_out :
  _guard1189 ? cond33_out :
  1'd0;
assign cond52_write_en = _guard1190;
assign cond52_clk = clk;
assign cond52_reset = reset;
assign cond52_in =
  _guard1191 ? idx_between_14_15_reg_out :
  1'd0;
assign cond56_write_en = _guard1192;
assign cond56_clk = clk;
assign cond56_reset = reset;
assign cond56_in =
  _guard1193 ? idx_between_8_12_reg_out :
  1'd0;
assign cond58_write_en = _guard1194;
assign cond58_clk = clk;
assign cond58_reset = reset;
assign cond58_in =
  _guard1195 ? idx_between_5_9_reg_out :
  1'd0;
assign fsm0_write_en = _guard1196;
assign fsm0_clk = clk;
assign fsm0_reset = reset;
assign fsm0_in =
  _guard1199 ? adder_out :
  _guard1202 ? 5'd0 :
  5'd0;
assign top_2_0_write_en = _guard1205;
assign top_2_0_clk = clk;
assign top_2_0_reset = reset;
assign top_2_0_in = top_1_0_out;
assign top_3_0_write_en = _guard1211;
assign top_3_0_clk = clk;
assign top_3_0_reset = reset;
assign top_3_0_in = top_2_0_out;
assign top_3_1_write_en = _guard1217;
assign top_3_1_clk = clk;
assign top_3_1_reset = reset;
assign top_3_1_in = top_2_1_out;
assign idx_write_en = _guard1225;
assign idx_clk = clk;
assign idx_reset = reset;
assign idx_in =
  _guard1228 ? 5'd0 :
  _guard1229 ? idx_add_out :
  'x;
assign idx_between_12_13_reg_write_en = _guard1234;
assign idx_between_12_13_reg_clk = clk;
assign idx_between_12_13_reg_reset = reset;
assign idx_between_12_13_reg_in =
  _guard1237 ? 1'd0 :
  _guard1238 ? idx_between_12_13_comb_out :
  'x;
assign idx_between_5_9_reg_write_en = _guard1243;
assign idx_between_5_9_reg_clk = clk;
assign idx_between_5_9_reg_reset = reset;
assign idx_between_5_9_reg_in =
  _guard1244 ? idx_between_5_9_comb_out :
  _guard1247 ? 1'd0 :
  'x;
assign index_lt_15_left = idx_add_out;
assign index_lt_15_right = 5'd15;
assign cond7_write_en = _guard1250;
assign cond7_clk = clk;
assign cond7_reset = reset;
assign cond7_in =
  _guard1251 ? idx_between_6_10_reg_out :
  1'd0;
assign cond_wire8_in =
  _guard1252 ? idx_between_10_11_reg_out :
  _guard1255 ? cond8_out :
  1'd0;
assign cond9_write_en = _guard1256;
assign cond9_clk = clk;
assign cond9_reset = reset;
assign cond9_in =
  _guard1257 ? idx_between_2_6_reg_out :
  1'd0;
assign cond14_write_en = _guard1258;
assign cond14_clk = clk;
assign cond14_reset = reset;
assign cond14_in =
  _guard1259 ? idx_between_3_7_reg_out :
  1'd0;
assign cond_wire20_in =
  _guard1262 ? cond20_out :
  _guard1263 ? idx_between_2_6_reg_out :
  1'd0;
assign cond27_write_en = _guard1264;
assign cond27_clk = clk;
assign cond27_reset = reset;
assign cond27_in =
  _guard1265 ? idx_between_11_12_reg_out :
  1'd0;
assign cond32_write_en = _guard1266;
assign cond32_clk = clk;
assign cond32_reset = reset;
assign cond32_in =
  _guard1267 ? idx_between_5_9_reg_out :
  1'd0;
assign cond_wire37_in =
  _guard1268 ? idx_between_3_7_reg_out :
  _guard1271 ? cond37_out :
  1'd0;
assign cond50_write_en = _guard1272;
assign cond50_clk = clk;
assign cond50_reset = reset;
assign cond50_in =
  _guard1273 ? idx_between_6_10_reg_out :
  1'd0;
assign cond_wire60_in =
  _guard1276 ? cond60_out :
  _guard1277 ? idx_between_9_13_reg_out :
  1'd0;
assign cond_wire64_in =
  _guard1280 ? cond64_out :
  _guard1281 ? idx_between_10_14_reg_out :
  1'd0;
assign wrapper_early_reset_static_seq_done_in = _guard1284;
assign top_0_1_write_en = _guard1287;
assign top_0_1_clk = clk;
assign top_0_1_reset = reset;
assign top_0_1_in = t1_read_data;
assign left_0_2_write_en = _guard1293;
assign left_0_2_clk = clk;
assign left_0_2_reset = reset;
assign left_0_2_in = left_0_1_out;
assign top_2_3_write_en = _guard1299;
assign top_2_3_clk = clk;
assign top_2_3_reset = reset;
assign top_2_3_in = top_1_3_out;
assign left_3_0_write_en = _guard1305;
assign left_3_0_clk = clk;
assign left_3_0_reset = reset;
assign left_3_0_in = l3_read_data;
assign idx_between_3_7_comb_left = index_ge_3_out;
assign idx_between_3_7_comb_right = index_lt_7_out;
assign idx_between_13_14_comb_left = index_ge_13_out;
assign idx_between_13_14_comb_right = index_lt_14_out;
assign index_lt_8_left = idx_add_out;
assign index_lt_8_right = 5'd8;
assign index_ge_4_left = idx_add_out;
assign index_ge_4_right = 5'd4;
assign index_lt_9_left = idx_add_out;
assign index_lt_9_right = 5'd9;
assign idx_between_14_15_reg_write_en = _guard1323;
assign idx_between_14_15_reg_clk = clk;
assign idx_between_14_15_reg_reset = reset;
assign idx_between_14_15_reg_in =
  _guard1324 ? idx_between_14_15_comb_out :
  _guard1327 ? 1'd0 :
  'x;
assign idx_between_9_10_reg_write_en = _guard1332;
assign idx_between_9_10_reg_clk = clk;
assign idx_between_9_10_reg_reset = reset;
assign idx_between_9_10_reg_in =
  _guard1333 ? idx_between_9_10_comb_out :
  _guard1336 ? 1'd0 :
  'x;
assign idx_between_1_5_reg_write_en = _guard1341;
assign idx_between_1_5_reg_clk = clk;
assign idx_between_1_5_reg_reset = reset;
assign idx_between_1_5_reg_in =
  _guard1344 ? 1'd0 :
  _guard1345 ? idx_between_1_5_comb_out :
  'x;
assign index_ge_1_left = idx_add_out;
assign index_ge_1_right = 5'd1;
assign index_lt_6_left = idx_add_out;
assign index_lt_6_right = 5'd6;
assign cond4_write_en = _guard1350;
assign cond4_clk = clk;
assign cond4_reset = reset;
assign cond4_in =
  _guard1351 ? idx_between_1_5_reg_out :
  1'd0;
assign cond5_write_en = _guard1352;
assign cond5_clk = clk;
assign cond5_reset = reset;
assign cond5_in =
  _guard1353 ? idx_between_2_6_reg_out :
  1'd0;
assign cond_wire6_in =
  _guard1356 ? cond6_out :
  _guard1357 ? idx_between_2_6_reg_out :
  1'd0;
assign cond20_write_en = _guard1358;
assign cond20_clk = clk;
assign cond20_reset = reset;
assign cond20_in =
  _guard1359 ? idx_between_2_6_reg_out :
  1'd0;
assign cond_wire36_in =
  _guard1362 ? cond36_out :
  _guard1363 ? idx_between_2_6_reg_out :
  1'd0;
assign cond46_write_en = _guard1364;
assign cond46_clk = clk;
assign cond46_reset = reset;
assign cond46_in =
  _guard1365 ? idx_between_5_9_reg_out :
  1'd0;
assign cond_wire62_in =
  _guard1366 ? idx_between_6_10_reg_out :
  _guard1369 ? cond62_out :
  1'd0;
assign cond63_write_en = _guard1370;
assign cond63_clk = clk;
assign cond63_reset = reset;
assign cond63_in =
  _guard1371 ? idx_between_6_10_reg_out :
  1'd0;
assign cond_wire66_in =
  _guard1372 ? idx_between_7_11_reg_out :
  _guard1375 ? cond66_out :
  1'd0;
assign adder0_left =
  _guard1376 ? fsm_out :
  1'd0;
assign adder0_right = _guard1377;
assign early_reset_static_seq_go_in = _guard1378;
assign top_0_2_write_en = _guard1381;
assign top_0_2_clk = clk;
assign top_0_2_reset = reset;
assign top_0_2_in = t2_read_data;
assign top_1_1_write_en = _guard1387;
assign top_1_1_clk = clk;
assign top_1_1_reset = reset;
assign top_1_1_in = top_0_1_out;
assign left_3_2_write_en = _guard1393;
assign left_3_2_clk = clk;
assign left_3_2_reset = reset;
assign left_3_2_in = left_3_1_out;
assign t0_add_left = 3'd1;
assign t0_add_right = t0_idx_out;
assign l0_add_left = 3'd1;
assign l0_add_right = l0_idx_out;
assign idx_between_4_8_comb_left = index_ge_4_out;
assign idx_between_4_8_comb_right = index_lt_8_out;
assign index_ge_9_left = idx_add_out;
assign index_ge_9_right = 5'd9;
assign idx_between_10_11_reg_write_en = _guard1417;
assign idx_between_10_11_reg_clk = clk;
assign idx_between_10_11_reg_reset = reset;
assign idx_between_10_11_reg_in =
  _guard1418 ? idx_between_10_11_comb_out :
  _guard1421 ? 1'd0 :
  'x;
assign index_ge_11_left = idx_add_out;
assign index_ge_11_right = 5'd11;
assign idx_between_11_15_comb_left = index_ge_11_out;
assign idx_between_11_15_comb_right = index_lt_15_out;
assign cond_wire2_in =
  _guard1426 ? idx_between_5_9_reg_out :
  _guard1429 ? cond2_out :
  1'd0;
assign cond_wire9_in =
  _guard1432 ? cond9_out :
  _guard1433 ? idx_between_2_6_reg_out :
  1'd0;
assign cond10_write_en = _guard1434;
assign cond10_clk = clk;
assign cond10_reset = reset;
assign cond10_in =
  _guard1435 ? idx_between_3_7_reg_out :
  1'd0;
assign cond_wire11_in =
  _guard1436 ? idx_between_3_7_reg_out :
  _guard1439 ? cond11_out :
  1'd0;
assign cond21_write_en = _guard1440;
assign cond21_clk = clk;
assign cond21_reset = reset;
assign cond21_in =
  _guard1441 ? idx_between_2_6_reg_out :
  1'd0;
assign cond24_write_en = _guard1442;
assign cond24_clk = clk;
assign cond24_reset = reset;
assign cond24_in =
  _guard1443 ? idx_between_3_7_reg_out :
  1'd0;
assign cond31_write_en = _guard1444;
assign cond31_clk = clk;
assign cond31_reset = reset;
assign cond31_in =
  _guard1445 ? idx_between_12_13_reg_out :
  1'd0;
assign cond36_write_en = _guard1446;
assign cond36_clk = clk;
assign cond36_reset = reset;
assign cond36_in =
  _guard1447 ? idx_between_2_6_reg_out :
  1'd0;
assign cond_wire41_in =
  _guard1448 ? idx_between_4_8_reg_out :
  _guard1451 ? cond41_out :
  1'd0;
assign cond_wire45_in =
  _guard1454 ? cond45_out :
  _guard1455 ? idx_between_5_9_reg_out :
  1'd0;
assign cond51_write_en = _guard1456;
assign cond51_clk = clk;
assign cond51_reset = reset;
assign cond51_in =
  _guard1457 ? idx_between_10_14_reg_out :
  1'd0;
assign cond_wire57_in =
  _guard1460 ? cond57_out :
  _guard1461 ? idx_between_12_13_reg_out :
  1'd0;
assign cond_wire58_in =
  _guard1464 ? cond58_out :
  _guard1465 ? idx_between_5_9_reg_out :
  1'd0;
assign cond61_write_en = _guard1466;
assign cond61_clk = clk;
assign cond61_reset = reset;
assign cond61_in =
  _guard1467 ? idx_between_13_14_reg_out :
  1'd0;
assign signal_reg_write_en = _guard1477;
assign signal_reg_clk = clk;
assign signal_reg_reset = reset;
assign signal_reg_in =
  _guard1483 ? 1'd1 :
  _guard1486 ? 1'd0 :
  1'd0;
assign pe_2_0_mul_ready =
  _guard1489 ? 1'd1 :
  _guard1492 ? 1'd0 :
  1'd0;
assign pe_2_0_clk = clk;
assign pe_2_0_top =
  _guard1505 ? top_2_0_out :
  32'd0;
assign pe_2_0_left =
  _guard1518 ? left_2_0_out :
  32'd0;
assign pe_2_0_reset = reset;
assign pe_2_0_go = _guard1531;
assign left_2_1_write_en = _guard1534;
assign left_2_1_clk = clk;
assign left_2_1_reset = reset;
assign left_2_1_in = left_2_0_out;
assign top_2_2_write_en = _guard1540;
assign top_2_2_clk = clk;
assign top_2_2_reset = reset;
assign top_2_2_in = top_1_2_out;
assign t1_add_left = 3'd1;
assign t1_add_right = t1_idx_out;
assign t3_idx_write_en = _guard1556;
assign t3_idx_clk = clk;
assign t3_idx_reset = reset;
assign t3_idx_in =
  _guard1559 ? t3_add_out :
  _guard1562 ? 3'd0 :
  'x;
assign index_lt_10_left = idx_add_out;
assign index_lt_10_right = 5'd10;
assign index_ge_2_left = idx_add_out;
assign index_ge_2_right = 5'd2;
assign cond_wire_in =
  _guard1567 ? idx_between_0_4_reg_out :
  _guard1570 ? cond_out :
  1'd0;
assign cond_wire15_in =
  _guard1573 ? cond15_out :
  _guard1574 ? idx_between_4_8_reg_out :
  1'd0;
assign cond16_write_en = _guard1575;
assign cond16_clk = clk;
assign cond16_reset = reset;
assign cond16_in =
  _guard1576 ? idx_between_4_8_reg_out :
  1'd0;
assign cond37_write_en = _guard1577;
assign cond37_clk = clk;
assign cond37_reset = reset;
assign cond37_in =
  _guard1578 ? idx_between_3_7_reg_out :
  1'd0;
assign cond_wire49_in =
  _guard1579 ? idx_between_6_10_reg_out :
  _guard1582 ? cond49_out :
  1'd0;
assign cond_wire55_in =
  _guard1583 ? idx_between_4_8_reg_out :
  _guard1586 ? cond55_out :
  1'd0;
assign pe_0_0_mul_ready =
  _guard1589 ? 1'd1 :
  _guard1592 ? 1'd0 :
  1'd0;
assign pe_0_0_clk = clk;
assign pe_0_0_top =
  _guard1605 ? top_0_0_out :
  32'd0;
assign pe_0_0_left =
  _guard1618 ? left_0_0_out :
  32'd0;
assign pe_0_0_reset = reset;
assign pe_0_0_go = _guard1631;
assign pe_3_3_mul_ready =
  _guard1634 ? 1'd1 :
  _guard1637 ? 1'd0 :
  1'd0;
assign pe_3_3_clk = clk;
assign pe_3_3_top =
  _guard1650 ? top_3_3_out :
  32'd0;
assign pe_3_3_left =
  _guard1663 ? left_3_3_out :
  32'd0;
assign pe_3_3_reset = reset;
assign pe_3_3_go = _guard1676;
assign top_3_3_write_en = _guard1679;
assign top_3_3_clk = clk;
assign top_3_3_reset = reset;
assign top_3_3_in = top_2_3_out;
assign t2_add_left = 3'd1;
assign t2_add_right = t2_idx_out;
assign idx_between_12_13_comb_left = index_ge_12_out;
assign idx_between_12_13_comb_right = index_lt_13_out;
assign index_lt_12_left = idx_add_out;
assign index_lt_12_right = 5'd12;
assign index_ge_5_left = idx_add_out;
assign index_ge_5_right = 5'd5;
assign index_ge_10_left = idx_add_out;
assign index_ge_10_right = 5'd10;
assign idx_between_7_11_comb_left = index_ge_7_out;
assign idx_between_7_11_comb_right = index_lt_11_out;
assign cond0_write_en = _guard1699;
assign cond0_clk = clk;
assign cond0_reset = reset;
assign cond0_in =
  _guard1700 ? idx_between_1_5_reg_out :
  1'd0;
assign cond_wire7_in =
  _guard1701 ? idx_between_6_10_reg_out :
  _guard1704 ? cond7_out :
  1'd0;
assign cond_wire10_in =
  _guard1705 ? idx_between_3_7_reg_out :
  _guard1708 ? cond10_out :
  1'd0;
assign cond_wire12_in =
  _guard1709 ? idx_between_7_11_reg_out :
  _guard1712 ? cond12_out :
  1'd0;
assign cond_wire17_in =
  _guard1713 ? idx_between_8_12_reg_out :
  _guard1716 ? cond17_out :
  1'd0;
assign cond_wire19_in =
  _guard1719 ? cond19_out :
  _guard1720 ? idx_between_1_5_reg_out :
  1'd0;
assign cond_wire23_in =
  _guard1723 ? cond23_out :
  _guard1724 ? idx_between_10_11_reg_out :
  1'd0;
assign cond_wire25_in =
  _guard1725 ? idx_between_3_7_reg_out :
  _guard1728 ? cond25_out :
  1'd0;
assign cond33_write_en = _guard1729;
assign cond33_clk = clk;
assign cond33_reset = reset;
assign cond33_in =
  _guard1730 ? idx_between_5_9_reg_out :
  1'd0;
assign cond_wire42_in =
  _guard1731 ? idx_between_4_8_reg_out :
  _guard1734 ? cond42_out :
  1'd0;
assign cond47_write_en = _guard1735;
assign cond47_clk = clk;
assign cond47_reset = reset;
assign cond47_in =
  _guard1736 ? idx_between_9_13_reg_out :
  1'd0;
assign cond48_write_en = _guard1737;
assign cond48_clk = clk;
assign cond48_reset = reset;
assign cond48_in =
  _guard1738 ? idx_between_13_14_reg_out :
  1'd0;
assign cond66_write_en = _guard1739;
assign cond66_clk = clk;
assign cond66_reset = reset;
assign cond66_in =
  _guard1740 ? idx_between_7_11_reg_out :
  1'd0;
assign early_reset_static_seq_done_in = ud_out;
assign top_0_3_write_en = _guard1743;
assign top_0_3_clk = clk;
assign top_0_3_reset = reset;
assign top_0_3_in = t3_read_data;
assign top_2_1_write_en = _guard1749;
assign top_2_1_clk = clk;
assign top_2_1_reset = reset;
assign top_2_1_in = top_1_1_out;
assign left_3_3_write_en = _guard1755;
assign left_3_3_clk = clk;
assign left_3_3_reset = reset;
assign left_3_3_in = left_3_2_out;
assign t2_idx_write_en = _guard1765;
assign t2_idx_clk = clk;
assign t2_idx_reset = reset;
assign t2_idx_in =
  _guard1768 ? t2_add_out :
  _guard1771 ? 3'd0 :
  'x;
assign l2_idx_write_en = _guard1778;
assign l2_idx_clk = clk;
assign l2_idx_reset = reset;
assign l2_idx_in =
  _guard1781 ? 3'd0 :
  _guard1784 ? l2_add_out :
  'x;
assign index_lt_7_left = idx_add_out;
assign index_lt_7_right = 5'd7;
assign index_ge_6_left = idx_add_out;
assign index_ge_6_right = 5'd6;
assign idx_between_11_12_comb_left = index_ge_11_out;
assign idx_between_11_12_comb_right = index_lt_12_out;
assign cond1_write_en = _guard1791;
assign cond1_clk = clk;
assign cond1_reset = reset;
assign cond1_in =
  _guard1792 ? idx_between_1_5_reg_out :
  1'd0;
assign cond2_write_en = _guard1793;
assign cond2_clk = clk;
assign cond2_reset = reset;
assign cond2_in =
  _guard1794 ? idx_between_5_9_reg_out :
  1'd0;
assign cond_wire5_in =
  _guard1797 ? cond5_out :
  _guard1798 ? idx_between_2_6_reg_out :
  1'd0;
assign cond22_write_en = _guard1799;
assign cond22_clk = clk;
assign cond22_reset = reset;
assign cond22_in =
  _guard1800 ? idx_between_6_10_reg_out :
  1'd0;
assign cond26_write_en = _guard1801;
assign cond26_clk = clk;
assign cond26_reset = reset;
assign cond26_in =
  _guard1802 ? idx_between_7_11_reg_out :
  1'd0;
assign cond_wire34_in =
  _guard1805 ? cond34_out :
  _guard1806 ? idx_between_9_13_reg_out :
  1'd0;
assign cond39_write_en = _guard1807;
assign cond39_clk = clk;
assign cond39_reset = reset;
assign cond39_in =
  _guard1808 ? idx_between_7_11_reg_out :
  1'd0;
assign cond49_write_en = _guard1809;
assign cond49_clk = clk;
assign cond49_reset = reset;
assign cond49_in =
  _guard1810 ? idx_between_6_10_reg_out :
  1'd0;
assign cond_wire52_in =
  _guard1813 ? cond52_out :
  _guard1814 ? idx_between_14_15_reg_out :
  1'd0;
assign cond_wire68_in =
  _guard1815 ? idx_between_15_16_reg_out :
  _guard1818 ? cond68_out :
  1'd0;
assign top_0_0_write_en = _guard1821;
assign top_0_0_clk = clk;
assign top_0_0_reset = reset;
assign top_0_0_in = t0_read_data;
assign pe_1_1_mul_ready =
  _guard1827 ? 1'd1 :
  _guard1830 ? 1'd0 :
  1'd0;
assign pe_1_1_clk = clk;
assign pe_1_1_top =
  _guard1843 ? top_1_1_out :
  32'd0;
assign pe_1_1_left =
  _guard1856 ? left_1_1_out :
  32'd0;
assign pe_1_1_reset = reset;
assign pe_1_1_go = _guard1869;
assign idx_between_8_12_comb_left = index_ge_8_out;
assign idx_between_8_12_comb_right = index_lt_12_out;
assign index_ge_13_left = idx_add_out;
assign index_ge_13_right = 5'd13;
assign idx_between_9_13_reg_write_en = _guard1878;
assign idx_between_9_13_reg_clk = clk;
assign idx_between_9_13_reg_reset = reset;
assign idx_between_9_13_reg_in =
  _guard1879 ? idx_between_9_13_comb_out :
  _guard1882 ? 1'd0 :
  'x;
assign idx_between_1_5_comb_left = index_ge_1_out;
assign idx_between_1_5_comb_right = index_lt_5_out;
assign idx_between_10_14_reg_write_en = _guard1889;
assign idx_between_10_14_reg_clk = clk;
assign idx_between_10_14_reg_reset = reset;
assign idx_between_10_14_reg_in =
  _guard1890 ? idx_between_10_14_comb_out :
  _guard1893 ? 1'd0 :
  'x;
assign idx_between_11_12_reg_write_en = _guard1898;
assign idx_between_11_12_reg_clk = clk;
assign idx_between_11_12_reg_reset = reset;
assign idx_between_11_12_reg_in =
  _guard1901 ? 1'd0 :
  _guard1902 ? idx_between_11_12_comb_out :
  'x;
assign idx_between_11_15_reg_write_en = _guard1907;
assign idx_between_11_15_reg_clk = clk;
assign idx_between_11_15_reg_reset = reset;
assign idx_between_11_15_reg_in =
  _guard1910 ? 1'd0 :
  _guard1911 ? idx_between_11_15_comb_out :
  'x;
assign cond_wire1_in =
  _guard1912 ? idx_between_1_5_reg_out :
  _guard1915 ? cond1_out :
  1'd0;
assign cond8_write_en = _guard1916;
assign cond8_clk = clk;
assign cond8_reset = reset;
assign cond8_in =
  _guard1917 ? idx_between_10_11_reg_out :
  1'd0;
assign cond12_write_en = _guard1918;
assign cond12_clk = clk;
assign cond12_reset = reset;
assign cond12_in =
  _guard1919 ? idx_between_7_11_reg_out :
  1'd0;
assign cond28_write_en = _guard1920;
assign cond28_clk = clk;
assign cond28_reset = reset;
assign cond28_in =
  _guard1921 ? idx_between_4_8_reg_out :
  1'd0;
assign cond_wire28_in =
  _guard1922 ? idx_between_4_8_reg_out :
  _guard1925 ? cond28_out :
  1'd0;
assign cond_wire53_in =
  _guard1926 ? idx_between_3_7_reg_out :
  _guard1929 ? cond53_out :
  1'd0;
assign cond55_write_en = _guard1930;
assign cond55_clk = clk;
assign cond55_reset = reset;
assign cond55_in =
  _guard1931 ? idx_between_4_8_reg_out :
  1'd0;
assign cond_wire65_in =
  _guard1934 ? cond65_out :
  _guard1935 ? idx_between_14_15_reg_out :
  1'd0;
assign wrapper_early_reset_static_seq_go_in = go;
assign left_0_1_write_en = _guard1938;
assign left_0_1_clk = clk;
assign left_0_1_reset = reset;
assign left_0_1_in = left_0_0_out;
assign pe_2_2_mul_ready =
  _guard1944 ? 1'd1 :
  _guard1947 ? 1'd0 :
  1'd0;
assign pe_2_2_clk = clk;
assign pe_2_2_top =
  _guard1960 ? top_2_2_out :
  32'd0;
assign pe_2_2_left =
  _guard1973 ? left_2_2_out :
  32'd0;
assign pe_2_2_reset = reset;
assign pe_2_2_go = _guard1986;
assign l2_add_left = 3'd1;
assign l2_add_right = l2_idx_out;
assign index_lt_14_left = idx_add_out;
assign index_lt_14_right = 5'd14;
assign index_lt_4_left = idx_add_out;
assign index_lt_4_right = 5'd4;
assign idx_between_2_6_reg_write_en = _guard2001;
assign idx_between_2_6_reg_clk = clk;
assign idx_between_2_6_reg_reset = reset;
assign idx_between_2_6_reg_in =
  _guard2004 ? 1'd0 :
  _guard2005 ? idx_between_2_6_comb_out :
  'x;
assign idx_between_2_6_comb_left = index_ge_2_out;
assign idx_between_2_6_comb_right = index_lt_6_out;
assign cond_wire14_in =
  _guard2008 ? idx_between_3_7_reg_out :
  _guard2011 ? cond14_out :
  1'd0;
assign cond_wire21_in =
  _guard2014 ? cond21_out :
  _guard2015 ? idx_between_2_6_reg_out :
  1'd0;
assign cond38_write_en = _guard2016;
assign cond38_clk = clk;
assign cond38_reset = reset;
assign cond38_in =
  _guard2017 ? idx_between_3_7_reg_out :
  1'd0;
assign cond42_write_en = _guard2018;
assign cond42_clk = clk;
assign cond42_reset = reset;
assign cond42_in =
  _guard2019 ? idx_between_4_8_reg_out :
  1'd0;
assign cond_wire51_in =
  _guard2022 ? cond51_out :
  _guard2023 ? idx_between_10_14_reg_out :
  1'd0;
assign cond59_write_en = _guard2024;
assign cond59_clk = clk;
assign cond59_reset = reset;
assign cond59_in =
  _guard2025 ? idx_between_5_9_reg_out :
  1'd0;
// COMPONENT END: main
endmodule

